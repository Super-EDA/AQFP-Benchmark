module sorter_48 ( a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ , b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ );
  input a_44_ , a_5_ , a_38_ , a_43_ , a_20_ , a_27_ , a_8_ , a_40_ , a_47_ , a_11_ , a_0_ , a_6_ , a_16_ , a_9_ , a_31_ , a_4_ , a_30_ , a_35_ , a_26_ , a_19_ , a_7_ , a_13_ , a_45_ , a_34_ , a_42_ , a_14_ , a_41_ , a_17_ , a_37_ , a_18_ , a_29_ , a_21_ , a_32_ , a_22_ , a_36_ , a_3_ , a_28_ , a_46_ , a_25_ , a_10_ , a_12_ , a_33_ , a_24_ , a_1_ , a_15_ , a_2_ , a_39_ , a_23_ ;
  output b_47_ , b_43_ , b_40_ , b_11_ , b_7_ , b_5_ , b_32_ , b_17_ , b_29_ , b_25_ , b_12_ , b_16_ , b_1_ , b_42_ , b_0_ , b_28_ , b_9_ , b_36_ , b_2_ , b_20_ , b_41_ , b_33_ , b_31_ , b_34_ , b_13_ , b_21_ , b_35_ , b_39_ , b_27_ , b_46_ , b_4_ , b_14_ , b_37_ , b_22_ , b_6_ , b_38_ , b_18_ , b_15_ , b_30_ , b_8_ , b_26_ , b_24_ , b_19_ , b_23_ , b_10_ , b_3_ , b_45_ , b_44_ ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 ;
  assign n49 = a_35_ & a_34_ ;
  assign n50 = a_33_ & n49 ;
  assign n51 = a_31_ | a_32_ ;
  assign n52 = a_30_ | n51 ;
  assign n53 = n50 & n52 ;
  assign n54 = a_35_ | a_34_ ;
  assign n55 = a_33_ | n54 ;
  assign n56 = a_31_ & a_32_ ;
  assign n57 = a_30_ & n56 ;
  assign n58 = n55 & n57 ;
  assign n59 = ( a_35_ & a_34_ ) | ( a_35_ & a_33_ ) | ( a_34_ & a_33_ ) ;
  assign n60 = ( a_31_ & a_30_ ) | ( a_31_ & a_32_ ) | ( a_30_ & a_32_ ) ;
  assign n61 = n59 & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n53 & n62 ;
  assign n64 = a_29_ & a_28_ ;
  assign n65 = a_27_ & n64 ;
  assign n66 = a_26_ | a_25_ ;
  assign n67 = a_24_ | n66 ;
  assign n68 = n65 | n67 ;
  assign n69 = ( a_27_ & a_29_ ) | ( a_27_ & a_28_ ) | ( a_29_ & a_28_ ) ;
  assign n70 = ( a_26_ & a_25_ ) | ( a_26_ & a_24_ ) | ( a_25_ & a_24_ ) ;
  assign n71 = n69 | n70 ;
  assign n72 = a_29_ | a_28_ ;
  assign n73 = a_27_ | n72 ;
  assign n74 = a_26_ & a_25_ ;
  assign n75 = a_24_ & n74 ;
  assign n76 = n73 | n75 ;
  assign n77 = n71 | n76 ;
  assign n78 = n68 | n77 ;
  assign n79 = n63 & n78 ;
  assign n80 = n50 | n52 ;
  assign n81 = n55 | n57 ;
  assign n82 = n59 | n60 ;
  assign n83 = n81 & n82 ;
  assign n84 = n80 & n83 ;
  assign n85 = n65 & n67 ;
  assign n86 = n69 & n70 ;
  assign n87 = n73 & n75 ;
  assign n88 = n86 | n87 ;
  assign n89 = n85 | n88 ;
  assign n90 = n84 & n89 ;
  assign n91 = n79 & n90 ;
  assign n92 = ( n53 & n58 ) | ( n53 & n61 ) | ( n58 & n61 ) ;
  assign n93 = ( n68 & n71 ) | ( n68 & n76 ) | ( n71 & n76 ) ;
  assign n94 = n92 & n93 ;
  assign n95 = ( n80 & n81 ) | ( n80 & n82 ) | ( n81 & n82 ) ;
  assign n96 = ( n85 & n86 ) | ( n85 & n87 ) | ( n86 & n87 ) ;
  assign n97 = n95 & n96 ;
  assign n98 = n94 & n97 ;
  assign n99 = n58 | n61 ;
  assign n100 = n53 | n99 ;
  assign n101 = n71 & n76 ;
  assign n102 = n68 & n101 ;
  assign n103 = n100 & n102 ;
  assign n104 = n81 | n82 ;
  assign n105 = n80 | n104 ;
  assign n106 = n86 & n87 ;
  assign n107 = n85 & n106 ;
  assign n108 = n105 & n107 ;
  assign n109 = n103 & n108 ;
  assign n110 = n98 & n109 ;
  assign n111 = n91 & n110 ;
  assign n112 = a_40_ & a_41_ ;
  assign n113 = a_39_ & n112 ;
  assign n114 = a_38_ | a_37_ ;
  assign n115 = a_36_ | n114 ;
  assign n116 = n113 & n115 ;
  assign n117 = a_40_ | a_41_ ;
  assign n118 = a_39_ | n117 ;
  assign n119 = a_38_ & a_37_ ;
  assign n120 = a_36_ & n119 ;
  assign n121 = n118 & n120 ;
  assign n122 = ( a_40_ & a_41_ ) | ( a_40_ & a_39_ ) | ( a_41_ & a_39_ ) ;
  assign n123 = ( a_38_ & a_37_ ) | ( a_38_ & a_36_ ) | ( a_37_ & a_36_ ) ;
  assign n124 = n122 & n123 ;
  assign n125 = n121 | n124 ;
  assign n126 = n116 | n125 ;
  assign n127 = ( a_44_ & a_43_ ) | ( a_44_ & a_42_ ) | ( a_43_ & a_42_ ) ;
  assign n128 = ( a_47_ & a_45_ ) | ( a_47_ & a_46_ ) | ( a_45_ & a_46_ ) ;
  assign n129 = n127 | n128 ;
  assign n130 = a_44_ & a_43_ ;
  assign n131 = a_42_ & n130 ;
  assign n132 = a_47_ | a_46_ ;
  assign n133 = a_45_ | n132 ;
  assign n134 = n131 | n133 ;
  assign n135 = n129 & n134 ;
  assign n136 = a_47_ & a_46_ ;
  assign n137 = a_45_ & n136 ;
  assign n138 = a_44_ | a_43_ ;
  assign n139 = a_42_ | n138 ;
  assign n140 = n137 | n139 ;
  assign n141 = n135 & n140 ;
  assign n142 = n126 | n141 ;
  assign n143 = n113 | n115 ;
  assign n144 = n118 | n120 ;
  assign n145 = n122 | n123 ;
  assign n146 = n144 | n145 ;
  assign n147 = n143 | n146 ;
  assign n148 = n127 & n128 ;
  assign n149 = n131 & n133 ;
  assign n150 = n148 & n149 ;
  assign n151 = n137 & n139 ;
  assign n152 = n150 & n151 ;
  assign n153 = n147 | n152 ;
  assign n154 = n142 | n153 ;
  assign n155 = n121 & n124 ;
  assign n156 = n116 & n155 ;
  assign n157 = n129 | n134 ;
  assign n158 = n140 | n157 ;
  assign n159 = n156 | n158 ;
  assign n160 = n144 & n145 ;
  assign n161 = n143 & n160 ;
  assign n162 = n148 | n149 ;
  assign n163 = n151 | n162 ;
  assign n164 = n161 | n163 ;
  assign n165 = n159 | n164 ;
  assign n166 = ( n116 & n121 ) | ( n116 & n124 ) | ( n121 & n124 ) ;
  assign n167 = ( n129 & n134 ) | ( n129 & n140 ) | ( n134 & n140 ) ;
  assign n168 = n166 | n167 ;
  assign n169 = ( n143 & n144 ) | ( n143 & n145 ) | ( n144 & n145 ) ;
  assign n170 = ( n148 & n149 ) | ( n148 & n151 ) | ( n149 & n151 ) ;
  assign n171 = n169 | n170 ;
  assign n172 = n168 | n171 ;
  assign n173 = n165 | n172 ;
  assign n174 = n154 | n173 ;
  assign n175 = n111 & n174 ;
  assign n176 = n63 | n78 ;
  assign n177 = n84 | n89 ;
  assign n178 = n176 & n177 ;
  assign n179 = n100 | n102 ;
  assign n180 = n105 | n107 ;
  assign n181 = n179 & n180 ;
  assign n182 = n92 | n93 ;
  assign n183 = n95 | n96 ;
  assign n184 = n182 & n183 ;
  assign n185 = n181 & n184 ;
  assign n186 = n178 & n185 ;
  assign n187 = n126 & n141 ;
  assign n188 = n147 & n152 ;
  assign n189 = n187 | n188 ;
  assign n190 = n156 & n158 ;
  assign n191 = n161 & n163 ;
  assign n192 = n190 | n191 ;
  assign n193 = n166 & n167 ;
  assign n194 = n169 & n170 ;
  assign n195 = n193 | n194 ;
  assign n196 = n192 | n195 ;
  assign n197 = n189 | n196 ;
  assign n198 = n186 & n197 ;
  assign n199 = n175 & n198 ;
  assign n200 = n79 | n90 ;
  assign n201 = n94 | n97 ;
  assign n202 = n103 | n108 ;
  assign n203 = n201 & n202 ;
  assign n204 = n200 & n203 ;
  assign n205 = n142 & n153 ;
  assign n206 = n159 & n164 ;
  assign n207 = n168 & n171 ;
  assign n208 = n206 | n207 ;
  assign n209 = n205 | n208 ;
  assign n210 = n204 & n209 ;
  assign n211 = n176 | n177 ;
  assign n212 = n179 | n180 ;
  assign n213 = n182 | n183 ;
  assign n214 = n212 & n213 ;
  assign n215 = n211 & n214 ;
  assign n216 = n187 & n188 ;
  assign n217 = n190 & n191 ;
  assign n218 = n193 & n194 ;
  assign n219 = n217 | n218 ;
  assign n220 = n216 | n219 ;
  assign n221 = n215 & n220 ;
  assign n222 = n210 & n221 ;
  assign n223 = n199 & n222 ;
  assign n224 = ( n91 & n98 ) | ( n91 & n109 ) | ( n98 & n109 ) ;
  assign n225 = ( n154 & n165 ) | ( n154 & n172 ) | ( n165 & n172 ) ;
  assign n226 = n224 & n225 ;
  assign n227 = ( n178 & n181 ) | ( n178 & n184 ) | ( n181 & n184 ) ;
  assign n228 = ( n189 & n192 ) | ( n189 & n195 ) | ( n192 & n195 ) ;
  assign n229 = n227 & n228 ;
  assign n230 = n226 & n229 ;
  assign n231 = ( n200 & n201 ) | ( n200 & n202 ) | ( n201 & n202 ) ;
  assign n232 = ( n205 & n206 ) | ( n205 & n207 ) | ( n206 & n207 ) ;
  assign n233 = n231 & n232 ;
  assign n234 = ( n211 & n212 ) | ( n211 & n213 ) | ( n212 & n213 ) ;
  assign n235 = ( n216 & n217 ) | ( n216 & n218 ) | ( n217 & n218 ) ;
  assign n236 = n234 & n235 ;
  assign n237 = n233 & n236 ;
  assign n238 = n230 & n237 ;
  assign n239 = n223 & n238 ;
  assign n240 = n98 | n109 ;
  assign n241 = n91 | n240 ;
  assign n242 = n165 & n172 ;
  assign n243 = n154 & n242 ;
  assign n244 = n241 & n243 ;
  assign n245 = n181 | n184 ;
  assign n246 = n178 | n245 ;
  assign n247 = n192 & n195 ;
  assign n248 = n189 & n247 ;
  assign n249 = n246 & n248 ;
  assign n250 = n244 & n249 ;
  assign n251 = n201 | n202 ;
  assign n252 = n200 | n251 ;
  assign n253 = n206 & n207 ;
  assign n254 = n205 & n253 ;
  assign n255 = n252 & n254 ;
  assign n256 = n212 | n213 ;
  assign n257 = n211 | n256 ;
  assign n258 = n217 & n218 ;
  assign n259 = n216 & n258 ;
  assign n260 = n257 & n259 ;
  assign n261 = n255 & n260 ;
  assign n262 = n250 & n261 ;
  assign n263 = n239 & n262 ;
  assign n264 = a_11_ & a_10_ ;
  assign n265 = a_9_ & n264 ;
  assign n266 = a_8_ | a_7_ ;
  assign n267 = a_6_ | n266 ;
  assign n268 = n265 & n267 ;
  assign n269 = a_11_ | a_10_ ;
  assign n270 = a_9_ | n269 ;
  assign n271 = a_8_ & a_7_ ;
  assign n272 = a_6_ & n271 ;
  assign n273 = n270 & n272 ;
  assign n274 = ( a_11_ & a_9_ ) | ( a_11_ & a_10_ ) | ( a_9_ & a_10_ ) ;
  assign n275 = ( a_8_ & a_6_ ) | ( a_8_ & a_7_ ) | ( a_6_ & a_7_ ) ;
  assign n276 = n274 & n275 ;
  assign n277 = n273 & n276 ;
  assign n278 = n268 & n277 ;
  assign n279 = a_5_ & a_4_ ;
  assign n280 = a_3_ & n279 ;
  assign n281 = a_1_ | a_2_ ;
  assign n282 = a_0_ | n281 ;
  assign n283 = n280 | n282 ;
  assign n284 = a_5_ | a_4_ ;
  assign n285 = a_3_ | n284 ;
  assign n286 = a_1_ & a_2_ ;
  assign n287 = a_0_ & n286 ;
  assign n288 = n285 | n287 ;
  assign n289 = ( a_5_ & a_4_ ) | ( a_5_ & a_3_ ) | ( a_4_ & a_3_ ) ;
  assign n290 = ( a_0_ & a_1_ ) | ( a_0_ & a_2_ ) | ( a_1_ & a_2_ ) ;
  assign n291 = n289 | n290 ;
  assign n292 = n288 | n291 ;
  assign n293 = n283 | n292 ;
  assign n294 = n278 & n293 ;
  assign n295 = n265 | n267 ;
  assign n296 = n270 | n272 ;
  assign n297 = n274 | n275 ;
  assign n298 = n296 & n297 ;
  assign n299 = n295 & n298 ;
  assign n300 = n280 & n282 ;
  assign n301 = n285 & n287 ;
  assign n302 = n289 & n290 ;
  assign n303 = n301 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = n299 & n304 ;
  assign n306 = n294 & n305 ;
  assign n307 = n273 | n276 ;
  assign n308 = n268 | n307 ;
  assign n309 = n288 & n291 ;
  assign n310 = n283 & n309 ;
  assign n311 = n308 & n310 ;
  assign n312 = n296 | n297 ;
  assign n313 = n295 | n312 ;
  assign n314 = n301 & n302 ;
  assign n315 = n300 & n314 ;
  assign n316 = n313 & n315 ;
  assign n317 = n311 & n316 ;
  assign n318 = ( n268 & n273 ) | ( n268 & n276 ) | ( n273 & n276 ) ;
  assign n319 = ( n283 & n288 ) | ( n283 & n291 ) | ( n288 & n291 ) ;
  assign n320 = n318 & n319 ;
  assign n321 = ( n295 & n296 ) | ( n295 & n297 ) | ( n296 & n297 ) ;
  assign n322 = ( n300 & n301 ) | ( n300 & n302 ) | ( n301 & n302 ) ;
  assign n323 = n321 & n322 ;
  assign n324 = n320 & n323 ;
  assign n325 = n317 & n324 ;
  assign n326 = n306 & n325 ;
  assign n327 = a_22_ & a_23_ ;
  assign n328 = a_21_ & n327 ;
  assign n329 = a_20_ | a_19_ ;
  assign n330 = a_18_ | n329 ;
  assign n331 = n328 | n330 ;
  assign n332 = a_22_ | a_23_ ;
  assign n333 = a_21_ | n332 ;
  assign n334 = a_20_ & a_19_ ;
  assign n335 = a_18_ & n334 ;
  assign n336 = n333 | n335 ;
  assign n337 = ( a_21_ & a_22_ ) | ( a_21_ & a_23_ ) | ( a_22_ & a_23_ ) ;
  assign n338 = ( a_20_ & a_19_ ) | ( a_20_ & a_18_ ) | ( a_19_ & a_18_ ) ;
  assign n339 = n337 | n338 ;
  assign n340 = n336 & n339 ;
  assign n341 = n331 & n340 ;
  assign n342 = a_16_ & a_17_ ;
  assign n343 = a_15_ & n342 ;
  assign n344 = a_13_ | a_14_ ;
  assign n345 = a_12_ | n344 ;
  assign n346 = n343 & n345 ;
  assign n347 = a_16_ | a_17_ ;
  assign n348 = a_15_ | n347 ;
  assign n349 = a_13_ & a_14_ ;
  assign n350 = a_12_ & n349 ;
  assign n351 = n348 & n350 ;
  assign n352 = ( a_16_ & a_17_ ) | ( a_16_ & a_15_ ) | ( a_17_ & a_15_ ) ;
  assign n353 = ( a_13_ & a_14_ ) | ( a_13_ & a_12_ ) | ( a_14_ & a_12_ ) ;
  assign n354 = n352 & n353 ;
  assign n355 = n351 | n354 ;
  assign n356 = n346 | n355 ;
  assign n357 = n341 | n356 ;
  assign n358 = n328 & n330 ;
  assign n359 = n333 & n335 ;
  assign n360 = n337 & n338 ;
  assign n361 = n359 & n360 ;
  assign n362 = n358 & n361 ;
  assign n363 = n348 | n350 ;
  assign n364 = n352 | n353 ;
  assign n365 = n363 | n364 ;
  assign n366 = n343 | n345 ;
  assign n367 = n365 | n366 ;
  assign n368 = n362 | n367 ;
  assign n369 = n357 | n368 ;
  assign n370 = n336 | n339 ;
  assign n371 = n331 | n370 ;
  assign n372 = n351 & n354 ;
  assign n373 = n346 & n372 ;
  assign n374 = n371 | n373 ;
  assign n375 = n359 | n360 ;
  assign n376 = n358 | n375 ;
  assign n377 = n363 & n364 ;
  assign n378 = n366 & n377 ;
  assign n379 = n376 | n378 ;
  assign n380 = n374 | n379 ;
  assign n381 = ( n331 & n336 ) | ( n331 & n339 ) | ( n336 & n339 ) ;
  assign n382 = ( n346 & n351 ) | ( n346 & n354 ) | ( n351 & n354 ) ;
  assign n383 = n381 | n382 ;
  assign n384 = ( n358 & n359 ) | ( n358 & n360 ) | ( n359 & n360 ) ;
  assign n385 = ( n363 & n364 ) | ( n363 & n366 ) | ( n364 & n366 ) ;
  assign n386 = n384 | n385 ;
  assign n387 = n383 | n386 ;
  assign n388 = n380 | n387 ;
  assign n389 = n369 | n388 ;
  assign n390 = n326 | n389 ;
  assign n391 = n278 | n293 ;
  assign n392 = n299 | n304 ;
  assign n393 = n391 & n392 ;
  assign n394 = n318 | n319 ;
  assign n395 = n321 | n322 ;
  assign n396 = n394 & n395 ;
  assign n397 = n308 | n310 ;
  assign n398 = n313 | n315 ;
  assign n399 = n397 & n398 ;
  assign n400 = n396 & n399 ;
  assign n401 = n393 & n400 ;
  assign n402 = n341 & n356 ;
  assign n403 = n362 & n367 ;
  assign n404 = n402 | n403 ;
  assign n405 = n371 & n373 ;
  assign n406 = n376 & n378 ;
  assign n407 = n405 | n406 ;
  assign n408 = n381 & n382 ;
  assign n409 = n384 & n385 ;
  assign n410 = n408 | n409 ;
  assign n411 = n407 | n410 ;
  assign n412 = n404 | n411 ;
  assign n413 = n401 | n412 ;
  assign n414 = n390 | n413 ;
  assign n415 = n311 | n316 ;
  assign n416 = n320 | n323 ;
  assign n417 = n415 & n416 ;
  assign n418 = n294 | n305 ;
  assign n419 = n417 & n418 ;
  assign n420 = n357 & n368 ;
  assign n421 = n374 & n379 ;
  assign n422 = n383 & n386 ;
  assign n423 = n421 | n422 ;
  assign n424 = n420 | n423 ;
  assign n425 = n419 | n424 ;
  assign n426 = n391 | n392 ;
  assign n427 = n394 | n395 ;
  assign n428 = n397 | n398 ;
  assign n429 = n427 & n428 ;
  assign n430 = n426 & n429 ;
  assign n431 = n402 & n403 ;
  assign n432 = n405 & n406 ;
  assign n433 = n408 & n409 ;
  assign n434 = n432 | n433 ;
  assign n435 = n431 | n434 ;
  assign n436 = n430 | n435 ;
  assign n437 = n425 | n436 ;
  assign n438 = n414 | n437 ;
  assign n439 = ( n306 & n317 ) | ( n306 & n324 ) | ( n317 & n324 ) ;
  assign n440 = ( n369 & n380 ) | ( n369 & n387 ) | ( n380 & n387 ) ;
  assign n441 = n439 | n440 ;
  assign n442 = ( n393 & n396 ) | ( n393 & n399 ) | ( n396 & n399 ) ;
  assign n443 = ( n404 & n407 ) | ( n404 & n410 ) | ( n407 & n410 ) ;
  assign n444 = n442 | n443 ;
  assign n445 = n441 | n444 ;
  assign n446 = ( n415 & n416 ) | ( n415 & n418 ) | ( n416 & n418 ) ;
  assign n447 = ( n420 & n421 ) | ( n420 & n422 ) | ( n421 & n422 ) ;
  assign n448 = n446 | n447 ;
  assign n449 = ( n426 & n427 ) | ( n426 & n428 ) | ( n427 & n428 ) ;
  assign n450 = ( n431 & n432 ) | ( n431 & n433 ) | ( n432 & n433 ) ;
  assign n451 = n449 | n450 ;
  assign n452 = n448 | n451 ;
  assign n453 = n445 | n452 ;
  assign n454 = n438 | n453 ;
  assign n455 = n317 | n324 ;
  assign n456 = n306 | n455 ;
  assign n457 = n380 & n387 ;
  assign n458 = n369 & n457 ;
  assign n459 = n456 | n458 ;
  assign n460 = n396 | n399 ;
  assign n461 = n393 | n460 ;
  assign n462 = n407 & n410 ;
  assign n463 = n404 & n462 ;
  assign n464 = n461 | n463 ;
  assign n465 = n459 | n464 ;
  assign n466 = n415 | n416 ;
  assign n467 = n418 | n466 ;
  assign n468 = n421 & n422 ;
  assign n469 = n420 & n468 ;
  assign n470 = n467 | n469 ;
  assign n471 = n427 | n428 ;
  assign n472 = n426 | n471 ;
  assign n473 = n432 & n433 ;
  assign n474 = n431 & n473 ;
  assign n475 = n472 | n474 ;
  assign n476 = n470 | n475 ;
  assign n477 = n465 | n476 ;
  assign n478 = n454 | n477 ;
  assign n479 = n263 | n478 ;
  assign n480 = n111 | n174 ;
  assign n481 = n186 | n197 ;
  assign n482 = n480 & n481 ;
  assign n483 = n204 | n209 ;
  assign n484 = n215 | n220 ;
  assign n485 = n483 & n484 ;
  assign n486 = n482 & n485 ;
  assign n487 = n224 | n225 ;
  assign n488 = n227 | n228 ;
  assign n489 = n487 & n488 ;
  assign n490 = n231 | n232 ;
  assign n491 = n234 | n235 ;
  assign n492 = n490 & n491 ;
  assign n493 = n489 & n492 ;
  assign n494 = n486 & n493 ;
  assign n495 = n241 | n243 ;
  assign n496 = n246 | n248 ;
  assign n497 = n495 & n496 ;
  assign n498 = n252 | n254 ;
  assign n499 = n257 | n259 ;
  assign n500 = n498 & n499 ;
  assign n501 = n497 & n500 ;
  assign n502 = n494 & n501 ;
  assign n503 = n326 & n389 ;
  assign n504 = n401 & n412 ;
  assign n505 = n503 | n504 ;
  assign n506 = n419 & n424 ;
  assign n507 = n430 & n435 ;
  assign n508 = n506 | n507 ;
  assign n509 = n505 | n508 ;
  assign n510 = n439 & n440 ;
  assign n511 = n442 & n443 ;
  assign n512 = n510 | n511 ;
  assign n513 = n446 & n447 ;
  assign n514 = n449 & n450 ;
  assign n515 = n513 | n514 ;
  assign n516 = n512 | n515 ;
  assign n517 = n509 | n516 ;
  assign n518 = n456 & n458 ;
  assign n519 = n461 & n463 ;
  assign n520 = n518 | n519 ;
  assign n521 = n467 & n469 ;
  assign n522 = n472 & n474 ;
  assign n523 = n521 | n522 ;
  assign n524 = n520 | n523 ;
  assign n525 = n517 | n524 ;
  assign n526 = n502 | n525 ;
  assign n527 = n479 | n526 ;
  assign n528 = n175 | n198 ;
  assign n529 = n210 | n221 ;
  assign n530 = n528 & n529 ;
  assign n531 = n226 | n229 ;
  assign n532 = n233 | n236 ;
  assign n533 = n531 & n532 ;
  assign n534 = n530 & n533 ;
  assign n535 = n244 | n249 ;
  assign n536 = n255 | n260 ;
  assign n537 = n535 & n536 ;
  assign n538 = n534 & n537 ;
  assign n539 = n390 & n413 ;
  assign n540 = n425 & n436 ;
  assign n541 = n539 | n540 ;
  assign n542 = n441 & n444 ;
  assign n543 = n448 & n451 ;
  assign n544 = n542 | n543 ;
  assign n545 = n541 | n544 ;
  assign n546 = n459 & n464 ;
  assign n547 = n470 & n475 ;
  assign n548 = n546 | n547 ;
  assign n549 = n545 | n548 ;
  assign n550 = n538 | n549 ;
  assign n551 = n480 | n481 ;
  assign n552 = n483 | n484 ;
  assign n553 = n551 & n552 ;
  assign n554 = n487 | n488 ;
  assign n555 = n490 | n491 ;
  assign n556 = n554 & n555 ;
  assign n557 = n553 & n556 ;
  assign n558 = n495 | n496 ;
  assign n559 = n498 | n499 ;
  assign n560 = n558 & n559 ;
  assign n561 = n557 & n560 ;
  assign n562 = n503 & n504 ;
  assign n563 = n506 & n507 ;
  assign n564 = n562 | n563 ;
  assign n565 = n510 & n511 ;
  assign n566 = n513 & n514 ;
  assign n567 = n565 | n566 ;
  assign n568 = n564 | n567 ;
  assign n569 = n518 & n519 ;
  assign n570 = n521 & n522 ;
  assign n571 = n569 | n570 ;
  assign n572 = n568 | n571 ;
  assign n573 = n561 | n572 ;
  assign n574 = n550 | n573 ;
  assign n575 = n527 | n574 ;
  assign n576 = n199 | n222 ;
  assign n577 = n230 | n237 ;
  assign n578 = n576 & n577 ;
  assign n579 = n250 | n261 ;
  assign n580 = n578 & n579 ;
  assign n581 = n414 & n437 ;
  assign n582 = n445 & n452 ;
  assign n583 = n581 | n582 ;
  assign n584 = n465 & n476 ;
  assign n585 = n583 | n584 ;
  assign n586 = n580 | n585 ;
  assign n587 = n482 | n485 ;
  assign n588 = n489 | n492 ;
  assign n589 = n587 & n588 ;
  assign n590 = n497 | n500 ;
  assign n591 = n589 & n590 ;
  assign n592 = n505 & n508 ;
  assign n593 = n512 & n515 ;
  assign n594 = n592 | n593 ;
  assign n595 = n520 & n523 ;
  assign n596 = n594 | n595 ;
  assign n597 = n591 | n596 ;
  assign n598 = n586 | n597 ;
  assign n599 = n528 | n529 ;
  assign n600 = n531 | n532 ;
  assign n601 = n599 & n600 ;
  assign n602 = n535 | n536 ;
  assign n603 = n601 & n602 ;
  assign n604 = n539 & n540 ;
  assign n605 = n542 & n543 ;
  assign n606 = n604 | n605 ;
  assign n607 = n546 & n547 ;
  assign n608 = n606 | n607 ;
  assign n609 = n603 | n608 ;
  assign n610 = n551 | n552 ;
  assign n611 = n554 | n555 ;
  assign n612 = n610 & n611 ;
  assign n613 = n558 | n559 ;
  assign n614 = n612 & n613 ;
  assign n615 = n562 & n563 ;
  assign n616 = n565 & n566 ;
  assign n617 = n615 | n616 ;
  assign n618 = n569 & n570 ;
  assign n619 = n617 | n618 ;
  assign n620 = n614 | n619 ;
  assign n621 = n609 | n620 ;
  assign n622 = n598 | n621 ;
  assign n623 = n575 | n622 ;
  assign n624 = ( n223 & n238 ) | ( n223 & n262 ) | ( n238 & n262 ) ;
  assign n625 = ( n438 & n453 ) | ( n438 & n477 ) | ( n453 & n477 ) ;
  assign n626 = n624 | n625 ;
  assign n627 = ( n486 & n493 ) | ( n486 & n501 ) | ( n493 & n501 ) ;
  assign n628 = ( n509 & n516 ) | ( n509 & n524 ) | ( n516 & n524 ) ;
  assign n629 = n627 | n628 ;
  assign n630 = n626 | n629 ;
  assign n631 = ( n530 & n533 ) | ( n530 & n537 ) | ( n533 & n537 ) ;
  assign n632 = ( n541 & n544 ) | ( n541 & n548 ) | ( n544 & n548 ) ;
  assign n633 = n631 | n632 ;
  assign n634 = ( n553 & n556 ) | ( n553 & n560 ) | ( n556 & n560 ) ;
  assign n635 = ( n564 & n567 ) | ( n564 & n571 ) | ( n567 & n571 ) ;
  assign n636 = n634 | n635 ;
  assign n637 = n633 | n636 ;
  assign n638 = n630 | n637 ;
  assign n639 = ( n576 & n577 ) | ( n576 & n579 ) | ( n577 & n579 ) ;
  assign n640 = ( n581 & n582 ) | ( n581 & n584 ) | ( n582 & n584 ) ;
  assign n641 = n639 | n640 ;
  assign n642 = ( n587 & n588 ) | ( n587 & n590 ) | ( n588 & n590 ) ;
  assign n643 = ( n592 & n593 ) | ( n592 & n595 ) | ( n593 & n595 ) ;
  assign n644 = n642 | n643 ;
  assign n645 = n641 | n644 ;
  assign n646 = ( n599 & n600 ) | ( n599 & n602 ) | ( n600 & n602 ) ;
  assign n647 = ( n604 & n605 ) | ( n604 & n607 ) | ( n605 & n607 ) ;
  assign n648 = n646 | n647 ;
  assign n649 = ( n610 & n611 ) | ( n610 & n613 ) | ( n611 & n613 ) ;
  assign n650 = ( n615 & n616 ) | ( n615 & n618 ) | ( n616 & n618 ) ;
  assign n651 = n649 | n650 ;
  assign n652 = n648 | n651 ;
  assign n653 = n645 | n652 ;
  assign n654 = n638 | n653 ;
  assign n655 = n223 | n238 ;
  assign n656 = n262 | n655 ;
  assign n657 = n438 & n453 ;
  assign n658 = n477 & n657 ;
  assign n659 = n656 | n658 ;
  assign n660 = n486 | n493 ;
  assign n661 = n501 | n660 ;
  assign n662 = n509 & n516 ;
  assign n663 = n524 & n662 ;
  assign n664 = n661 | n663 ;
  assign n665 = n659 | n664 ;
  assign n666 = n530 | n533 ;
  assign n667 = n537 | n666 ;
  assign n668 = n541 & n544 ;
  assign n669 = n548 & n668 ;
  assign n670 = n667 | n669 ;
  assign n671 = n553 | n556 ;
  assign n672 = n560 | n671 ;
  assign n673 = n564 & n567 ;
  assign n674 = n571 & n673 ;
  assign n675 = n672 | n674 ;
  assign n676 = n670 | n675 ;
  assign n677 = n665 | n676 ;
  assign n678 = n576 | n577 ;
  assign n679 = n579 | n678 ;
  assign n680 = n581 & n582 ;
  assign n681 = n584 & n680 ;
  assign n682 = n679 | n681 ;
  assign n683 = n587 | n588 ;
  assign n684 = n590 | n683 ;
  assign n685 = n592 & n593 ;
  assign n686 = n595 & n685 ;
  assign n687 = n684 | n686 ;
  assign n688 = n682 | n687 ;
  assign n689 = n599 | n600 ;
  assign n690 = n602 | n689 ;
  assign n691 = n604 & n605 ;
  assign n692 = n607 & n691 ;
  assign n693 = n690 | n692 ;
  assign n694 = n610 | n611 ;
  assign n695 = n613 | n694 ;
  assign n696 = n615 & n616 ;
  assign n697 = n618 & n696 ;
  assign n698 = n695 | n697 ;
  assign n699 = n693 | n698 ;
  assign n700 = n688 | n699 ;
  assign n701 = n677 | n700 ;
  assign n702 = n654 | n701 ;
  assign n703 = n623 | n702 ;
  assign n704 = n575 & n622 ;
  assign n705 = n638 & n653 ;
  assign n706 = n677 & n700 ;
  assign n707 = ( n704 & n705 ) | ( n704 & n706 ) | ( n705 & n706 ) ;
  assign n708 = n527 & n574 ;
  assign n709 = n598 & n621 ;
  assign n710 = n708 | n709 ;
  assign n711 = n630 & n637 ;
  assign n712 = n645 & n652 ;
  assign n713 = n711 | n712 ;
  assign n714 = n665 & n676 ;
  assign n715 = n688 & n699 ;
  assign n716 = n714 | n715 ;
  assign n717 = ( n710 & n713 ) | ( n710 & n716 ) | ( n713 & n716 ) ;
  assign n718 = n263 & n478 ;
  assign n719 = n502 & n525 ;
  assign n720 = n718 & n719 ;
  assign n721 = n538 & n549 ;
  assign n722 = n561 & n572 ;
  assign n723 = n721 & n722 ;
  assign n724 = n720 | n723 ;
  assign n725 = n580 & n585 ;
  assign n726 = n591 & n596 ;
  assign n727 = n725 & n726 ;
  assign n728 = n603 & n608 ;
  assign n729 = n614 & n619 ;
  assign n730 = n728 & n729 ;
  assign n731 = n727 | n730 ;
  assign n732 = n724 | n731 ;
  assign n733 = n624 & n625 ;
  assign n734 = n627 & n628 ;
  assign n735 = n733 & n734 ;
  assign n736 = n631 & n632 ;
  assign n737 = n634 & n635 ;
  assign n738 = n736 & n737 ;
  assign n739 = n735 | n738 ;
  assign n740 = n639 & n640 ;
  assign n741 = n642 & n643 ;
  assign n742 = n740 & n741 ;
  assign n743 = n646 & n647 ;
  assign n744 = n649 & n650 ;
  assign n745 = n743 & n744 ;
  assign n746 = n742 | n745 ;
  assign n747 = n739 | n746 ;
  assign n748 = n656 & n658 ;
  assign n749 = n661 & n663 ;
  assign n750 = n748 & n749 ;
  assign n751 = n667 & n669 ;
  assign n752 = n672 & n674 ;
  assign n753 = n751 & n752 ;
  assign n754 = n750 | n753 ;
  assign n755 = n679 & n681 ;
  assign n756 = n684 & n686 ;
  assign n757 = n755 & n756 ;
  assign n758 = n690 & n692 ;
  assign n759 = n695 & n697 ;
  assign n760 = n758 & n759 ;
  assign n761 = n757 | n760 ;
  assign n762 = n754 | n761 ;
  assign n763 = n747 | n762 ;
  assign n764 = n732 | n763 ;
  assign n765 = n724 & n731 ;
  assign n766 = n739 & n746 ;
  assign n767 = n754 & n761 ;
  assign n768 = ( n765 & n766 ) | ( n765 & n767 ) | ( n766 & n767 ) ;
  assign n769 = n720 & n723 ;
  assign n770 = n727 & n730 ;
  assign n771 = n769 | n770 ;
  assign n772 = n735 & n738 ;
  assign n773 = n742 & n745 ;
  assign n774 = n772 | n773 ;
  assign n775 = n750 & n753 ;
  assign n776 = n757 & n760 ;
  assign n777 = n775 | n776 ;
  assign n778 = n774 | n777 ;
  assign n779 = n771 | n778 ;
  assign n780 = n479 & n526 ;
  assign n781 = n550 & n573 ;
  assign n782 = n780 | n781 ;
  assign n783 = n586 & n597 ;
  assign n784 = n609 & n620 ;
  assign n785 = n783 | n784 ;
  assign n786 = n782 & n785 ;
  assign n787 = n626 & n629 ;
  assign n788 = n633 & n636 ;
  assign n789 = n787 | n788 ;
  assign n790 = n641 & n644 ;
  assign n791 = n648 & n651 ;
  assign n792 = n790 | n791 ;
  assign n793 = n789 & n792 ;
  assign n794 = n659 & n664 ;
  assign n795 = n670 & n675 ;
  assign n796 = n794 | n795 ;
  assign n797 = n682 & n687 ;
  assign n798 = n693 & n698 ;
  assign n799 = n797 | n798 ;
  assign n800 = n796 & n799 ;
  assign n801 = n793 | n800 ;
  assign n802 = n786 | n801 ;
  assign n803 = n718 | n719 ;
  assign n804 = n721 | n722 ;
  assign n805 = n803 & n804 ;
  assign n806 = n725 | n726 ;
  assign n807 = n728 | n729 ;
  assign n808 = n806 & n807 ;
  assign n809 = n805 | n808 ;
  assign n810 = n733 | n734 ;
  assign n811 = n736 | n737 ;
  assign n812 = n810 & n811 ;
  assign n813 = n740 | n741 ;
  assign n814 = n743 | n744 ;
  assign n815 = n813 & n814 ;
  assign n816 = n812 | n815 ;
  assign n817 = n748 | n749 ;
  assign n818 = n751 | n752 ;
  assign n819 = n817 & n818 ;
  assign n820 = n755 | n756 ;
  assign n821 = n758 | n759 ;
  assign n822 = n820 & n821 ;
  assign n823 = n819 | n822 ;
  assign n824 = n816 | n823 ;
  assign n825 = n809 | n824 ;
  assign n826 = n780 & n781 ;
  assign n827 = n783 & n784 ;
  assign n828 = n826 | n827 ;
  assign n829 = n787 & n788 ;
  assign n830 = n790 & n791 ;
  assign n831 = n829 | n830 ;
  assign n832 = n794 & n795 ;
  assign n833 = n797 & n798 ;
  assign n834 = n832 | n833 ;
  assign n835 = n831 | n834 ;
  assign n836 = n828 | n835 ;
  assign n837 = n826 & n827 ;
  assign n838 = n829 & n830 ;
  assign n839 = n832 & n833 ;
  assign n840 = ( n837 & n838 ) | ( n837 & n839 ) | ( n838 & n839 ) ;
  assign n841 = n805 & n808 ;
  assign n842 = n812 & n815 ;
  assign n843 = n819 & n822 ;
  assign n844 = n842 & n843 ;
  assign n845 = n841 & n844 ;
  assign n846 = ( n809 & n816 ) | ( n809 & n823 ) | ( n816 & n823 ) ;
  assign n847 = n769 & n770 ;
  assign n848 = n772 & n773 ;
  assign n849 = n775 & n776 ;
  assign n850 = ( n847 & n848 ) | ( n847 & n849 ) | ( n848 & n849 ) ;
  assign n851 = n705 & n706 ;
  assign n852 = n704 & n851 ;
  assign n853 = n848 & n849 ;
  assign n854 = n847 & n853 ;
  assign n855 = ( n828 & n831 ) | ( n828 & n834 ) | ( n831 & n834 ) ;
  assign n856 = n747 & n762 ;
  assign n857 = n732 & n856 ;
  assign n858 = n708 & n709 ;
  assign n859 = n711 & n712 ;
  assign n860 = n714 & n715 ;
  assign n861 = n859 & n860 ;
  assign n862 = n858 & n861 ;
  assign n863 = n848 | n849 ;
  assign n864 = n847 | n863 ;
  assign n865 = n803 | n804 ;
  assign n866 = n806 | n807 ;
  assign n867 = n865 & n866 ;
  assign n868 = n810 | n811 ;
  assign n869 = n813 | n814 ;
  assign n870 = n868 & n869 ;
  assign n871 = n817 | n818 ;
  assign n872 = n820 | n821 ;
  assign n873 = n871 & n872 ;
  assign n874 = n870 | n873 ;
  assign n875 = n867 | n874 ;
  assign n876 = n713 | n716 ;
  assign n877 = n710 | n876 ;
  assign n878 = n782 | n785 ;
  assign n879 = n789 | n792 ;
  assign n880 = n796 | n799 ;
  assign n881 = n879 & n880 ;
  assign n882 = n878 & n881 ;
  assign n883 = ( n786 & n793 ) | ( n786 & n800 ) | ( n793 & n800 ) ;
  assign n884 = ( n878 & n879 ) | ( n878 & n880 ) | ( n879 & n880 ) ;
  assign n885 = ( n841 & n842 ) | ( n841 & n843 ) | ( n842 & n843 ) ;
  assign n886 = n865 | n866 ;
  assign n887 = n868 | n869 ;
  assign n888 = n871 | n872 ;
  assign n889 = n887 & n888 ;
  assign n890 = n886 & n889 ;
  assign n891 = n879 | n880 ;
  assign n892 = n878 | n891 ;
  assign n893 = n713 & n716 ;
  assign n894 = n710 & n893 ;
  assign n895 = n831 & n834 ;
  assign n896 = n828 & n895 ;
  assign n897 = ( n623 & n654 ) | ( n623 & n701 ) | ( n654 & n701 ) ;
  assign n898 = ( n771 & n774 ) | ( n771 & n777 ) | ( n774 & n777 ) ;
  assign n899 = n842 | n843 ;
  assign n900 = n841 | n899 ;
  assign n901 = ( n858 & n859 ) | ( n858 & n860 ) | ( n859 & n860 ) ;
  assign n902 = ( n886 & n887 ) | ( n886 & n888 ) | ( n887 & n888 ) ;
  assign n903 = n766 & n767 ;
  assign n904 = n765 & n903 ;
  assign n905 = n859 | n860 ;
  assign n906 = n858 | n905 ;
  assign n907 = n870 & n873 ;
  assign n908 = n867 & n907 ;
  assign n909 = n816 & n823 ;
  assign n910 = n809 & n909 ;
  assign n911 = n793 & n800 ;
  assign n912 = n786 & n911 ;
  assign n913 = n766 | n767 ;
  assign n914 = n765 | n913 ;
  assign n915 = n838 | n839 ;
  assign n916 = n837 | n915 ;
  assign n917 = n838 & n839 ;
  assign n918 = n837 & n917 ;
  assign n919 = ( n867 & n870 ) | ( n867 & n873 ) | ( n870 & n873 ) ;
  assign n920 = n887 | n888 ;
  assign n921 = n886 | n920 ;
  assign n922 = ( n732 & n747 ) | ( n732 & n762 ) | ( n747 & n762 ) ;
  assign n923 = n774 & n777 ;
  assign n924 = n771 & n923 ;
  assign n925 = n654 & n701 ;
  assign n926 = n623 & n925 ;
  assign n927 = n705 | n706 ;
  assign n928 = n704 | n927 ;
  assign b_47_ = n703 ;
  assign b_43_ = n707 ;
  assign b_40_ = n717 ;
  assign b_11_ = n764 ;
  assign b_7_ = n768 ;
  assign b_5_ = n779 ;
  assign b_32_ = n802 ;
  assign b_17_ = n825 ;
  assign b_29_ = n836 ;
  assign b_25_ = n840 ;
  assign b_12_ = n845 ;
  assign b_16_ = n846 ;
  assign b_1_ = n850 ;
  assign b_42_ = n852 ;
  assign b_0_ = n854 ;
  assign b_28_ = n855 ;
  assign b_9_ = n857 ;
  assign b_36_ = n862 ;
  assign b_2_ = n864 ;
  assign b_20_ = n875 ;
  assign b_41_ = n877 ;
  assign b_33_ = n882 ;
  assign b_31_ = n883 ;
  assign b_34_ = n884 ;
  assign b_13_ = n885 ;
  assign b_21_ = n890 ;
  assign b_35_ = n892 ;
  assign b_39_ = n894 ;
  assign b_27_ = n896 ;
  assign b_46_ = n897 ;
  assign b_4_ = n898 ;
  assign b_14_ = n900 ;
  assign b_37_ = n901 ;
  assign b_22_ = n902 ;
  assign b_6_ = n904 ;
  assign b_38_ = n906 ;
  assign b_18_ = n908 ;
  assign b_15_ = n910 ;
  assign b_30_ = n912 ;
  assign b_8_ = n914 ;
  assign b_26_ = n916 ;
  assign b_24_ = n918 ;
  assign b_19_ = n919 ;
  assign b_23_ = n921 ;
  assign b_10_ = n922 ;
  assign b_3_ = n924 ;
  assign b_45_ = n926 ;
  assign b_44_ = n928 ;
endmodule