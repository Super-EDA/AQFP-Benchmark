module multiplier (
    a_0,
    a_1,
    a_2,
    a_3,
    a_4,
    a_5,
    a_6,
    a_7,
    b_0,
    b_1,
    b_2,
    b_3,
    b_4,
    b_5,
    b_6,
    b_7,
    s_0,
    s_1,
    s_2,
    s_3,
    s_4,
    s_5,
    s_6,
    s_7,
    s_8,
    s_9,
    s_10,
    s_11,
    s_12,
    s_13,
    s_14,
    s_15
);
  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;
  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  output s_0;
  output s_1;
  output s_2;
  output s_3;
  output s_4;
  output s_5;
  output s_6;
  output s_7;
  output s_8;
  output s_9;
  output s_10;
  output s_11;
  output s_12;
  output s_13;
  output s_14;
  output s_15;
  wire n17;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  assign n17  = a_1 & b_0;
  assign n18  = b_1 & a_0;
  assign n19  = n17 & n18;
  assign n20  = n17 | n18;
  assign n21  = ~n19 & n20;
  assign n22  = a_1 & b_6;
  assign n23  = b_4 & a_2;
  assign n24  = b_3 & a_3;
  assign n25  = n23 & n24;
  assign n26  = a_1 & b_5;
  assign n27  = n23 | n24;
  assign n28  = ~n25 & n27;
  assign n29  = n26 & n28;
  assign n30  = n25 | n29;
  assign n31  = n22 & n30;
  assign n32  = b_7 & a_0;
  assign n33  = n22 | n30;
  assign n34  = ~n31 & n33;
  assign n35  = n32 & n34;
  assign n36  = n31 | n35;
  assign n37  = a_1 & b_7;
  assign n38  = a_2 & b_6;
  assign n39  = b_4 & a_3;
  assign n40  = a_4 & b_3;
  assign n41  = n39 & n40;
  assign n42  = n39 | n40;
  assign n43  = ~n41 & n42;
  assign n44  = a_2 & b_5;
  assign n45  = n43 & n44;
  assign n46  = n41 | n45;
  assign n47  = n38 & n46;
  assign n48  = n38 | n46;
  assign n49  = ~n47 & n48;
  assign n50  = n37 & n49;
  assign n51  = n37 | n49;
  assign n52  = ~n50 & n51;
  assign n53  = b_5 & a_3;
  assign n54  = b_4 & a_4;
  assign n55  = a_5 & b_3;
  assign n56  = n54 & n55;
  assign n57  = n54 | n55;
  assign n58  = ~n56 & n57;
  assign n59  = n53 & n58;
  assign n60  = n53 | n58;
  assign n61  = ~n59 & n60;
  assign n62  = b_1 & a_6;
  assign n63  = a_7 & b_0;
  assign n64  = n62 & n63;
  assign n65  = b_2 & a_5;
  assign n66  = n62 | n63;
  assign n67  = ~n64 & n66;
  assign n68  = n65 & n67;
  assign n69  = n64 | n68;
  assign n70  = b_1 & a_7;
  assign n71  = a_6 & b_2;
  assign n72  = n70 | n71;
  assign n73  = b_2 & a_7;
  assign n74  = n62 & n73;
  assign n75  = n72 & ~n74;
  assign n76  = n69 & n75;
  assign n77  = n69 | n75;
  assign n78  = ~n76 & n77;
  assign n79  = n61 & n78;
  assign n80  = n61 | n78;
  assign n81  = ~n79 & n80;
  assign n82  = n65 | n67;
  assign n83  = ~n68 & n82;
  assign n84  = a_5 & b_0;
  assign n85  = n62 & n84;
  assign n86  = a_4 & b_2;
  assign n87  = b_1 & a_5;
  assign n88  = a_6 & b_0;
  assign n89  = n87 | n88;
  assign n90  = ~n85 & n89;
  assign n91  = n86 & n90;
  assign n92  = n85 | n91;
  assign n93  = n83 & n92;
  assign n94  = n43 | n44;
  assign n95  = ~n45 & n94;
  assign n96  = n83 | n92;
  assign n97  = ~n93 & n96;
  assign n98  = n95 & n97;
  assign n99  = n93 | n98;
  assign n100 = n81 & n99;
  assign n101 = n81 | n99;
  assign n102 = ~n100 & n101;
  assign n103 = n52 & n102;
  assign n104 = n52 | n102;
  assign n105 = ~n103 & n104;
  assign n106 = n95 | n97;
  assign n107 = ~n98 & n106;
  assign n108 = n86 | n90;
  assign n109 = ~n91 & n108;
  assign n110 = b_1 & a_4;
  assign n111 = n84 & n110;
  assign n112 = b_2 & a_3;
  assign n113 = n84 | n110;
  assign n114 = ~n111 & n113;
  assign n115 = n112 & n114;
  assign n116 = n111 | n115;
  assign n117 = n109 & n116;
  assign n118 = n26 | n28;
  assign n119 = ~n29 & n118;
  assign n120 = n109 | n116;
  assign n121 = ~n117 & n120;
  assign n122 = n119 & n121;
  assign n123 = n117 | n122;
  assign n124 = n107 & n123;
  assign n125 = n32 | n34;
  assign n126 = ~n35 & n125;
  assign n127 = n107 | n123;
  assign n128 = ~n124 & n127;
  assign n129 = n126 & n128;
  assign n130 = n124 | n129;
  assign n131 = n105 & n130;
  assign n132 = n105 | n130;
  assign n133 = ~n131 & n132;
  assign n134 = n36 & n133;
  assign n135 = n36 | n133;
  assign n136 = ~n134 & n135;
  assign n137 = n126 | n128;
  assign n138 = ~n129 & n137;
  assign n139 = n119 | n121;
  assign n140 = ~n122 & n139;
  assign n141 = n112 | n114;
  assign n142 = ~n115 & n141;
  assign n143 = a_4 & b_0;
  assign n144 = b_1 & a_3;
  assign n145 = n143 & n144;
  assign n146 = a_2 & b_2;
  assign n147 = n143 | n144;
  assign n148 = ~n145 & n147;
  assign n149 = n146 & n148;
  assign n150 = n145 | n149;
  assign n151 = n142 & n150;
  assign n152 = b_5 & a_0;
  assign n153 = b_4 & a_1;
  assign n154 = a_2 & b_3;
  assign n155 = n153 | n154;
  assign n156 = n153 & n154;
  assign n157 = n155 & ~n156;
  assign n158 = n152 & n157;
  assign n159 = n152 | n157;
  assign n160 = ~n158 & n159;
  assign n161 = n142 | n150;
  assign n162 = ~n151 & n161;
  assign n163 = n160 & n162;
  assign n164 = n151 | n163;
  assign n165 = n140 & n164;
  assign n166 = b_6 & a_0;
  assign n167 = n156 | n158;
  assign n168 = n166 & n167;
  assign n169 = n166 | n167;
  assign n170 = ~n168 & n169;
  assign n171 = n140 | n164;
  assign n172 = ~n165 & n171;
  assign n173 = n170 & n172;
  assign n174 = n165 | n173;
  assign n175 = n138 & n174;
  assign n176 = n138 | n174;
  assign n177 = ~n175 & n176;
  assign n178 = n168 & n177;
  assign n179 = n175 | n178;
  assign n180 = n136 | n179;
  assign n181 = n136 & n179;
  assign n182 = n180 & ~n181;
  assign n183 = n168 | n177;
  assign n184 = ~n178 & n183;
  assign n185 = n170 | n172;
  assign n186 = ~n173 & n185;
  assign n187 = n160 | n162;
  assign n188 = ~n163 & n187;
  assign n189 = n146 | n148;
  assign n190 = ~n149 & n189;
  assign n191 = a_2 & b_1;
  assign n192 = b_0 & a_3;
  assign n193 = n191 & n192;
  assign n194 = a_1 & b_2;
  assign n195 = n191 | n192;
  assign n196 = ~n193 & n195;
  assign n197 = n194 & n196;
  assign n198 = n193 | n197;
  assign n199 = n190 & n198;
  assign n200 = a_1 & b_3;
  assign n201 = b_4 & a_0;
  assign n202 = n200 | n201;
  assign n203 = b_3 & a_0;
  assign n204 = n153 & n203;
  assign n205 = n202 & ~n204;
  assign n206 = n190 | n198;
  assign n207 = ~n199 & n206;
  assign n208 = n205 & n207;
  assign n209 = n199 | n208;
  assign n210 = n188 & n209;
  assign n211 = n188 | n209;
  assign n212 = ~n210 & n211;
  assign n213 = n204 & n212;
  assign n214 = n210 | n213;
  assign n215 = n186 & n214;
  assign n216 = n184 & n215;
  assign n217 = n184 | n215;
  assign n218 = ~n216 & n217;
  assign n219 = n186 | n214;
  assign n220 = ~n215 & n219;
  assign n221 = n204 | n212;
  assign n222 = ~n213 & n221;
  assign n223 = n205 | n207;
  assign n224 = ~n208 & n223;
  assign n225 = a_1 & b_1;
  assign n226 = a_2 & b_0;
  assign n227 = n225 & n226;
  assign n228 = b_2 & a_0;
  assign n229 = n225 | n226;
  assign n230 = ~n227 & n229;
  assign n231 = n228 & n230;
  assign n232 = n227 | n231;
  assign n233 = n194 | n196;
  assign n234 = ~n197 & n233;
  assign n235 = n232 & n234;
  assign n236 = n232 | n234;
  assign n237 = ~n235 & n236;
  assign n238 = n203 & n237;
  assign n239 = n235 | n238;
  assign n240 = n224 & n239;
  assign n241 = n222 & n240;
  assign n242 = n220 & n241;
  assign n243 = n220 | n241;
  assign n244 = ~n242 & n243;
  assign n245 = n222 | n240;
  assign n246 = ~n241 & n245;
  assign n247 = n224 | n239;
  assign n248 = ~n240 & n247;
  assign n249 = n228 | n230;
  assign n250 = ~n231 & n249;
  assign n251 = n19 & n250;
  assign n252 = n203 | n237;
  assign n253 = ~n238 & n252;
  assign n254 = n251 & n253;
  assign n255 = n248 & n254;
  assign n256 = n246 & n255;
  assign n257 = n244 & n256;
  assign n258 = n242 | n257;
  assign n259 = n218 & n258;
  assign n260 = n216 | n259;
  assign n261 = n182 & n260;
  assign n262 = n182 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n251 | n253;
  assign n265 = ~n254 & n264;
  assign n266 = n246 | n255;
  assign n267 = ~n256 & n266;
  assign n268 = n181 | n261;
  assign n269 = n131 | n134;
  assign n270 = n47 | n50;
  assign n271 = a_2 & b_7;
  assign n272 = b_6 & a_3;
  assign n273 = n56 | n59;
  assign n274 = n272 & n273;
  assign n275 = n272 | n273;
  assign n276 = ~n274 & n275;
  assign n277 = n271 & n276;
  assign n278 = n271 | n276;
  assign n279 = ~n277 & n278;
  assign n280 = a_4 & b_5;
  assign n281 = b_4 & a_5;
  assign n282 = a_6 & b_3;
  assign n283 = n281 | n282;
  assign n284 = b_4 & a_6;
  assign n285 = n55 & n284;
  assign n286 = n283 & ~n285;
  assign n287 = n280 & n286;
  assign n288 = n280 | n286;
  assign n289 = ~n287 & n288;
  assign n290 = ~n62 & n73;
  assign n291 = n289 & n290;
  assign n292 = n289 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = n76 | n79;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n279 & n297;
  assign n299 = n279 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = n100 | n103;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n270 & n304;
  assign n306 = n270 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = n269 & n307;
  assign n309 = n269 | n307;
  assign n310 = ~n308 & n309;
  assign n311 = n268 | n310;
  assign n312 = n268 & n310;
  assign n313 = n311 & ~n312;
  assign n314 = n19 | n250;
  assign n315 = ~n251 & n314;
  assign n316 = n285 | n287;
  assign n317 = a_4 & b_6;
  assign n318 = n316 & n317;
  assign n319 = b_7 & a_3;
  assign n320 = n316 | n317;
  assign n321 = ~n318 & n320;
  assign n322 = n319 & n321;
  assign n323 = n318 | n322;
  assign n324 = a_7 & b_5;
  assign n325 = n284 & n324;
  assign n326 = b_4 & a_7;
  assign n327 = a_6 & b_5;
  assign n328 = n326 | n327;
  assign n329 = ~n325 & n328;
  assign n330 = b_7 & a_4;
  assign n331 = n282 & n326;
  assign n332 = a_5 & b_5;
  assign n333 = a_7 & b_3;
  assign n334 = n284 | n333;
  assign n335 = ~n331 & n334;
  assign n336 = n332 & n335;
  assign n337 = n331 | n336;
  assign n338 = a_5 & b_6;
  assign n339 = n337 & n338;
  assign n340 = n337 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = n330 & n341;
  assign n343 = n330 | n341;
  assign n344 = ~n342 & n343;
  assign n345 = n329 & n344;
  assign n346 = n329 | n344;
  assign n347 = ~n345 & n346;
  assign n348 = n74 | n291;
  assign n349 = n332 | n335;
  assign n350 = ~n336 & n349;
  assign n351 = n348 & n350;
  assign n352 = n348 | n350;
  assign n353 = ~n351 & n352;
  assign n354 = n319 | n321;
  assign n355 = ~n322 & n354;
  assign n356 = n353 & n355;
  assign n357 = n351 | n356;
  assign n358 = n347 & n357;
  assign n359 = n347 | n357;
  assign n360 = ~n358 & n359;
  assign n361 = n323 & n360;
  assign n362 = n323 | n360;
  assign n363 = ~n361 & n362;
  assign n364 = n295 | n298;
  assign n365 = n353 | n355;
  assign n366 = ~n356 & n365;
  assign n367 = n364 & n366;
  assign n368 = n274 | n277;
  assign n369 = n364 | n366;
  assign n370 = ~n367 & n369;
  assign n371 = n368 & n370;
  assign n372 = n367 | n371;
  assign n373 = n363 & n372;
  assign n374 = n363 | n372;
  assign n375 = ~n373 & n374;
  assign n376 = n302 | n305;
  assign n377 = n368 | n370;
  assign n378 = ~n371 & n377;
  assign n379 = n376 & n378;
  assign n380 = n268 | n308;
  assign n381 = n309 & n380;
  assign n382 = n376 | n378;
  assign n383 = ~n379 & n382;
  assign n384 = n381 & n383;
  assign n385 = n379 | n384;
  assign n386 = n375 | n385;
  assign n387 = n375 & n385;
  assign n388 = n386 & ~n387;
  assign n389 = a_6 & b_6;
  assign n390 = b_7 & a_7;
  assign n391 = n389 & n390;
  assign n392 = ~n389 & n390;
  assign n393 = a_7 & b_6;
  assign n394 = b_7 & a_6;
  assign n395 = n393 | n394;
  assign n396 = ~n391 & n395;
  assign n397 = b_7 & a_5;
  assign n398 = b_6 & n325;
  assign n399 = n325 | n389;
  assign n400 = ~n398 & n399;
  assign n401 = n397 & n400;
  assign n402 = n397 | n400;
  assign n403 = ~n401 & n402;
  assign n404 = n324 & n403;
  assign n405 = n396 & n404;
  assign n406 = n398 | n401;
  assign n407 = n396 | n404;
  assign n408 = ~n405 & n407;
  assign n409 = n406 & n408;
  assign n410 = n405 | n409;
  assign n411 = n392 & n410;
  assign n412 = n391 | n411;
  assign n413 = n392 | n410;
  assign n414 = ~n411 & n413;
  assign n415 = n406 | n408;
  assign n416 = ~n409 & n415;
  assign n417 = n324 | n403;
  assign n418 = ~n404 & n417;
  assign n419 = n345 & n418;
  assign n420 = n339 | n342;
  assign n421 = n345 | n418;
  assign n422 = ~n419 & n421;
  assign n423 = n420 & n422;
  assign n424 = n419 | n423;
  assign n425 = n416 & n424;
  assign n426 = n416 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n420 | n422;
  assign n429 = ~n423 & n428;
  assign n430 = n358 | n361;
  assign n431 = n429 & n430;
  assign n432 = n429 | n430;
  assign n433 = ~n431 & n432;
  assign n434 = n373 | n387;
  assign n435 = n433 & n434;
  assign n436 = n431 | n435;
  assign n437 = n427 & n436;
  assign n438 = n425 | n437;
  assign n439 = n414 & n438;
  assign n440 = n412 | n439;
  assign n441 = n248 | n254;
  assign n442 = ~n255 & n441;
  assign n443 = n381 | n383;
  assign n444 = ~n384 & n443;
  assign n445 = n414 | n438;
  assign n446 = ~n439 & n445;
  assign n447 = n218 | n258;
  assign n448 = ~n259 & n447;
  assign n449 = n427 | n436;
  assign n450 = ~n437 & n449;
  assign n451 = n433 | n434;
  assign n452 = ~n435 & n451;
  assign n453 = n244 | n256;
  assign n454 = ~n257 & n453;
  assign n455 = b_0 & a_0;
  assign s_1  = n21;
  assign s_8  = n263;
  assign s_3  = n265;
  assign s_5  = n267;
  assign s_9  = n313;
  assign s_2  = n315;
  assign s_11 = n388;
  assign s_15 = n440;
  assign s_4  = n442;
  assign s_10 = n444;
  assign s_14 = n446;
  assign s_7  = n448;
  assign s_13 = n450;
  assign s_12 = n452;
  assign s_6  = n454;
  assign s_0  = n455;
endmodule
