module c1355 (G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355);
  input G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9;
  output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;
  wire _w_1994,_w_1992,_w_1991,_w_1989,_w_1986,_w_1981,_w_1980,_w_1975,_w_1973,_w_1972,_w_1970,_w_1964,_w_1962,_w_1960,_w_1959,_w_1958,_w_1957,_w_1954,_w_1952,_w_1946,_w_1940,_w_1971,_w_1939,_w_1936,_w_1934,_w_1933,_w_1956,_w_1929,_w_1925,_w_1924,_w_1923,_w_1921,_w_1919,_w_1917,_w_1916,_w_1915,_w_1913,_w_1909,_w_1908,_w_1904,_w_1903,_w_1902,_w_1899,_w_1984,_w_1888,_w_1886,_w_1883,_w_1880,_w_1879,_w_1877,_w_1875,_w_1874,_w_1872,_w_1920,_w_1870,_w_1869,_w_1867,_w_1865,_w_1862,_w_1861,_w_1859,_w_1858,_w_1856,_w_1852,_w_1851,_w_1850,_w_1849,_w_1846,_w_1845,_w_1841,_w_1840,_w_1839,_w_1838,_w_1836,_w_1887,_w_1829,_w_1828,_w_1827,_w_1826,_w_1825,_w_1823,_w_1820,_w_1819,_w_1818,_w_1816,_w_1811,_w_1810,_w_1808,_w_1804,_w_1835,_w_1803,_w_1800,_w_1799,_w_1795,_w_1794,_w_1792,_w_1791,_w_1790,_w_1789,_w_1911,_w_1786,_w_1785,_w_1873,_w_1853,_w_1784,_w_1783,_w_1782,_w_1781,_w_1778,_w_1777,_w_1776,_w_1772,_w_1770,_w_1768,_w_1766,_w_1763,_w_1762,_w_1760,_w_1759,_w_1758,_w_1756,_w_1876,_w_1755,_w_1747,_w_1963,_w_1745,_w_1743,_w_1731,_w_1727,_w_1938,_w_1726,_w_1725,_w_1720,_w_1719,_w_1718,_w_1717,_w_1716,_w_1812,_w_1712,_w_1711,_w_1707,_w_1706,_w_1704,_w_1703,_w_1700,_w_1698,_w_1966,_w_1697,_w_1696,_w_1694,_w_1691,_w_1690,_w_1687,_w_1686,_w_1685,_w_1680,_w_1676,_w_1674,_w_1673,_w_1670,_w_1668,_w_1666,_w_1665,_w_1657,_w_1655,_w_1654,_w_1653,_w_1652,_w_1650,_w_1649,_w_1647,_w_1639,_w_1637,_w_1634,_w_1633,_w_1630,_w_1626,_w_1624,_w_1623,_w_1621,_w_1618,_w_1614,_w_1612,_w_1627,_w_1610,_w_1607,_w_1606,_w_1605,_w_1604,_w_1603,_w_1601,_w_1599,_w_1597,_w_1595,_w_1592,_w_1590,_w_1589,_w_1976,_w_1588,_w_1927,_w_1587,_w_1582,_w_1581,_w_1580,_w_1837,_w_1576,_w_1575,_w_1574,_w_1572,_w_1570,_w_1567,_w_1645,_w_1563,_w_1561,_w_1559,_w_1558,_w_1557,_w_1556,_w_1552,_w_1551,_w_1550,_w_1543,_w_1542,_w_1541,_w_1539,_w_1538,_w_1555,_w_1537,_w_1535,_w_1534,_w_1544,_w_1533,_w_1530,_w_1529,_w_1524,_w_1831,_w_1522,_w_1520,_w_1519,_w_1518,_w_1798,_w_1516,_w_1513,_w_1511,_w_1507,_w_1505,_w_1504,_w_1503,_w_1502,_w_1501,_w_1692,_w_1500,_w_1495,_w_1494,_w_1761,_w_1493,_w_1492,_w_1491,_w_1490,_w_1489,_w_1488,_w_1806,_w_1486,_w_1482,_w_1481,_w_1809,_w_1479,_w_1478,_w_1476,_w_1474,_w_1471,_w_1470,_w_1469,_w_1467,_w_1461,_w_1458,_w_1456,_w_1455,_w_1451,_w_1448,_w_1444,_w_1855,_w_1443,_w_1440,_w_1439,_w_1648,_w_1438,_w_1434,_w_1433,_w_1431,_w_1427,_w_1425,_w_1424,_w_1421,_w_1496,_w_1420,_w_1656,_w_1419,_w_1416,_w_1415,_w_1414,_w_1754,_w_1732,_w_1437,_w_1412,_w_1868,_w_1410,_w_1407,_w_1406,_w_1405,_w_1402,_w_1400,_w_1399,_w_1395,_w_1394,_w_1393,_w_1616,_w_1392,_w_1995,_w_1515,_w_1391,_w_1390,_w_1389,_w_1387,_w_1974,_w_1386,_w_1383,_w_1547,_w_1381,_w_1379,_w_1377,_w_1678,_w_1376,_w_1373,_w_1371,_w_1705,_w_1454,_w_1370,_w_1369,_w_1713,_w_1368,_w_1367,_w_1947,_w_1366,_w_1365,_w_1364,_w_1363,_w_1950,_w_1362,_w_1361,_w_1360,_w_1358,_w_1356,_w_1355,_w_1677,_w_1353,_w_1350,_w_1348,_w_1736,_w_1347,_w_1346,_w_1345,_w_1343,_w_1342,_w_1430,_w_1339,_w_1807,_w_1337,_w_1336,_w_1335,_w_1598,_w_1344,_w_1333,_w_1332,_w_1330,_w_1699,_w_1329,_w_1327,_w_1325,_w_1324,_w_1321,_w_1320,_w_1319,_w_1318,_w_1317,_w_1937,_w_1315,_w_1312,_w_1310,_w_1305,_w_1303,_w_1301,_w_1300,_w_1299,_w_1297,_w_1296,_w_1295,_w_1689,_w_1294,_w_1293,_w_1292,_w_1290,_w_1288,_w_1546,_w_1287,_w_1521,_w_1286,_w_1283,_w_1282,_w_1955,_w_1280,_w_1277,_w_1276,_w_1275,_w_1272,_w_1485,_w_1270,_w_1708,_w_1269,_w_1468,_w_1267,_w_1264,_w_1263,_w_1748,_w_1262,_w_1261,_w_1259,_w_1688,_w_1257,_w_1256,_w_1255,_w_1254,_w_1253,_w_1459,_w_1251,_w_1250,_w_1248,_w_1244,_w_1242,_w_1241,_w_1240,_w_1237,_w_1487,_w_1236,_w_1235,_w_1596,_w_1233,_w_1232,_w_1231,_w_1230,_w_1228,_w_1224,_w_1222,_w_1428,_w_1221,_w_1409,_w_1243,_w_1220,_w_1480,_w_1217,_w_1900,_w_1735,_w_1215,_w_1214,_w_1212,_w_1211,_w_1210,_w_1209,_w_1208,_w_1206,_w_1204,_w_1734,_w_1352,_w_1202,_w_1200,_w_1197,_w_1196,_w_1585,_w_1194,_w_1191,_w_1190,_w_1817,_w_1187,_w_1186,_w_1185,_w_1432,_w_1184,_w_1219,_w_1183,_w_1632,_w_1181,_w_1180,_w_1179,_w_1176,_w_1174,_w_1173,_w_1171,_w_1170,_w_1168,_w_1664,_w_1166,_w_1751,_w_1165,_w_1396,_w_1163,_w_1161,_w_1160,_w_1159,_w_1483,_w_1158,_w_1157,_w_1156,_w_1246,_w_1155,_w_1152,_w_1949,_w_1150,_w_1617,_w_1146,_w_1144,_w_1140,_w_1139,_w_1138,_w_1137,_w_1134,_w_1132,_w_1131,_w_1129,_w_1127,_w_1126,_w_1125,_w_1124,_w_1123,_w_1121,_w_1120,_w_1117,_w_1216,_w_1115,_w_1114,_w_1112,_w_1111,_w_1110,_w_1663,_w_1109,n249_9,n249_4,G16_0,n249_3,_w_1848,n249_6,n42,G23_1,n251_0,_w_1928,_w_1730,_w_1193,n185_0,n266_1,n144,n269_1,n96,_w_1864,_w_1151,n272_10,n272_6,n272_4,n48_0,n272_3,n272_2,_w_1814,_w_1658,n257_1,_w_1805,n427,_w_1757,G26_7,_w_1285,n279_1,n279_0,_w_1660,_w_1912,n281_3,_w_1843,n294_1,_w_1961,_w_1435,_w_1113,n316_2,_w_1832,_w_1638,n399,n318_3,_w_1894,_w_1475,_w_1417,n318_0,n336_1,n336_0,_w_1354,n249_8,n337_1,n337_0,n345_1,n272_7,n366_0,n370_0,_w_1797,n152_3,_w_1442,n379_2,_w_1833,_w_1584,_w_1068,G5_0,n112_1,n379_0,_w_1943,n232,_w_1988,n405_1,_w_1644,G18_6,n429,n134_0,n49,n425,_w_1942,_w_1473,n304_1,n61,n411,n409,G17_7,_w_1930,_w_1628,_w_1465,n405,n172_7,n397,n362_1,n386,n381,_w_1662,_w_1273,n380,n97_0,n78,_w_1266,n255,n374,n100,n379,G18_7,n237_1,n370,n367,_w_1693,_w_1560,_w_1527,n366,n345,_w_1910,_w_1201,n250_0,n363,n138,_w_1545,n360,n196_0,n359,n207,n424,n91_1,n357,n356,n355,n248,n376,_w_1830,n81_0,n143,G17_6,_w_1130,n346,n343,n121_0,_w_1854,n166_1,_w_1147,n191_3,n420,n212,n338,n272_1,n337,G12_7,_w_1460,n336,n332,n281_2,n146,_w_1302,G30_0,n152_0,n260_0,n316_1,_w_1095,n328,_w_1096,n327,n402,n100_3,n208,n257_0,_w_1323,n416,_w_1622,n393,G15_6,_w_1177,G5_3,n320,_w_1066,_w_1506,n318,n358,G23_0,_w_1154,n310,n239,_w_1188,_w_1092,n306,n304,n199,n300,n252_1,_w_1779,G41_8,_w_1813,_w_1540,_w_1309,n372,_w_1635,n296,n371,n292,n215,_w_1229,G1_6,n284,n397_1,n153_3,n72_1,n269_0,n283,n268,n282,n359_3,n318_1,n324,n351,G17_4,n281,n392_1,G24_2,_w_1723,n302,n279,n182,_w_1701,G26_2,G20_7,n278,n233,n327_0,n272_11,_w_1148,n276,_w_1477,n407,_w_1549,n274,_w_1341,n273,n229_6,_w_1885,n415_0,n272,n191_7,n55,n397_0,n269,n137_1,n251_1,_w_1714,n266,n421,n265,G28_1,G20_5,_w_1108,n317,n124_2,n262,_w_1834,n259,n160_1,_w_1226,n258,n257,n403,_w_1905,n250,G26_5,_w_1891,n114,_w_1278,_w_1172,_w_1071,_w_1671,n300_0,_w_1554,n246,_w_1331,n202_2,n378,_w_1462,n245,n238,n217_1,G32_2,n342,_w_1822,n235,_w_1398,G27_2,n103,_w_1967,n172_5,n236,G23_5,G17_5,n231,n240_1,n359_2,_w_1523,n230,n190,n375,n227,n417,n153,n274_0,n84_0,_w_1374,_w_1931,n186,n93,n163_0,n89,n87,_w_1384,n85,n161,_w_1328,n240,n84,_w_1133,n60_0,n401_0,_w_1351,G14_6,_w_1340,_w_1249,n152_6,_w_1577,n228,n80,_w_1162,n281_1,n414,_w_1357,G19_6,n298,n109,_w_1593,G2_2,n156,_w_1824,n347,_w_1602,n173_1,n68,_w_1907,n65,n64,_w_1213,n45_0,_w_1145,n361,n147,n145,_w_1884,n313,n51_0,_w_1105,n294,n218,n60,n146_1,G30_6,_w_1695,n59,_w_1801,G26_0,n299,_w_1304,n211,n88_0,n58,_w_1586,n263_0,n56,G5_6,_w_1463,G21_3,n73,n427_1,n157_1,n53,_w_1225,n249_5,n122,n260,_w_1090,n264,_w_1968,n152_8,n272_5,n45,n329,G11_5,n312,_w_1764,n47,n74,_w_1239,n370_1,n251,n71,_w_1260,n305,G31_0,_w_1382,n54,n195,G11_7,n261,n51_2,n70,G17_2,n191,n229_8,n288,n158,_w_1667,_w_1422,n282_0,n272_0,n72,_w_1388,_w_1892,n183,G3_6,_w_1724,n323_1,G31_2,_w_1195,n79,n414_1,n107,n160,_w_1738,n410,n54_1,n308_1,G4_4,_w_1897,n364,n366_1,_w_1418,n124,_w_1769,n197,n94,n117,n81,_w_1951,G14_7,n252_0,G12_6,G9_3,n325,G5_4,n69,_w_1227,n231_0,G13_3,n281_0,_w_1118,n45_1,n237_0,n119,G12_0,_w_1613,G13_5,n392,_w_1889,n165,_w_1844,n100_2,n109_1,_w_1629,n277,n76,_w_1314,n48,n282_1,n409_0,_w_1821,_w_1453,n77,n280_1,n134_1,_w_1525,n210,n199_0,n57,n132,n196,_w_1568,n82,n396_0,_w_1948,n272_9,n90,_w_1722,_w_1898,G17_3,n243_0,n97_1,n286,_w_1896,_w_1192,n113,n106,_w_1895,G10_7,n75,n172,n360_1,_w_1088,n205,n131_1,n280,n67,G28_6,n83,n279_2,_w_1636,_w_1252,n249_1,n111,n128_0,_w_1528,G13_7,_w_1932,n91,n341,n98,G32_6,n193_0,n301,n66_0,G5_2,G22_7,n202_3,n249,n321,G12_1,n396_3,_w_1646,_w_1149,n389,_w_1548,n409_1,_w_1093,n423_1,n243_1,G3_0,_w_1372,_w_1223,n379_1,n406,_w_1436,n52,_w_1401,n254_0,n428,_w_1737,G15_5,n423,n384_1,_w_1744,n115_0,G7_3,n50,G31_1,_w_1793,n345_0,G5_1,G32_5,_w_1306,n208_1,n388_1,_w_1532,n115_3,_w_1978,_w_1746,n222,n200,_w_1965,n203,_w_1289,n66_1,_w_1615,_w_1107,n99,_w_1135,n139,n211_0,n318_2,n101,n105,n163,_w_1484,n405_0,G2_4,_w_1796,_w_1274,n390,n223,n118_0,n187,n112,_w_1573,n294_0,n242,n221,G28_7,n243,n359_0,_w_1578,n349,n360_0,G27_6,n154,n178,_w_1446,n246_1,_w_1709,_w_1271,n384_0,n78_3,_w_1787,n120,n123,n126,n127,_w_1234,n256,n172_6,_w_1099,n198,n362,n241,_w_1205,_w_1198,n128,n125,_w_1085,n44,n129,n130,n175,n224,_w_1510,n336_2,n172_0,n271,n133,G21_6,n134,_w_1452,n75_0,n208_0,n135,n118,n136,n216,_w_1609,G18_5,n385,n316_3,_w_1514,n267,_w_1265,n204,_w_1728,n137,n226_1,G1_2,_w_1413,n141,_w_1742,n249_0,_w_1098,_w_1815,_w_1403,_w_1207,n419,_w_1517,_w_1408,n63,n150,n226,n234_1,n191_2,n362_0,_w_1182,G29_3,n384,n151,G24_0,n280_0,n110,n333,_w_1397,G11_4,n152,n249_2,G19_2,n217_0,_w_1702,_w_1279,n152_7,n180,n155,_w_1122,n414_0,G25_7,n157,_w_1741,n184,n396,_w_1385,n193,n75_1,n159,n179_1,_w_1326,_w_1189,n185,G27_5,n162,n60_1,G26_1,_w_1914,_w_1863,n380_0,_w_1969,n194,_w_1316,n327_1,n164,n166,_w_1775,_w_1313,n354,n171,n312_0,n176_1,_w_1426,n177,_w_1457,n368,n179,_w_1641,n349_1,n353,_w_1178,n181,n300_1,_w_1983,n188,n339,n413,G2_6,_w_1944,n189,n201,_w_1375,n246_0,n374_0,n148,n137_2,_w_1102,n314,n97,n66,n78_1,n115,G29_1,_w_1659,n142,G1_3,n209,n88,n213,G41_7,n230_1,n174,n78_4,n217,n219,n172_8,n220,_w_1128,n295,n106_0,n225,n299_0,_w_1531,n234_0,n231_1,n230_0,_w_1116,G28_2,_w_1566,n131,n229_1,n229_2,_w_1378,n414_3,n229_3,_w_1977,n229_5,n229_7,_w_1164,n323,G23_6,n226_0,_w_1579,n319_0,n263_1,n319_1,_w_1411,G8_1,_w_1175,G8_2,_w_1536,G8_3,G8_4,n272_12,n88_1,_w_1359,n149,G8_6,G3_7,G8_7,n206,_w_1094,_w_1979,n87_0,n87_1,_w_1788,_w_1143,n87_2,n388_0,n240_0,_w_1640,_w_1512,n84_1,G15_1,_w_1075,G15_2,n168,G3_1,G15_3,G15_7,n163_1,n414_2,G16_1,n78_0,n350,n124_0,_w_1860,n78_2,G16_6,G2_7,n78_6,n78_7,n361_0,n361_1,n361_2,n361_3,G20_6,n173_0,n299_1,_w_1611,n115_4,n394,n299_3,_w_1918,n290,G16_7,_w_1631,_w_1142,_w_1078,_w_1077,n103_1,n125_0,n214_2,_w_1247,n125_1,_w_1625,n380_1,n140_1,_w_1945,n94_1,G27_0,G29_7,n182_1,n57_1,_w_1423,n286_1,n331_0,n51_1,_w_1322,n51_3,_w_1081,n54_0,_w_1941,G19_0,G19_1,_w_1953,n63_0,G19_5,_w_1167,n188_1,G19_7,n312_1,G2_3,_w_1672,n249_7,n308_0,n191_0,n191_1,n229_0,n191_5,n191_6,n116,n191_8,n323_0,n72_0,_w_1715,_w_1070,n160_0,_w_1682,_w_1084,_w_1338,n140,G7_0,_w_1893,_w_1733,G7_1,n69_1,n103_0,G7_2,G7_4,n396_2,G7_5,n244,G16_5,G7_7,n128_1,G5_5,n247,G14_0,G5_7,G24_6,G41_1,n309,G41_2,n274_1,G41_3,_w_1203,G26_4,_w_1311,G14_2,_w_1773,_w_1729,n109_0,G41_5,G41_6,_w_1683,_w_1526,G9_6,G9_0,_w_1881,G15_4,G41_9,_w_1583,n359_1,G6_0,n316_0,n401,G17_1,G6_1,G19_4,G6_2,_w_1562,G4_6,_w_1749,G6_4,n170,G6_5,G6_6,_w_1404,n223_0,n108,G6_7,_w_1447,G26_6,_w_1565,n124_3,n81_1,n279_3,G32_0,_w_1104,G11_0,G32_1,G28_3,_w_1334,G32_3,_w_1291,n331_1,G32_4,_w_1906,G31_3,G31_4,_w_1600,_w_1466,G31_5,_w_1153,G31_6,_w_1752,n423_0,n298_0,n427_0,G9_1,n298_2,n298_3,G30_1,G4_3,n229_4,n62,G30_2,G30_3,G30_4,G30_5,G14_3,n260_1,G30_7,_w_1449,n287,_w_1065,n392_0,_w_1268,n214,G3_3,n299_2,n102,G3_4,G27_1,n104,G27_3,_w_1882,n341_1,G27_4,_w_1238,G13_0,n401_1,G21_1,n115_1,n229,G27_7,n316,G28_0,G28_4,G28_5,n331,n290_1,n48_1,_w_1740,_w_1079,n63_3,G26_3,G6_3,n176_0,n57_0,_w_1985,n275,G25_0,G25_1,n185_1,G25_2,G25_3,G24_3,G25_4,G25_5,_w_1987,G25_6,G24_1,_w_1871,G24_4,G24_5,n286_0,n51,G10_0,G32_7,n172_1,_w_1441,n172_3,n115_7,n205_0,_w_1847,_w_1258,n43,G18_1,n205_1,n272_8,G31_7,G23_2,_w_1619,_w_1281,n374_1,G23_3,_w_1669,G19_3,n169_1,G23_4,_w_1802,G22_4,G23_7,n169_0,_w_1661,_w_1429,_w_1298,n349_0,n192_1,n91_0,_w_1982,n341_0,_w_1681,G1_4,n290_0,_w_1643,G29_0,G3_5,G29_2,G22_3,_w_1771,G29_4,_w_1721,G9_4,_w_1564,_w_1380,G13_6,n250_1,n291,n86,G29_5,_w_1710,G29_6,_w_1842,G8_0,n182_0,n335,G22_0,n192,G22_1,_w_1499,G22_2,n379_3,n308,n46,G22_5,G22_6,G21_0,n169,n298_1,G4_5,G21_2,_w_1445,G8_5,G7_6,G21_7,n304_0,G20_0,n254,n382,G20_1,_w_1569,G20_2,_w_1497,G20_3,_w_1774,G20_4,_w_1308,G2_0,G2_1,G2_5,n140_0,n270,G18_0,_w_1750,n266_0,G18_3,G18_4,G17_0,_w_1684,n143_0,_w_1087,G16_2,G16_3,G16_4,_w_1620,G9_2,n112_0,_w_1890,_w_1141,G9_5,G15_0,G9_7,_w_1901,_w_1767,_w_1509,_w_1169,G11_1,n419_1,G11_2,_w_1765,n94_0,n191_4,G11_3,n152_5,G11_6,_w_1753,_w_1119,G10_1,_w_1651,G10_2,_w_1866,_w_1608,G10_3,G4_7,G10_4,G10_5,G10_6,n252,G1_0,_w_1591,_w_1508,n202,G41_4,G1_1,n176,G21_4,G1_5,G1_7,n106_1,_w_1594,_w_1245,n87_3,n100_0,_w_1675,n124_1,G21_5,n100_1,n172_4,n199_1,n42_0,_w_1464,n42_1,_w_1076,n223_1,G4_2,_w_1199,n154_0,n154_1,G4_0,G4_1,G41_0,n121_1,n146_0,_w_1307,n196_1,G13_1,G13_2,_w_1993,G13_4,_w_1990,n263,G14_1,G14_4,n336_3,G14_5,n118_1,n172_2,n188_0,n137_0,_w_1935,n137_3,n419_0,_w_1922,_w_1878,_w_1136,G18_2,n254_1,n63_1,_w_1450,n253,n63_2,n202_0,_w_1571,n202_1,n237,n149_0,_w_1739,n149_1,n152_1,n173,n131_0,n152_2,_w_1069,n152_4,n153_0,_w_1349,_w_1284,n153_1,_w_1101,_w_1472,n153_2,G12_2,n167,G12_3,G12_4,G12_5,G3_2,n157_0,n396_1,n193_1,n415_1,n143_1,_w_1780,n388,n214_0,n214_1,n78_5,n214_3,n166_0,n92,n179_0,n192_0,_w_1642,G24_7,n115_2,n115_5,n234,n115_6,_w_1553,n415,n115_8,n319,n220_0,n220_1,_w_1679,_w_1067,_w_1072,_w_1926,_w_1073,n69_0,_w_1074,_w_1080,_w_1857,_w_1082,_w_1218,_w_1083,n95,n398,_w_1086,_w_1089,n78_8,_w_1091,n121,_w_1097,n211_1,_w_1100,_w_1498,_w_1103,_w_1106;

  bfr _b_1574(.a(_w_1995),.q(_w_1994));
  bfr _b_1573(.a(G40),.q(_w_1995));
  bfr _b_1572(.a(_w_1993),.q(_w_1992));
  bfr _b_1568(.a(_w_1989),.q(_w_1988));
  bfr _b_1566(.a(_w_1987),.q(_w_1986));
  bfr _b_1565(.a(G36),.q(_w_1987));
  bfr _b_1563(.a(_w_1984),.q(_w_1983));
  bfr _b_1562(.a(G34),.q(_w_1984));
  bfr _b_1560(.a(_w_1981),.q(n172_2));
  bfr _b_1559(.a(_w_1980),.q(G24_5));
  bfr _b_1556(.a(_w_1977),.q(_w_1978));
  bfr _b_1555(.a(_w_1976),.q(_w_1977));
  bfr _b_1554(.a(_w_1975),.q(_w_1976));
  bfr _b_1553(.a(_w_1974),.q(_w_1975));
  bfr _b_1551(.a(_w_1972),.q(_w_1973));
  bfr _b_1550(.a(_w_1971),.q(_w_1972));
  bfr _b_1546(.a(_w_1967),.q(_w_1968));
  bfr _b_1544(.a(_w_1965),.q(_w_1966));
  bfr _b_1542(.a(_w_1963),.q(_w_1964));
  bfr _b_1539(.a(_w_1960),.q(_w_1961));
  bfr _b_1537(.a(_w_1958),.q(_w_1959));
  bfr _b_1536(.a(_w_1957),.q(G26_5));
  bfr _b_1535(.a(_w_1956),.q(_w_1957));
  bfr _b_1534(.a(_w_1955),.q(_w_1956));
  bfr _b_1533(.a(_w_1954),.q(_w_1955));
  bfr _b_1541(.a(_w_1962),.q(_w_1963));
  bfr _b_1528(.a(_w_1949),.q(_w_1950));
  bfr _b_1526(.a(_w_1947),.q(_w_1948));
  bfr _b_1524(.a(_w_1945),.q(_w_1946));
  bfr _b_1523(.a(_w_1944),.q(_w_1945));
  bfr _b_1522(.a(_w_1943),.q(_w_1944));
  bfr _b_1521(.a(_w_1942),.q(_w_1943));
  bfr _b_1520(.a(_w_1941),.q(_w_1942));
  bfr _b_1519(.a(_w_1940),.q(_w_1941));
  bfr _b_1516(.a(_w_1937),.q(_w_1938));
  bfr _b_1515(.a(_w_1936),.q(_w_1937));
  bfr _b_1513(.a(_w_1934),.q(G27_5));
  bfr _b_1512(.a(_w_1933),.q(_w_1934));
  bfr _b_1510(.a(_w_1931),.q(_w_1932));
  bfr _b_1509(.a(_w_1930),.q(_w_1931));
  bfr _b_1507(.a(_w_1928),.q(_w_1929));
  bfr _b_1506(.a(_w_1927),.q(_w_1928));
  bfr _b_1504(.a(_w_1925),.q(_w_1926));
  bfr _b_1503(.a(_w_1924),.q(_w_1925));
  bfr _b_1502(.a(_w_1923),.q(_w_1924));
  bfr _b_1500(.a(_w_1921),.q(_w_1922));
  bfr _b_1499(.a(_w_1920),.q(_w_1921));
  bfr _b_1497(.a(_w_1918),.q(_w_1919));
  bfr _b_1496(.a(_w_1917),.q(_w_1918));
  bfr _b_1493(.a(_w_1914),.q(_w_1915));
  bfr _b_1491(.a(_w_1912),.q(_w_1913));
  bfr _b_1489(.a(_w_1910),.q(_w_1911));
  bfr _b_1480(.a(_w_1901),.q(_w_1902));
  bfr _b_1479(.a(_w_1900),.q(_w_1901));
  bfr _b_1475(.a(_w_1896),.q(_w_1897));
  bfr _b_1474(.a(_w_1895),.q(_w_1896));
  bfr _b_1473(.a(_w_1894),.q(_w_1895));
  bfr _b_1472(.a(_w_1893),.q(_w_1894));
  bfr _b_1470(.a(_w_1891),.q(_w_1892));
  bfr _b_1468(.a(_w_1889),.q(_w_1890));
  bfr _b_1467(.a(_w_1888),.q(_w_1889));
  bfr _b_1466(.a(_w_1887),.q(n115_2));
  bfr _b_1465(.a(_w_1886),.q(n298_1));
  bfr _b_1463(.a(_w_1884),.q(_w_1885));
  bfr _b_1462(.a(_w_1883),.q(_w_1884));
  bfr _b_1459(.a(_w_1880),.q(_w_1881));
  bfr _b_1458(.a(_w_1879),.q(_w_1880));
  bfr _b_1456(.a(_w_1877),.q(_w_1878));
  bfr _b_1455(.a(_w_1876),.q(_w_1877));
  bfr _b_1454(.a(_w_1875),.q(_w_1876));
  bfr _b_1453(.a(_w_1874),.q(_w_1875));
  bfr _b_1450(.a(_w_1871),.q(_w_1872));
  bfr _b_1449(.a(_w_1870),.q(_w_1871));
  bfr _b_1444(.a(_w_1865),.q(_w_1866));
  bfr _b_1461(.a(_w_1882),.q(G7_5));
  bfr _b_1441(.a(_w_1862),.q(_w_1863));
  bfr _b_1440(.a(_w_1861),.q(_w_1862));
  bfr _b_1431(.a(_w_1852),.q(_w_1853));
  bfr _b_1429(.a(_w_1850),.q(_w_1851));
  bfr _b_1427(.a(_w_1848),.q(G8_5));
  bfr _b_1426(.a(_w_1847),.q(_w_1848));
  bfr _b_1548(.a(_w_1969),.q(_w_1970));
  bfr _b_1424(.a(_w_1845),.q(_w_1846));
  bfr _b_1422(.a(_w_1843),.q(_w_1844));
  bfr _b_1420(.a(_w_1841),.q(_w_1842));
  bfr _b_1419(.a(_w_1840),.q(_w_1841));
  bfr _b_1418(.a(_w_1839),.q(_w_1840));
  bfr _b_1417(.a(_w_1838),.q(_w_1839));
  bfr _b_1416(.a(_w_1837),.q(_w_1838));
  bfr _b_1571(.a(G39),.q(_w_1993));
  bfr _b_1412(.a(_w_1833),.q(_w_1834));
  bfr _b_1410(.a(_w_1831),.q(_w_1832));
  bfr _b_1409(.a(_w_1830),.q(_w_1831));
  bfr _b_1408(.a(_w_1829),.q(_w_1830));
  bfr _b_1407(.a(_w_1828),.q(_w_1829));
  bfr _b_1406(.a(_w_1827),.q(_w_1828));
  bfr _b_1405(.a(_w_1826),.q(_w_1827));
  bfr _b_1404(.a(_w_1825),.q(_w_1826));
  bfr _b_1403(.a(_w_1824),.q(n229_2));
  bfr _b_1402(.a(_w_1823),.q(_w_1824));
  bfr _b_1399(.a(_w_1820),.q(_w_1821));
  bfr _b_1398(.a(_w_1819),.q(_w_1820));
  bfr _b_1396(.a(_w_1817),.q(_w_1818));
  bfr _b_1391(.a(_w_1812),.q(_w_1813));
  bfr _b_1388(.a(_w_1809),.q(_w_1810));
  bfr _b_1387(.a(_w_1808),.q(_w_1809));
  bfr _b_1384(.a(_w_1805),.q(n274_1));
  bfr _b_1381(.a(_w_1802),.q(n316_1));
  bfr _b_1380(.a(_w_1801),.q(_w_1802));
  bfr _b_1378(.a(_w_1799),.q(_w_1800));
  bfr _b_1377(.a(_w_1798),.q(G25_5));
  bfr _b_1413(.a(_w_1834),.q(_w_1835));
  bfr _b_1375(.a(_w_1796),.q(_w_1797));
  bfr _b_1374(.a(_w_1795),.q(_w_1796));
  bfr _b_1371(.a(_w_1792),.q(_w_1793));
  bfr _b_1369(.a(_w_1790),.q(_w_1791));
  bfr _b_1366(.a(_w_1787),.q(_w_1788));
  bfr _b_1364(.a(_w_1785),.q(_w_1786));
  bfr _b_1359(.a(_w_1780),.q(_w_1781));
  bfr _b_1357(.a(_w_1778),.q(_w_1779));
  bfr _b_1356(.a(_w_1777),.q(_w_1778));
  bfr _b_1355(.a(_w_1776),.q(_w_1777));
  bfr _b_1354(.a(_w_1775),.q(G1355));
  bfr _b_1351(.a(_w_1772),.q(_w_1773));
  bfr _b_1350(.a(_w_1771),.q(_w_1772));
  bfr _b_1349(.a(_w_1770),.q(_w_1771));
  bfr _b_1348(.a(_w_1769),.q(_w_1770));
  bfr _b_1347(.a(_w_1768),.q(_w_1769));
  bfr _b_1460(.a(_w_1881),.q(_w_1882));
  bfr _b_1345(.a(_w_1766),.q(_w_1767));
  bfr _b_1341(.a(_w_1762),.q(_w_1763));
  bfr _b_1337(.a(_w_1758),.q(_w_1759));
  bfr _b_1336(.a(_w_1757),.q(_w_1758));
  bfr _b_1335(.a(_w_1756),.q(_w_1757));
  bfr _b_1334(.a(_w_1755),.q(_w_1756));
  bfr _b_1330(.a(_w_1751),.q(_w_1752));
  bfr _b_1329(.a(_w_1750),.q(_w_1751));
  bfr _b_1325(.a(_w_1746),.q(_w_1747));
  bfr _b_1332(.a(_w_1753),.q(_w_1754));
  bfr _b_1322(.a(_w_1743),.q(_w_1744));
  bfr _b_1321(.a(_w_1742),.q(_w_1743));
  bfr _b_1320(.a(_w_1741),.q(_w_1742));
  bfr _b_1525(.a(_w_1946),.q(_w_1947));
  bfr _b_1319(.a(_w_1740),.q(_w_1741));
  bfr _b_1314(.a(_w_1735),.q(_w_1736));
  bfr _b_1312(.a(_w_1733),.q(_w_1734));
  bfr _b_1397(.a(_w_1818),.q(_w_1819));
  bfr _b_1311(.a(_w_1732),.q(_w_1733));
  bfr _b_1307(.a(_w_1728),.q(_w_1729));
  bfr _b_1306(.a(_w_1727),.q(_w_1728));
  bfr _b_1305(.a(_w_1726),.q(_w_1727));
  bfr _b_1303(.a(_w_1724),.q(G1345));
  bfr _b_1302(.a(_w_1723),.q(G1343));
  bfr _b_1301(.a(_w_1722),.q(G1342));
  bfr _b_1300(.a(_w_1721),.q(G1351));
  bfr _b_1298(.a(_w_1719),.q(n272));
  bfr _b_1297(.a(_w_1718),.q(_w_1719));
  bfr _b_1295(.a(_w_1716),.q(_w_1717));
  bfr _b_1294(.a(_w_1715),.q(_w_1716));
  bfr _b_1292(.a(_w_1713),.q(_w_1714));
  bfr _b_1291(.a(_w_1712),.q(_w_1713));
  bfr _b_1290(.a(_w_1711),.q(_w_1712));
  bfr _b_1289(.a(_w_1710),.q(_w_1711));
  bfr _b_1514(.a(_w_1935),.q(_w_1936));
  bfr _b_1287(.a(_w_1708),.q(_w_1709));
  bfr _b_1286(.a(_w_1707),.q(_w_1708));
  bfr _b_1283(.a(_w_1704),.q(_w_1705));
  bfr _b_1282(.a(_w_1703),.q(_w_1704));
  bfr _b_1279(.a(_w_1700),.q(_w_1701));
  bfr _b_1276(.a(_w_1697),.q(_w_1698));
  bfr _b_1275(.a(_w_1696),.q(_w_1697));
  bfr _b_1274(.a(_w_1695),.q(_w_1696));
  bfr _b_1278(.a(_w_1699),.q(_w_1700));
  bfr _b_1272(.a(_w_1693),.q(n316_3));
  bfr _b_1268(.a(_w_1689),.q(G1346));
  bfr _b_1277(.a(_w_1698),.q(_w_1699));
  bfr _b_1267(.a(_w_1688),.q(n250_1));
  bfr _b_1259(.a(_w_1680),.q(_w_1681));
  bfr _b_1254(.a(_w_1675),.q(_w_1676));
  bfr _b_1251(.a(_w_1672),.q(_w_1673));
  bfr _b_1250(.a(_w_1671),.q(_w_1672));
  bfr _b_1249(.a(_w_1670),.q(_w_1671));
  bfr _b_1248(.a(_w_1669),.q(_w_1670));
  bfr _b_1372(.a(_w_1793),.q(_w_1794));
  bfr _b_1246(.a(_w_1667),.q(_w_1668));
  bfr _b_1245(.a(_w_1666),.q(_w_1667));
  bfr _b_1242(.a(_w_1663),.q(_w_1664));
  bfr _b_1241(.a(_w_1662),.q(_w_1663));
  bfr _b_1239(.a(_w_1660),.q(n379));
  bfr _b_1324(.a(_w_1745),.q(_w_1746));
  bfr _b_1235(.a(_w_1656),.q(_w_1657));
  bfr _b_1234(.a(_w_1655),.q(_w_1656));
  bfr _b_1233(.a(_w_1654),.q(_w_1655));
  bfr _b_1361(.a(_w_1782),.q(_w_1783));
  bfr _b_1232(.a(_w_1653),.q(_w_1654));
  bfr _b_1230(.a(_w_1651),.q(_w_1652));
  bfr _b_1229(.a(_w_1650),.q(_w_1651));
  bfr _b_1228(.a(_w_1649),.q(_w_1650));
  bfr _b_1227(.a(_w_1648),.q(n154));
  bfr _b_1224(.a(_w_1645),.q(_w_1646));
  bfr _b_1222(.a(_w_1643),.q(_w_1644));
  bfr _b_1221(.a(_w_1642),.q(_w_1643));
  bfr _b_1270(.a(_w_1691),.q(n336));
  bfr _b_1263(.a(_w_1684),.q(G1344));
  bfr _b_1220(.a(_w_1641),.q(_w_1642));
  bfr _b_1219(.a(_w_1640),.q(_w_1641));
  bfr _b_1443(.a(_w_1864),.q(_w_1865));
  bfr _b_1216(.a(_w_1637),.q(_w_1638));
  bfr _b_1214(.a(_w_1635),.q(_w_1636));
  bfr _b_1213(.a(_w_1634),.q(_w_1635));
  bfr _b_1265(.a(_w_1686),.q(_w_1687));
  bfr _b_1212(.a(_w_1633),.q(_w_1634));
  bfr _b_1211(.a(_w_1632),.q(_w_1633));
  bfr _b_1207(.a(_w_1628),.q(_w_1629));
  bfr _b_1206(.a(_w_1627),.q(_w_1628));
  bfr _b_1204(.a(_w_1625),.q(_w_1626));
  bfr _b_1482(.a(_w_1903),.q(_w_1904));
  bfr _b_1203(.a(_w_1624),.q(_w_1625));
  bfr _b_1201(.a(_w_1622),.q(_w_1623));
  bfr _b_1200(.a(_w_1621),.q(_w_1622));
  bfr _b_1549(.a(_w_1970),.q(_w_1971));
  bfr _b_1199(.a(_w_1620),.q(G1341));
  bfr _b_1198(.a(_w_1619),.q(n254));
  bfr _b_1196(.a(_w_1617),.q(_w_1618));
  bfr _b_1194(.a(_w_1615),.q(_w_1616));
  bfr _b_1193(.a(_w_1614),.q(_w_1615));
  bfr _b_1192(.a(_w_1613),.q(n125));
  bfr _b_1191(.a(_w_1612),.q(_w_1613));
  bfr _b_1190(.a(_w_1611),.q(_w_1612));
  bfr _b_1189(.a(_w_1610),.q(_w_1611));
  bfr _b_1188(.a(_w_1609),.q(G23_5));
  bfr _b_1187(.a(_w_1608),.q(_w_1609));
  bfr _b_1186(.a(_w_1607),.q(_w_1608));
  bfr _b_1389(.a(_w_1810),.q(n272_8));
  bfr _b_1183(.a(_w_1604),.q(_w_1605));
  bfr _b_1180(.a(_w_1601),.q(_w_1602));
  bfr _b_1179(.a(_w_1600),.q(_w_1601));
  bfr _b_1177(.a(_w_1598),.q(_w_1599));
  bfr _b_1176(.a(_w_1597),.q(_w_1598));
  bfr _b_1174(.a(_w_1595),.q(_w_1596));
  bfr _b_1173(.a(_w_1594),.q(_w_1595));
  bfr _b_1171(.a(_w_1592),.q(_w_1593));
  bfr _b_1169(.a(_w_1590),.q(_w_1591));
  bfr _b_1168(.a(_w_1589),.q(_w_1590));
  bfr _b_1167(.a(_w_1588),.q(_w_1589));
  bfr _b_1166(.a(_w_1587),.q(_w_1588));
  bfr _b_1163(.a(_w_1584),.q(_w_1585));
  bfr _b_1162(.a(_w_1583),.q(_w_1584));
  bfr _b_1161(.a(_w_1582),.q(_w_1583));
  bfr _b_1159(.a(_w_1580),.q(_w_1581));
  bfr _b_1158(.a(_w_1579),.q(_w_1580));
  bfr _b_1156(.a(_w_1577),.q(_w_1578));
  bfr _b_1154(.a(_w_1575),.q(_w_1576));
  bfr _b_1153(.a(_w_1574),.q(_w_1575));
  bfr _b_1152(.a(_w_1573),.q(_w_1574));
  bfr _b_1150(.a(_w_1571),.q(_w_1572));
  bfr _b_1148(.a(_w_1569),.q(_w_1570));
  bfr _b_1147(.a(_w_1568),.q(_w_1569));
  bfr _b_1144(.a(_w_1565),.q(_w_1566));
  bfr _b_1142(.a(_w_1563),.q(_w_1564));
  bfr _b_1141(.a(_w_1562),.q(_w_1563));
  bfr _b_1140(.a(_w_1561),.q(n230_1));
  bfr _b_1138(.a(_w_1559),.q(_w_1560));
  bfr _b_1137(.a(_w_1558),.q(_w_1559));
  bfr _b_1136(.a(_w_1557),.q(_w_1558));
  bfr _b_1134(.a(_w_1555),.q(_w_1556));
  bfr _b_1133(.a(_w_1554),.q(n251_1));
  bfr _b_1132(.a(_w_1553),.q(_w_1554));
  bfr _b_1293(.a(_w_1714),.q(_w_1715));
  bfr _b_1131(.a(_w_1552),.q(_w_1553));
  bfr _b_1129(.a(_w_1550),.q(_w_1551));
  bfr _b_1127(.a(_w_1548),.q(_w_1549));
  bfr _b_1126(.a(_w_1547),.q(G1348));
  bfr _b_1125(.a(_w_1546),.q(G18_5));
  bfr _b_1124(.a(_w_1545),.q(_w_1546));
  bfr _b_1160(.a(_w_1581),.q(_w_1582));
  bfr _b_1122(.a(_w_1543),.q(_w_1544));
  bfr _b_1120(.a(_w_1541),.q(_w_1542));
  bfr _b_1119(.a(_w_1540),.q(_w_1541));
  bfr _b_1118(.a(_w_1539),.q(_w_1540));
  bfr _b_1116(.a(_w_1537),.q(_w_1538));
  bfr _b_1115(.a(_w_1536),.q(_w_1537));
  bfr _b_1114(.a(_w_1535),.q(_w_1536));
  bfr _b_1113(.a(_w_1534),.q(_w_1535));
  bfr _b_1111(.a(_w_1532),.q(_w_1533));
  bfr _b_1110(.a(_w_1531),.q(_w_1532));
  bfr _b_1109(.a(_w_1530),.q(_w_1531));
  spl4L g172_s_2(.a(n172_4),.q0(n172_5),.q1(n172_6),.q2(n172_7),.q3(n172_8));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(n140_1));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(n75_1));
  spl3L G24_s_1(.a(G24_2),.q0(G24_3),.q1(G24_4),.q2(_w_1958));
  and_bi g174(.a(n100_2),.b(n173_0),.q(n174));
  bfr _b_1273(.a(_w_1694),.q(_w_1695));
  bfr _b_861(.a(_w_1282),.q(_w_1283));
  spl3L G24_s_0(.a(G24),.q0(G24_0),.q1(G24_1),.q2(G24_2));
  spl3L G25_s_0(.a(G25),.q0(G25_0),.q1(G25_1),.q2(G25_2));
  bfr _b_1486(.a(_w_1907),.q(_w_1908));
  bfr _b_1014(.a(_w_1435),.q(_w_1436));
  bfr _b_1085(.a(_w_1506),.q(_w_1507));
  spl2 G26_s_2(.a(G26_5),.q0(G26_6),.q1(G26_7));
  spl3L G26_s_1(.a(G26_2),.q0(G26_3),.q1(G26_4),.q2(_w_1935));
  bfr _b_665(.a(_w_1086),.q(_w_1087));
  spl2 g388_s_0(.a(n388),.q0(n388_0),.q1(n388_1));
  bfr _b_1471(.a(_w_1892),.q(_w_1893));
  spl3L G28_s_0(.a(G28),.q0(G28_0),.q1(G28_1),.q2(G28_2));
  spl3L G27_s_1(.a(G27_2),.q0(G27_3),.q1(G27_4),.q2(_w_1912));
  spl3L G3_s_1(.a(G3_2),.q0(G3_3),.q1(G3_4),.q2(_w_1888));
  bfr _b_958(.a(_w_1379),.q(_w_1380));
  spl3L G3_s_0(.a(G3),.q0(G3_0),.q1(G3_1),.q2(G3_2));
  spl3L g115_s_0(.a(n115),.q0(n115_0),.q1(n115_1),.q2(_w_1887));
  or_bb g176(.a(n174),.b(n175),.q(n176));
  bfr _b_1098(.a(_w_1519),.q(n229_4));
  bfr _b_1373(.a(_w_1794),.q(_w_1795));
  spl2 g423_s_0(.a(n423),.q0(n423_0),.q1(n423_1));
  bfr _b_1313(.a(_w_1734),.q(_w_1735));
  or_bb g241(.a(n237_0),.b(n240_0),.q(n241));
  spl3L G32_s_0(.a(G32),.q0(G32_0),.q1(G32_1),.q2(G32_2));
  spl3L G20_s_0(.a(G20),.q0(G20_0),.q1(G20_1),.q2(G20_2));
  spl2 G6_s_2(.a(G6_5),.q0(G6_6),.q1(G6_7));
  spl4L G41_s_0(.a(G41),.q0(G41_0),.q1(G41_1),.q2(G41_2),.q3(G41_3));
  spl3L G5_s_0(.a(G5),.q0(G5_0),.q1(G5_1),.q2(G5_2));
  bfr _b_1328(.a(_w_1749),.q(G1352));
  spl3L G7_s_1(.a(G7_2),.q0(G7_3),.q1(G7_4),.q2(_w_1859));
  spl2 g226_s_0(.a(n226),.q0(n226_0),.q1(n226_1));
  bfr _b_860(.a(_w_1281),.q(_w_1282));
  spl2 g160_s_0(.a(n160),.q0(n160_0),.q1(n160_1));
  and_bi g367(.a(G18_6),.b(n366_0),.q(n367));
  spl2 g94_s_0(.a(n94),.q0(n94_0),.q1(n94_1));
  bfr _b_1498(.a(_w_1919),.q(_w_1920));
  or_bb g249(.a(n247),.b(n248),.q(_w_1856));
  and_bb g281(.a(n153_3),.b(n280_0),.q(n281));
  bfr _b_1428(.a(_w_1849),.q(_w_1850));
  bfr _b_1376(.a(_w_1797),.q(_w_1798));
  bfr _b_1039(.a(_w_1460),.q(_w_1461));
  bfr _b_1567(.a(G37),.q(_w_1989));
  spl4L g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1),.q2(n299_2),.q3(n299_3));
  spl4L g78_s_2(.a(n78_4),.q0(n78_5),.q1(n78_6),.q2(n78_7),.q3(n78_8));
  bfr _b_924(.a(_w_1345),.q(_w_1346));
  spl2 g78_s_1(.a(n78_2),.q0(n78_3),.q1(_w_1849));
  and_bi g175(.a(n173_1),.b(n100_3),.q(n175));
  spl4L g414_s_0(.a(n414),.q0(n414_0),.q1(n414_1),.q2(n414_2),.q3(n414_3));
  spl2 g405_s_0(.a(n405),.q0(n405_0),.q1(n405_1));
  and_bb g345(.a(n249_9),.b(n336_2),.q(n345));
  spl3L G15_s_0(.a(G15),.q0(G15_0),.q1(G15_1),.q2(G15_2));
  spl2 g240_s_0(.a(n240),.q0(n240_0),.q1(n240_1));
  spl3L G8_s_1(.a(G8_2),.q0(G8_3),.q1(G8_4),.q2(_w_1825));
  or_bb g342(.a(G14_6),.b(n341_0),.q(n342));
  spl3L g229_s_0(.a(n229),.q0(n229_0),.q1(n229_1),.q2(_w_1822));
  spl4L g249_s_2(.a(n249_5),.q0(n249_6),.q1(n249_7),.q2(n249_8),.q3(n249_9));
  bfr _b_788(.a(_w_1209),.q(_w_1210));
  spl3L g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1),.q2(_w_1858));
  spl2 g249_s_1(.a(n249_3),.q0(n249_4),.q1(_w_1814));
  spl2 g384_s_0(.a(n384),.q0(n384_0),.q1(n384_1));
  bfr _b_993(.a(_w_1414),.q(_w_1415));
  bfr _b_1304(.a(_w_1725),.q(n414));
  spl4L g249_s_0(.a(n249),.q0(n249_0),.q1(n249_1),.q2(n249_2),.q3(n249_3));
  spl2 g252_s_0(.a(n252),.q0(n252_0),.q1(_w_1811));
  spl2 g45_s_0(.a(n45),.q0(n45_0),.q1(n45_1));
  spl4L g318_s_0(.a(n318),.q0(n318_0),.q1(n318_1),.q2(n318_2),.q3(n318_3));
  and_bi g248(.a(n234_1),.b(n246_1),.q(n248));
  bfr _b_1338(.a(_w_1759),.q(_w_1760));
  spl2 g260_s_0(.a(n260),.q0(n260_0),.q1(n260_1));
  spl2 g272_s_1(.a(n272_1),.q0(n272_2),.q1(_w_1806));
  and_bi g291(.a(G3_6),.b(n290_0),.q(n291));
  spl2 g274_s_0(.a(n274),.q0(n274_0),.q1(_w_1803));
  or_bb g237(.a(n235),.b(n236),.q(n237));
  bfr _b_990(.a(_w_1411),.q(_w_1412));
  bfr _b_813(.a(_w_1234),.q(_w_1235));
  spl2 g337_s_0(.a(n337),.q0(n337_0),.q1(n337_1));
  spl2 g323_s_0(.a(n323),.q0(n323_0),.q1(n323_1));
  spl3L G25_s_1(.a(G25_2),.q0(G25_3),.q1(G25_4),.q2(_w_1776));
  bfr _b_1178(.a(_w_1599),.q(_w_1600));
  spl2 g360_s_0(.a(n360),.q0(n360_0),.q1(n360_1));
  spl2 g359_s_1(.a(n359_1),.q0(n359_2),.q1(n359_3));
  bfr _b_1296(.a(_w_1717),.q(G6_5));
  bfr _b_1058(.a(_w_1479),.q(_w_1480));
  spl2 g279_s_0(.a(n279),.q0(n279_0),.q1(n279_1));
  bfr _b_1316(.a(_w_1737),.q(_w_1738));
  and_bb g195(.a(G29_1),.b(G30_1),.q(n195));
  bfr _b_1451(.a(_w_1872),.q(_w_1873));
  bfr _b_1393(.a(_w_1814),.q(_w_1815));
  bfr _b_1343(.a(_w_1764),.q(_w_1765));
  bfr _b_795(.a(_w_1216),.q(_w_1217));
  spl2 G31_s_2(.a(G31_5),.q0(G31_6),.q1(G31_7));
  spl2 g266_s_0(.a(n266),.q0(n266_0),.q1(n266_1));
  spl2 g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1));
  spl2 g380_s_0(.a(n380),.q0(n380_0),.q1(n380_1));
  spl3L G8_s_0(.a(G8),.q0(G8_0),.q1(G8_1),.q2(G8_2));
  or_bi g430(.a(n429),.b(n428),.q(_w_1775));
  and_bb g427(.a(n152_8),.b(n414_3),.q(n427));
  and_bi g425(.a(n423_1),.b(G31_7),.q(n425));
  spl2 g366_s_0(.a(n366),.q0(n366_0),.q1(n366_1));
  and_bi g424(.a(G31_6),.b(n423_0),.q(n424));
  and_bb g429(.a(G32_7),.b(n427_1),.q(n429));
  spl3L G29_s_0(.a(G29),.q0(G29_0),.q1(G29_1),.q2(G29_2));
  spl3L G21_s_0(.a(G21),.q0(G21_0),.q1(G21_1),.q2(G21_2));
  bfr _b_1540(.a(_w_1961),.q(_w_1962));
  bfr _b_681(.a(_w_1102),.q(_w_1103));
  bfr _b_1068(.a(_w_1489),.q(_w_1490));
  and_bi g420(.a(G30_6),.b(n419_0),.q(n420));
  or_bi g418(.a(n417),.b(n416),.q(_w_1749));
  spl2 g282_s_0(.a(n282),.q0(n282_0),.q1(n282_1));
  bfr _b_787(.a(_w_1208),.q(_w_1209));
  bfr _b_1415(.a(_w_1836),.q(_w_1837));
  bfr _b_942(.a(_w_1363),.q(_w_1364));
  spl3L G19_s_1(.a(G19_2),.q0(G19_3),.q1(G19_4),.q2(_w_1726));
  and_bb g415(.a(n172_8),.b(n414_0),.q(n415));
  and_bb g414(.a(n359_3),.b(n413),.q(_w_1725));
  and_bb g413(.a(n250_1),.b(n272_7),.q(n413));
  spl2 G28_s_2(.a(G28_5),.q0(G28_6),.q1(G28_7));
  and_bi g85(.a(n84_0),.b(n81_0),.q(n85));
  or_bb g261(.a(G16_0),.b(G8_0),.q(n261));
  spl3L G22_s_0(.a(G22),.q0(G22_0),.q1(G22_1),.q2(G22_2));
  spl2 G27_s_2(.a(G27_5),.q0(G27_6),.q1(G27_7));
  bfr _b_698(.a(_w_1119),.q(_w_1120));
  bfr _b_1240(.a(_w_1661),.q(_w_1662));
  and_bi g398(.a(G25_6),.b(n397_0),.q(n398));
  and_bb g397(.a(n172_7),.b(n396_0),.q(n397));
  bfr _b_1490(.a(_w_1911),.q(G3_5));
  and_bi g394(.a(n392_1),.b(G24_7),.q(n394));
  and_bb g366(.a(n191_5),.b(n361_1),.q(n366));
  spl2 g118_s_0(.a(n118),.q0(n118_0),.q1(n118_1));
  and_bi g390(.a(n388_1),.b(G23_7),.q(n390));
  or_bb g152(.a(n150),.b(n151),.q(n152));
  and_ii g387(.a(n385),.b(n386),.q(_w_1724));
  bfr _b_1260(.a(_w_1681),.q(_w_1682));
  and_bi g406(.a(G27_6),.b(n405_0),.q(n406));
  bfr _b_691(.a(_w_1112),.q(_w_1113));
  and_ii g377(.a(n375),.b(n376),.q(_w_1723));
  and_bb g374(.a(n152_5),.b(n361_3),.q(n374));
  bfr _b_914(.a(_w_1335),.q(_w_1336));
  spl2 g243_s_0(.a(n243),.q0(n243_0),.q1(n243_1));
  bfr _b_1035(.a(_w_1456),.q(_w_1457));
  and_bi g371(.a(G19_6),.b(n370_0),.q(n371));
  and_bi g61(.a(n60_0),.b(n57_0),.q(n61));
  and_bb g242(.a(n237_1),.b(n240_1),.q(n242));
  bfr _b_957(.a(_w_1378),.q(_w_1379));
  and_bb g370(.a(n115_5),.b(n361_2),.q(n370));
  bfr _b_1033(.a(_w_1454),.q(_w_1455));
  and_bi g368(.a(n366_1),.b(G18_7),.q(n368));
  bfr _b_1342(.a(_w_1763),.q(_w_1764));
  and_ii g365(.a(n363),.b(n364),.q(_w_1720));
  and_bi g364(.a(n362_1),.b(G17_7),.q(n364));
  or_bb g272(.a(n270),.b(n271),.q(_w_1718));
  or_bb g359(.a(n355),.b(n358),.q(n359));
  bfr _b_655(.a(_w_1076),.q(n192_1));
  bfr _b_818(.a(_w_1239),.q(_w_1240));
  bfr _b_1552(.a(_w_1973),.q(_w_1974));
  bfr _b_981(.a(_w_1402),.q(_w_1403));
  bfr _b_1105(.a(_w_1526),.q(_w_1527));
  or_bb g121(.a(n119),.b(n120),.q(n121));
  or_bb g354(.a(n115_3),.b(n152_3),.q(n354));
  and_ii g326(.a(n324),.b(n325),.q(G1333));
  and_bi g283(.a(G1_6),.b(n282_0),.q(n283));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  or_bi g352(.a(n351),.b(n350),.q(G1339));
  spl2 G5_s_2(.a(G5_5),.q0(G5_6),.q1(G5_7));
  and_bb g244(.a(n214_2),.b(n243_0),.q(n244));
  spl2 G13_s_2(.a(G13_5),.q0(G13_6),.q1(G13_7));
  or_bb g350(.a(G16_6),.b(n349_0),.q(n350));
  bfr _b_770(.a(_w_1191),.q(_w_1192));
  bfr _b_940(.a(_w_1361),.q(_w_1362));
  and_bb g349(.a(n272_12),.b(n336_3),.q(n349));
  and_ii g373(.a(n371),.b(n372),.q(_w_1722));
  or_bb g183(.a(n179_0),.b(n182_0),.q(n183));
  spl2 g237_s_0(.a(n237),.q0(n237_0),.q1(n237_1));
  and_bi g347(.a(n345_1),.b(G15_7),.q(n347));
  and_bi g246(.a(n245),.b(n244),.q(n246));
  bfr _b_1121(.a(_w_1542),.q(_w_1543));
  spl2 g176_s_0(.a(n176),.q0(n176_0),.q1(n176_1));
  bfr _b_695(.a(_w_1116),.q(_w_1117));
  and_bb g343(.a(G14_7),.b(n341_1),.q(n343));
  spl4L G41_s_2(.a(G41_3),.q0(G41_6),.q1(G41_7),.q2(G41_8),.q3(G41_9));
  and_bi g255(.a(n63_2),.b(n254_0),.q(n255));
  bfr _b_1425(.a(_w_1846),.q(_w_1847));
  spl2 G25_s_2(.a(G25_5),.q0(G25_6),.q1(G25_7));
  and_bb g339(.a(G13_7),.b(n337_1),.q(n339));
  bfr _b_690(.a(_w_1111),.q(_w_1112));
  or_bb g338(.a(G13_6),.b(n337_0),.q(n338));
  spl4L g229_s_2(.a(n229_4),.q0(n229_5),.q1(n229_6),.q2(n229_7),.q3(n229_8));
  and_bb g336(.a(n279_3),.b(n335),.q(_w_1691));
  and_bb g335(.a(n298_2),.b(n316_2),.q(n335));
  bfr _b_1269(.a(_w_1690),.q(n272_5));
  bfr _b_1087(.a(_w_1508),.q(G30_5));
  bfr _b_1501(.a(_w_1922),.q(_w_1923));
  and_ii g334(.a(n332),.b(n333),.q(G1335));
  and_bi g333(.a(n331_1),.b(G12_7),.q(n333));
  and_bb g184(.a(n179_1),.b(n182_1),.q(n184));
  bfr _b_1040(.a(_w_1461),.q(_w_1462));
  and_bi g332(.a(G12_6),.b(n331_0),.q(n332));
  bfr _b_965(.a(_w_1386),.q(_w_1387));
  or_bb g54(.a(n52),.b(n53),.q(n54));
  bfr _b_1264(.a(_w_1685),.q(G1347));
  spl2 G24_s_2(.a(G24_5),.q0(G24_6),.q1(G24_7));
  spl2 g57_s_0(.a(n57),.q0(n57_0),.q1(n57_1));
  and_ii g330(.a(n328),.b(n329),.q(G1334));
  spl2 G11_s_2(.a(G11_5),.q0(G11_6),.q1(G11_7));
  bfr _b_1210(.a(_w_1631),.q(_w_1632));
  bfr _b_898(.a(_w_1319),.q(_w_1320));
  spl3L G14_s_0(.a(G14),.q0(G14_0),.q1(G14_1),.q2(G14_2));
  and_bi g328(.a(G11_6),.b(n327_0),.q(n328));
  spl3L G19_s_0(.a(G19),.q0(G19_0),.q1(G19_1),.q2(G19_2));
  bfr _b_1243(.a(_w_1664),.q(_w_1665));
  and_bi g324(.a(G10_6),.b(n323_0),.q(n324));
  and_bb g405(.a(n115_7),.b(n396_2),.q(n405));
  and_bi g402(.a(G26_6),.b(n401_0),.q(n402));
  and_bb g56(.a(G22_1),.b(G23_1),.q(n56));
  and_bb g337(.a(n336_0),.b(n78_8),.q(n337));
  bfr _b_1430(.a(_w_1851),.q(_w_1852));
  bfr _b_780(.a(_w_1201),.q(_w_1202));
  and_bb g327(.a(n249_8),.b(n318_2),.q(n327));
  bfr _b_1092(.a(_w_1513),.q(_w_1514));
  bfr _b_1545(.a(_w_1966),.q(_w_1967));
  spl2 g327_s_0(.a(n327),.q0(n327_0),.q1(n327_1));
  spl2 g169_s_0(.a(n169),.q0(n169_0),.q1(n169_1));
  bfr _b_838(.a(_w_1259),.q(_w_1260));
  and_ii g322(.a(n320),.b(n321),.q(G1332));
  spl2 G30_s_2(.a(G30_5),.q0(G30_6),.q1(G30_7));
  and_ii g391(.a(n389),.b(n390),.q(_w_1689));
  bfr _b_1370(.a(_w_1791),.q(_w_1792));
  bfr _b_1323(.a(_w_1744),.q(_w_1745));
  bfr _b_1226(.a(_w_1647),.q(_w_1648));
  spl2 g173_s_0(.a(n173),.q0(n173_0),.q1(n173_1));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(_w_1686));
  and_bi g320(.a(G9_6),.b(n319_0),.q(n320));
  spl4L g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1),.q2(n361_2),.q3(n361_3));
  and_ii g395(.a(n393),.b(n394),.q(_w_1685));
  and_bi g96(.a(G11_4),.b(G9_4),.q(n96));
  bfr _b_1143(.a(_w_1564),.q(_w_1565));
  and_bb g319(.a(n318_0),.b(n78_7),.q(n319));
  spl2 g345_s_0(.a(n345),.q0(n345_0),.q1(n345_1));
  and_bi g314(.a(n312_1),.b(G8_7),.q(n314));
  and_bb g312(.a(n272_10),.b(n299_3),.q(n312));
  bfr _b_1281(.a(_w_1702),.q(_w_1703));
  and_ii g311(.a(n309),.b(n310),.q(G1330));
  and_bi g127(.a(n125_1),.b(n124_1),.q(n127));
  bfr _b_1197(.a(_w_1618),.q(_w_1619));
  bfr _b_985(.a(_w_1406),.q(_w_1407));
  and_bb g362(.a(n172_5),.b(n361_0),.q(n362));
  spl4L g191_s_2(.a(n191_4),.q0(n191_5),.q1(n191_6),.q2(n191_7),.q3(n191_8));
  bfr _b_1481(.a(_w_1902),.q(_w_1903));
  and_bi g263(.a(n261),.b(n262),.q(n263));
  bfr _b_657(.a(_w_1078),.q(_w_1079));
  bfr _b_984(.a(_w_1405),.q(_w_1406));
  and_bb g341(.a(n229_8),.b(n336_1),.q(n341));
  bfr _b_1047(.a(_w_1468),.q(_w_1469));
  and_bi g310(.a(n308_1),.b(G7_7),.q(n310));
  bfr _b_1123(.a(_w_1544),.q(_w_1545));
  and_bi g196(.a(n194),.b(n195),.q(n196));
  or_bb g78(.a(n76),.b(n77),.q(n78));
  and_bi g309(.a(G7_6),.b(n308_0),.q(n309));
  and_ii g307(.a(n305),.b(n306),.q(G1329));
  bfr _b_1395(.a(_w_1816),.q(_w_1817));
  bfr _b_1151(.a(_w_1572),.q(_w_1573));
  bfr _b_1139(.a(_w_1560),.q(_w_1561));
  and_bi g219(.a(G6_1),.b(G10_1),.q(n219));
  spl2 g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1));
  bfr _b_1530(.a(_w_1951),.q(_w_1952));
  bfr _b_1401(.a(_w_1822),.q(_w_1823));
  bfr _b_692(.a(_w_1113),.q(_w_1114));
  bfr _b_1063(.a(_w_1484),.q(_w_1485));
  and_bi g305(.a(G6_6),.b(n304_0),.q(n305));
  bfr _b_1247(.a(_w_1668),.q(_w_1669));
  or_bb g356(.a(n153_0),.b(n298_0),.q(n356));
  and_bb g378(.a(n252_1),.b(n272_6),.q(n378));
  spl2 g84_s_0(.a(n84),.q0(n84_0),.q1(n84_1));
  bfr _b_944(.a(_w_1365),.q(_w_1366));
  bfr _b_970(.a(_w_1391),.q(_w_1392));
  and_ii g383(.a(n381),.b(n382),.q(_w_1684));
  spl2 g146_s_0(.a(n146),.q0(n146_0),.q1(n146_1));
  spl3L G28_s_1(.a(G28_2),.q0(G28_3),.q1(G28_4),.q2(_w_1661));
  and_bb g300(.a(n299_0),.b(n78_6),.q(n300));
  or_bb g92(.a(G10_3),.b(G12_3),.q(n92));
  and_bb g379(.a(n359_2),.b(n378),.q(_w_1660));
  and_bb g299(.a(n280_1),.b(n298_3),.q(n299));
  and_bb g167(.a(n124_2),.b(n166_0),.q(n167));
  and_bb g417(.a(G29_7),.b(n415_1),.q(n417));
  bfr _b_1045(.a(_w_1466),.q(_w_1467));
  and_bb g162(.a(G17_4),.b(G29_4),.q(n162));
  and_bi g158(.a(G21_3),.b(G25_3),.q(n158));
  spl2 g121_s_0(.a(n121),.q0(n121_0),.q1(n121_1));
  bfr _b_797(.a(_w_1218),.q(_w_1219));
  bfr _b_1339(.a(_w_1760),.q(_w_1761));
  and_bi g58(.a(G21_0),.b(G24_0),.q(n58));
  bfr _b_908(.a(_w_1329),.q(_w_1330));
  and_bi g190(.a(n176_1),.b(n188_1),.q(n190));
  bfr _b_1135(.a(_w_1556),.q(_w_1557));
  bfr _b_700(.a(_w_1121),.q(_w_1122));
  bfr _b_1386(.a(_w_1807),.q(_w_1808));
  bfr _b_1244(.a(_w_1665),.q(_w_1666));
  bfr _b_873(.a(_w_1294),.q(_w_1295));
  spl3L G6_s_1(.a(G6_2),.q0(G6_3),.q1(G6_4),.q2(_w_1694));
  spl2 g279_s_1(.a(n279_1),.q0(n279_2),.q1(n279_3));
  and_bi g105(.a(G31_4),.b(G27_4),.q(n105));
  spl4L g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1),.q2(n137_2),.q3(n137_3));
  or_bb g428(.a(G32_6),.b(n427_0),.q(n428));
  and_bb g423(.a(n115_8),.b(n414_2),.q(n423));
  bfr _b_1447(.a(_w_1868),.q(_w_1869));
  bfr _b_1073(.a(_w_1494),.q(_w_1495));
  and_bi g155(.a(n87_2),.b(n154_0),.q(n155));
  spl2 g359_s_0(.a(n359),.q0(n359_0),.q1(n359_1));
  bfr _b_714(.a(_w_1135),.q(_w_1136));
  spl2 g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1));
  bfr _b_703(.a(_w_1124),.q(_w_1125));
  bfr _b_744(.a(_w_1165),.q(_w_1166));
  and_ii g289(.a(n287),.b(n288),.q(G1325));
  bfr _b_1445(.a(_w_1866),.q(_w_1867));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(n88_1));
  bfr _b_814(.a(_w_1235),.q(_w_1236));
  and_bi g421(.a(n419_1),.b(G30_7),.q(n421));
  and_bb g147(.a(n137_0),.b(n146_0),.q(n147));
  and_bi g240(.a(n238),.b(n239),.q(n240));
  bfr _b_1044(.a(_w_1465),.q(_w_1466));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(n112_1));
  bfr _b_1145(.a(_w_1566),.q(_w_1567));
  spl2 g269_s_0(.a(n269),.q0(n269_0),.q1(n269_1));
  and_bi g151(.a(n128_1),.b(n149_1),.q(n151));
  and_bb g318(.a(n316_3),.b(n317),.q(n318));
  bfr _b_880(.a(_w_1301),.q(_w_1302));
  bfr _b_1130(.a(_w_1551),.q(_w_1552));
  bfr _b_890(.a(_w_1311),.q(_w_1312));
  or_bb g144(.a(n140_0),.b(n143_0),.q(n144));
  and_bi g140(.a(n138),.b(n139),.q(n140));
  or_bb g138(.a(G20_3),.b(G24_3),.q(n138));
  and_bi g329(.a(n327_1),.b(G11_7),.q(n329));
  and_bb g88(.a(_w_1992),.b(G41_4),.q(_w_1649));
  or_bb g137(.a(n135),.b(n136),.q(n137));
  and_bb g154(.a(_w_1988),.b(G41_6),.q(_w_1645));
  spl3L G27_s_0(.a(G27),.q0(G27_0),.q1(G27_1),.q2(G27_2));
  or_bb g353(.a(n192_0),.b(n316_0),.q(n353));
  bfr _b_794(.a(_w_1215),.q(_w_1216));
  bfr _b_1028(.a(_w_1449),.q(_w_1450));
  and_bi g200(.a(n199_0),.b(n196_0),.q(n200));
  and_bi g90(.a(n88_1),.b(n87_1),.q(n90));
  and_bi g95(.a(G9_3),.b(G11_3),.q(n95));
  and_bi g209(.a(G26_0),.b(G27_0),.q(n209));
  spl3L G15_s_1(.a(G15_2),.q0(G15_3),.q1(G15_4),.q2(_w_1621));
  or_bb g160(.a(n158),.b(n159),.q(n160));
  and_ii g369(.a(n367),.b(n368),.q(_w_1620));
  spl2 g316_s_0(.a(n316),.q0(n316_0),.q1(_w_1799));
  bfr _b_1106(.a(_w_1527),.q(_w_1528));
  and_bb g254(.a(_w_1986),.b(G41_9),.q(_w_1617));
  spl4L g51_s_0(.a(n51),.q0(n51_0),.q1(n51_1),.q2(n51_2),.q3(n51_3));
  bfr _b_1483(.a(_w_1904),.q(_w_1905));
  bfr _b_737(.a(_w_1158),.q(_w_1159));
  and_bb g130(.a(G14_4),.b(G16_4),.q(n130));
  bfr _b_967(.a(_w_1388),.q(_w_1389));
  or_bb g129(.a(G14_3),.b(G16_3),.q(n129));
  and_bi g53(.a(n42_1),.b(n51_1),.q(n53));
  bfr _b_1117(.a(_w_1538),.q(_w_1539));
  or_bb g187(.a(n137_3),.b(n185_1),.q(n187));
  or_bb g168(.a(n124_3),.b(n166_1),.q(n168));
  and_bi g296(.a(n294_1),.b(G4_7),.q(n296));
  or_bb g128(.a(n126),.b(n127),.q(n128));
  and_bb g193(.a(_w_1983),.b(G41_8),.q(_w_1614));
  bfr _b_926(.a(_w_1347),.q(_w_1348));
  and_bi g126(.a(n124_0),.b(n125_0),.q(n126));
  bfr _b_1531(.a(_w_1952),.q(_w_1953));
  and_bb g125(.a(_w_1994),.b(G41_5),.q(_w_1610));
  bfr _b_696(.a(_w_1117),.q(_w_1118));
  bfr _b_1362(.a(_w_1783),.q(_w_1784));
  bfr _b_1215(.a(_w_1636),.q(_w_1637));
  and_bi g375(.a(G20_6),.b(n374_0),.q(n375));
  or_bb g194(.a(G29_0),.b(G30_0),.q(n194));
  and_bi g123(.a(n118_1),.b(n121_1),.q(n123));
  and_bi g399(.a(n397_1),.b(G25_7),.q(n399));
  bfr _b_1253(.a(_w_1674),.q(_w_1675));
  and_bi g381(.a(G21_6),.b(n380_0),.q(n381));
  and_bi g325(.a(n323_1),.b(G10_7),.q(n325));
  and_bi g119(.a(G6_3),.b(G5_3),.q(n119));
  bfr _b_844(.a(_w_1265),.q(_w_1266));
  bfr _b_1318(.a(_w_1739),.q(_w_1740));
  and_bi g256(.a(n254_1),.b(n63_3),.q(n256));
  and_bi g118(.a(n116),.b(n117),.q(n118));
  and_ii g297(.a(n295),.b(n296),.q(G1327));
  bfr _b_921(.a(_w_1342),.q(_w_1343));
  or_bb g279(.a(n273),.b(n278),.q(n279));
  spl2 g319_s_0(.a(n319),.q0(n319_0),.q1(n319_1));
  spl3L G30_s_0(.a(G30),.q0(G30_0),.q1(G30_1),.q2(G30_2));
  spl2 g312_s_0(.a(n312),.q0(n312_0),.q1(n312_1));
  and_bi g250(.a(n230_0),.b(n249_0),.q(n250));
  bfr _b_853(.a(_w_1274),.q(_w_1275));
  spl3L g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1),.q2(_w_1981));
  spl3L G23_s_1(.a(G23_2),.q0(G23_3),.q1(G23_4),.q2(_w_1587));
  bfr _b_1379(.a(_w_1800),.q(_w_1801));
  spl2 g397_s_0(.a(n397),.q0(n397_0),.q1(n397_1));
  or_bb g225(.a(n214_1),.b(n223_1),.q(n225));
  bfr _b_1056(.a(_w_1477),.q(_w_1478));
  or_bb g234(.a(n232),.b(n233),.q(n234));
  or_bb g111(.a(n100_1),.b(n109_1),.q(n111));
  and_bb g110(.a(n100_0),.b(n109_0),.q(n110));
  and_ii g408(.a(n406),.b(n407),.q(_w_1586));
  and_bb g222(.a(n217_1),.b(n220_1),.q(n222));
  or_bb g220(.a(n218),.b(n219),.q(n220));
  and_bi g150(.a(n149_0),.b(n128_0),.q(n150));
  or_bb g63(.a(n61),.b(n62),.q(n63));
  or_bb g164(.a(n160_0),.b(n163_0),.q(n164));
  and_bi g113(.a(n112_0),.b(n91_0),.q(n113));
  and_bi g201(.a(n196_1),.b(n199_1),.q(n201));
  spl3L G26_s_0(.a(G26),.q0(G26_0),.q1(G26_1),.q2(G26_2));
  bfr _b_821(.a(_w_1242),.q(_w_1243));
  and_bi g306(.a(n304_1),.b(G6_7),.q(n306));
  bfr _b_1439(.a(_w_1860),.q(_w_1861));
  bfr _b_1363(.a(_w_1784),.q(_w_1785));
  bfr _b_1288(.a(_w_1709),.q(_w_1710));
  bfr _b_1091(.a(_w_1512),.q(n78_2));
  and_bb g102(.a(G19_4),.b(G23_4),.q(n102));
  bfr _b_1327(.a(_w_1748),.q(G19_5));
  bfr _b_1280(.a(_w_1701),.q(_w_1702));
  spl2 G2_s_2(.a(G2_5),.q0(G2_6),.q1(G2_7));
  spl2 g257_s_0(.a(n257),.q0(n257_0),.q1(n257_1));
  bfr _b_1042(.a(_w_1463),.q(_w_1464));
  bfr _b_1043(.a(_w_1464),.q(_w_1465));
  and_bi g135(.a(n134_0),.b(n131_0),.q(n135));
  and_bi g66(.a(n64),.b(n65),.q(n66));
  and_bi g389(.a(G23_6),.b(n388_0),.q(n389));
  or_bb g64(.a(G13_0),.b(G5_0),.q(n64));
  and_bi g321(.a(n319_1),.b(G9_7),.q(n321));
  or_bb g161(.a(G17_3),.b(G29_3),.q(n161));
  bfr _b_1484(.a(_w_1905),.q(_w_1906));
  and_bb g294(.a(n272_9),.b(n281_3),.q(n294));
  and_bi g46(.a(G20_0),.b(G18_0),.q(n46));
  and_bi g62(.a(n57_1),.b(n60_1),.q(n62));
  bfr _b_1077(.a(_w_1498),.q(_w_1499));
  spl2 G3_s_2(.a(G3_5),.q0(G3_6),.q1(G3_7));
  spl2 g251_s_0(.a(n251),.q0(n251_0),.q1(_w_1548));
  or_bb g91(.a(n89),.b(n90),.q(n91));
  and_bi g313(.a(G8_6),.b(n312_0),.q(n313));
  and_bi g156(.a(n154_1),.b(n87_3),.q(n156));
  bfr _b_1079(.a(_w_1500),.q(_w_1501));
  and_bi g75(.a(n74),.b(n73),.q(n75));
  spl2 g263_s_0(.a(n263),.q0(n263_0),.q1(n263_1));
  and_bi g217(.a(n215),.b(n216),.q(n217));
  bfr _b_1564(.a(G35),.q(_w_1985));
  bfr _b_1414(.a(_w_1835),.q(_w_1836));
  and_bb g73(.a(n63_0),.b(n72_0),.q(n73));
  and_bi g407(.a(n405_1),.b(G27_7),.q(n407));
  and_bb g108(.a(n103_1),.b(n106_1),.q(n108));
  and_bi g47(.a(G18_1),.b(G20_1),.q(n47));
  and_bi g45(.a(n43),.b(n44),.q(n45));
  bfr _b_875(.a(_w_1296),.q(_w_1297));
  and_bi g197(.a(G32_0),.b(G31_0),.q(n197));
  spl2 G16_s_2(.a(G16_5),.q0(G16_6),.q1(G16_7));
  spl2 g166_s_0(.a(n166),.q0(n166_0),.q1(n166_1));
  bfr _b_1237(.a(_w_1658),.q(_w_1659));
  and_bi g203(.a(n202_0),.b(n193_0),.q(n203));
  bfr _b_713(.a(_w_1134),.q(_w_1135));
  bfr _b_820(.a(_w_1241),.q(_w_1242));
  or_bb g43(.a(G17_0),.b(G19_0),.q(n43));
  and_bi g182(.a(n180),.b(n181),.q(n182));
  or_bb g191(.a(n189),.b(n190),.q(n191));
  bfr _b_1255(.a(_w_1676),.q(_w_1677));
  spl2 G8_s_2(.a(G8_5),.q0(G8_6),.q1(G8_7));
  bfr _b_722(.a(_w_1143),.q(_w_1144));
  bfr _b_831(.a(_w_1252),.q(G9_5));
  bfr _b_867(.a(_w_1288),.q(_w_1289));
  bfr _b_1023(.a(_w_1444),.q(_w_1445));
  and_bi g258(.a(G12_0),.b(G4_0),.q(n258));
  spl2 g81_s_0(.a(n81),.q0(n81_0),.q1(n81_1));
  bfr _b_1435(.a(_w_1856),.q(_w_1857));
  and_bi g133(.a(G15_4),.b(G13_4),.q(n133));
  bfr _b_1057(.a(_w_1478),.q(_w_1479));
  bfr _b_1423(.a(_w_1844),.q(_w_1845));
  and_bb g396(.a(n230_1),.b(n360_1),.q(n396));
  bfr _b_1432(.a(_w_1853),.q(_w_1854));
  and_bi g393(.a(G24_6),.b(n392_0),.q(n393));
  and_bi g269(.a(n268),.b(n267),.q(n269));
  and_bi g287(.a(G2_6),.b(n286_0),.q(n287));
  bfr _b_1266(.a(_w_1687),.q(_w_1688));
  bfr _b_1172(.a(_w_1593),.q(_w_1594));
  and_bi g49(.a(n48_0),.b(n45_0),.q(n49));
  and_bi g376(.a(n374_1),.b(G20_7),.q(n376));
  and_bb g165(.a(n160_1),.b(n163_1),.q(n165));
  bfr _b_999(.a(_w_1420),.q(_w_1421));
  and_bi g302(.a(n300_1),.b(G5_7),.q(n302));
  bfr _b_733(.a(_w_1154),.q(_w_1155));
  and_bi g178(.a(G18_4),.b(G26_4),.q(n178));
  bfr _b_1434(.a(_w_1855),.q(n78_4));
  and_bb g186(.a(n137_2),.b(n185_0),.q(n186));
  bfr _b_1025(.a(_w_1446),.q(_w_1447));
  bfr _b_863(.a(_w_1284),.q(_w_1285));
  bfr _b_726(.a(_w_1147),.q(_w_1148));
  bfr _b_1027(.a(_w_1448),.q(_w_1449));
  and_bi g59(.a(G24_1),.b(G21_1),.q(n59));
  and_bi g141(.a(G32_3),.b(G28_3),.q(n141));
  or_bb g55(.a(G22_0),.b(G23_0),.q(n55));
  bfr _b_1258(.a(_w_1679),.q(_w_1680));
  spl2 g217_s_0(.a(n217),.q0(n217_0),.q1(n217_1));
  or_bb g245(.a(n214_3),.b(n243_1),.q(n245));
  bfr _b_1170(.a(_w_1591),.q(_w_1592));
  and_bb g42(.a(_w_1982),.b(G41_0),.q(_w_1520));
  bfr _b_738(.a(_w_1159),.q(_w_1160));
  and_bi g235(.a(G11_0),.b(G15_0),.q(n235));
  and_bi g149(.a(n148),.b(n147),.q(n149));
  bfr _b_767(.a(_w_1188),.q(_w_1189));
  and_bi g77(.a(n54_1),.b(n75_1),.q(n77));
  bfr _b_1149(.a(_w_1570),.q(_w_1571));
  bfr _b_1086(.a(_w_1507),.q(_w_1508));
  bfr _b_1082(.a(_w_1503),.q(_w_1504));
  bfr _b_1557(.a(_w_1978),.q(_w_1979));
  spl2 g308_s_0(.a(n308),.q0(n308_0),.q1(n308_1));
  bfr _b_1165(.a(_w_1586),.q(G1350));
  and_bi g218(.a(G10_0),.b(G6_0),.q(n218));
  and_bi g57(.a(n55),.b(n56),.q(n57));
  bfr _b_859(.a(_w_1280),.q(_w_1281));
  and_bi g132(.a(G13_3),.b(G15_3),.q(n132));
  bfr _b_1231(.a(_w_1652),.q(n88));
  bfr _b_647(.a(_w_1068),.q(_w_1069));
  bfr _b_1128(.a(_w_1549),.q(_w_1550));
  spl2 g229_s_1(.a(n229_2),.q0(n229_3),.q1(_w_1513));
  spl3L G31_s_0(.a(G31),.q0(G31_0),.q1(G31_1),.q2(G31_2));
  bfr _b_899(.a(_w_1320),.q(_w_1321));
  or_bb g180(.a(G22_3),.b(G30_3),.q(n180));
  and_bi g83(.a(G2_4),.b(G1_4),.q(n83));
  spl2 g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1));
  spl3L g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1),.q2(_w_1510));
  bfr _b_1476(.a(_w_1897),.q(_w_1898));
  bfr _b_1048(.a(_w_1469),.q(_w_1470));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(n280_1));
  and_ii g404(.a(n402),.b(n403),.q(_w_1509));
  and_bb g308(.a(n249_7),.b(n299_2),.q(n308));
  bfr _b_731(.a(_w_1152),.q(_w_1153));
  and_bi g251(.a(n78_1),.b(n229_1),.q(n251));
  and_bi g112(.a(n111),.b(n110),.q(n112));
  and_bi g270(.a(n269_0),.b(n257_0),.q(n270));
  spl3L G23_s_0(.a(G23),.q0(G23_0),.q1(G23_1),.q2(G23_2));
  and_ii g315(.a(n313),.b(n314),.q(G1331));
  spl2 g230_s_0(.a(n230),.q0(n230_0),.q1(_w_1555));
  and_bi g298(.a(n152_1),.b(n115_1),.q(n298));
  spl3L G30_s_1(.a(G30_2),.q0(G30_3),.q1(G30_4),.q2(_w_1486));
  and_bi g163(.a(n161),.b(n162),.q(n163));
  and_bb g65(.a(G13_1),.b(G5_1),.q(n65));
  and_bi g50(.a(n45_1),.b(n48_1),.q(n50));
  or_bb g84(.a(n82),.b(n83),.q(n84));
  bfr _b_668(.a(_w_1089),.q(_w_1090));
  bfr _b_1529(.a(_w_1950),.q(_w_1951));
  or_bi g340(.a(n339),.b(n338),.q(G1336));
  bfr _b_964(.a(_w_1385),.q(_w_1386));
  or_bb g143(.a(n141),.b(n142),.q(n143));
  bfr _b_1181(.a(_w_1602),.q(_w_1603));
  bfr _b_1103(.a(_w_1524),.q(_w_1525));
  spl2 g125_s_0(.a(n125),.q0(n125_0),.q1(n125_1));
  and_bb g265(.a(n260_1),.b(n263_1),.q(n265));
  and_bb g207(.a(G25_1),.b(G28_1),.q(n207));
  and_bb g360(.a(n274_1),.b(n359_0),.q(n360));
  bfr _b_769(.a(_w_1190),.q(_w_1191));
  bfr _b_1310(.a(_w_1731),.q(_w_1732));
  and_bb g93(.a(G10_4),.b(G12_4),.q(n93));
  and_bi g271(.a(n257_1),.b(n269_1),.q(n271));
  spl2 g143_s_0(.a(n143),.q0(n143_0),.q1(n143_1));
  bfr _b_1457(.a(_w_1878),.q(_w_1879));
  and_bi g122(.a(n121_0),.b(n118_0),.q(n122));
  and_bi g86(.a(n81_1),.b(n84_1),.q(n86));
  spl2 g392_s_0(.a(n392),.q0(n392_0),.q1(n392_1));
  bfr _b_833(.a(_w_1254),.q(_w_1255));
  bfr _b_935(.a(_w_1356),.q(_w_1357));
  bfr _b_742(.a(_w_1163),.q(_w_1164));
  or_bb g134(.a(n132),.b(n133),.q(n134));
  spl2 g72_s_0(.a(n72),.q0(n72_0),.q1(n72_1));
  and_bi g89(.a(n87_0),.b(n88_0),.q(n89));
  bfr _b_652(.a(_w_1073),.q(_w_1074));
  and_bi g52(.a(n51_0),.b(n42_0),.q(n52));
  and_bi g363(.a(G17_6),.b(n362_0),.q(n363));
  and_bi g76(.a(n75_0),.b(n54_0),.q(n76));
  bfr _b_1271(.a(_w_1692),.q(_w_1693));
  or_bb g107(.a(n103_0),.b(n106_0),.q(n107));
  bfr _b_666(.a(_w_1087),.q(_w_1088));
  bfr _b_832(.a(_w_1253),.q(_w_1254));
  spl2 G32_s_2(.a(G32_5),.q0(G32_6),.q1(G32_7));
  spl2 g172_s_1(.a(n172_2),.q0(n172_3),.q1(_w_1653));
  or_bb g100(.a(n98),.b(n99),.q(n100));
  bfr _b_1561(.a(G33),.q(_w_1982));
  bfr _b_730(.a(_w_1151),.q(_w_1152));
  bfr _b_1256(.a(_w_1677),.q(_w_1678));
  bfr _b_765(.a(_w_1186),.q(_w_1187));
  and_bi g103(.a(n101),.b(n102),.q(n103));
  and_bi g72(.a(n70),.b(n71),.q(n72));
  and_bi g99(.a(n94_1),.b(n97_1),.q(n99));
  bfr _b_1052(.a(_w_1473),.q(_w_1474));
  spl2 g286_s_0(.a(n286),.q0(n286_0),.q1(n286_1));
  spl3L G11_s_1(.a(G11_2),.q0(G11_3),.q1(G11_4),.q2(_w_1750));
  and_bi g208(.a(n206),.b(n207),.q(n208));
  spl2 G41_s_1(.a(G41_2),.q0(G41_4),.q1(G41_5));
  and_bi g213(.a(n208_1),.b(n211_1),.q(n213));
  and_bi g169(.a(n168),.b(n167),.q(n169));
  and_bi g170(.a(n169_0),.b(n157_0),.q(n170));
  bfr _b_1218(.a(_w_1639),.q(_w_1640));
  and_bb g290(.a(n249_6),.b(n281_2),.q(n290));
  and_ii g285(.a(n283),.b(n284),.q(G1324));
  bfr _b_1317(.a(_w_1738),.q(_w_1739));
  spl2 g370_s_0(.a(n370),.q0(n370_0),.q1(n370_1));
  and_bi g171(.a(n157_1),.b(n169_1),.q(n171));
  bfr _b_1000(.a(_w_1421),.q(_w_1422));
  spl2 G7_s_2(.a(G7_5),.q0(G7_6),.q1(G7_7));
  spl3L G18_s_1(.a(G18_2),.q0(G18_3),.q1(G18_4),.q2(_w_1524));
  spl2 G15_s_2(.a(G15_5),.q0(G15_6),.q1(G15_7));
  bfr _b_1081(.a(_w_1502),.q(_w_1503));
  bfr _b_1340(.a(_w_1761),.q(_w_1762));
  and_bb g173(.a(_w_1990),.b(G41_7),.q(_w_1459));
  and_ii g426(.a(n424),.b(n425),.q(_w_1458));
  bfr _b_882(.a(_w_1303),.q(_w_1304));
  bfr _b_1257(.a(_w_1678),.q(_w_1679));
  and_bi g252(.a(n251_0),.b(n249_1),.q(n252));
  or_bb g179(.a(n177),.b(n178),.q(n179));
  bfr _b_1344(.a(_w_1765),.q(_w_1766));
  and_bb g317(.a(n153_2),.b(n279_2),.q(n317));
  and_ii g412(.a(n410),.b(n411),.q(_w_1721));
  bfr _b_915(.a(_w_1336),.q(_w_1337));
  and_bi g131(.a(n129),.b(n130),.q(n131));
  and_bb g216(.a(G14_1),.b(G2_1),.q(n216));
  and_bi g228(.a(n205_1),.b(n226_1),.q(n228));
  and_bi g358(.a(n356),.b(n357),.q(n358));
  bfr _b_1157(.a(_w_1578),.q(_w_1579));
  spl2 g246_s_0(.a(n246),.q0(n246_0),.q1(n246_1));
  and_bi g230(.a(n229_0),.b(n78_0),.q(n230));
  bfr _b_707(.a(_w_1128),.q(_w_1129));
  spl2 g103_s_0(.a(n103),.q0(n103_0),.q1(n103_1));
  bfr _b_996(.a(_w_1417),.q(_w_1418));
  and_bi g346(.a(G15_6),.b(n345_0),.q(n346));
  bfr _b_1517(.a(_w_1938),.q(_w_1939));
  or_bb g264(.a(n260_0),.b(n263_0),.q(n264));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(_w_1453));
  and_bi g185(.a(n183),.b(n184),.q(n185));
  and_bi g188(.a(n187),.b(n186),.q(n188));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  and_bi g166(.a(n164),.b(n165),.q(n166));
  and_bb g409(.a(n152_7),.b(n396_3),.q(n409));
  and_bi g273(.a(n253),.b(n272_4),.q(n273));
  bfr _b_1495(.a(_w_1916),.q(_w_1917));
  spl4L g124_s_0(.a(n124),.q0(n124_0),.q1(n124_1),.q2(n124_2),.q3(n124_3));
  or_bb g157(.a(n155),.b(n156),.q(n157));
  and_bb g331(.a(n272_11),.b(n318_3),.q(n331));
  and_bb g380(.a(n172_6),.b(n379_0),.q(n380));
  bfr _b_772(.a(_w_1193),.q(_w_1194));
  or_bb g199(.a(n197),.b(n198),.q(n199));
  and_bi g292(.a(n290_1),.b(G3_7),.q(n292));
  bfr _b_786(.a(_w_1207),.q(_w_1208));
  and_bb g401(.a(n191_7),.b(n396_1),.q(n401));
  and_bb g392(.a(n152_6),.b(n379_3),.q(n392));
  and_bb g117(.a(G7_4),.b(G8_4),.q(n117));
  bfr _b_684(.a(_w_1105),.q(_w_1106));
  bfr _b_912(.a(_w_1333),.q(_w_1334));
  or_bb g202(.a(n200),.b(n201),.q(n202));
  bfr _b_1175(.a(_w_1596),.q(_w_1597));
  bfr _b_660(.a(_w_1081),.q(_w_1082));
  and_bi g226(.a(n225),.b(n224),.q(n226));
  spl2 g362_s_0(.a(n362),.q0(n362_0),.q1(n362_1));
  and_ii g400(.a(n398),.b(n399),.q(_w_1547));
  spl2 g157_s_0(.a(n157),.q0(n157_0),.q1(n157_1));
  and_bi g198(.a(G31_1),.b(G32_1),.q(n198));
  bfr _b_688(.a(_w_1109),.q(_w_1110));
  and_bi g204(.a(n193_1),.b(n202_1),.q(n204));
  bfr _b_760(.a(_w_1181),.q(_w_1182));
  and_bi g372(.a(n370_1),.b(G19_7),.q(n372));
  bfr _b_922(.a(_w_1343),.q(_w_1344));
  bfr _b_928(.a(_w_1349),.q(_w_1350));
  bfr _b_1532(.a(_w_1953),.q(_w_1954));
  bfr _b_1464(.a(_w_1885),.q(_w_1886));
  bfr _b_1309(.a(_w_1730),.q(_w_1731));
  and_bi g82(.a(G1_3),.b(G2_3),.q(n82));
  and_bi g301(.a(G5_6),.b(n300_0),.q(n301));
  bfr _b_943(.a(_w_1364),.q(_w_1365));
  bfr _b_1112(.a(_w_1533),.q(_w_1534));
  or_bb g206(.a(G25_0),.b(G28_0),.q(n206));
  spl2 G23_s_2(.a(G23_5),.q0(G23_6),.q1(G23_7));
  or_bb g106(.a(n104),.b(n105),.q(n106));
  or_bb g115(.a(n113),.b(n114),.q(n115));
  spl2 g272_s_0(.a(n272),.q0(n272_0),.q1(n272_1));
  and_bi g288(.a(n286_1),.b(G2_7),.q(n288));
  bfr _b_1083(.a(_w_1504),.q(_w_1505));
  or_bb g74(.a(n63_1),.b(n72_1),.q(n74));
  and_bi g210(.a(G27_1),.b(G26_1),.q(n210));
  or_bb g253(.a(n250_0),.b(n252_0),.q(n253));
  bfr _b_1433(.a(_w_1854),.q(_w_1855));
  spl2 G19_s_2(.a(G19_5),.q0(G19_6),.q1(G19_7));
  spl2 g211_s_0(.a(n211),.q0(n211_0),.q1(n211_1));
  bfr _b_1358(.a(_w_1779),.q(_w_1780));
  bfr _b_706(.a(_w_1127),.q(_w_1128));
  bfr _b_1543(.a(_w_1964),.q(_w_1965));
  or_bb g70(.a(n66_0),.b(n69_0),.q(n70));
  and_bi g382(.a(n380_1),.b(G21_7),.q(n382));
  bfr _b_1236(.a(_w_1657),.q(_w_1658));
  and_bi g67(.a(G1_0),.b(G9_0),.q(n67));
  or_bb g214(.a(n212),.b(n213),.q(n214));
  bfr _b_1360(.a(_w_1781),.q(_w_1782));
  and_bb g384(.a(n191_6),.b(n379_1),.q(n384));
  bfr _b_858(.a(_w_1279),.q(_w_1280));
  spl3L G32_s_1(.a(G32_2),.q0(G32_3),.q1(G32_4),.q2(_w_1430));
  and_bi g274(.a(n249_2),.b(n272_0),.q(n274));
  spl3L G13_s_0(.a(G13),.q0(G13_0),.q1(G13_1),.q2(G13_2));
  spl4L g87_s_0(.a(n87),.q0(n87_0),.q1(n87_1),.q2(n87_2),.q3(n87_3));
  spl2 g272_s_2(.a(n272_3),.q0(n272_4),.q1(_w_1690));
  or_bb g116(.a(G7_3),.b(G8_3),.q(n116));
  or_bb g215(.a(G14_0),.b(G2_0),.q(n215));
  bfr _b_790(.a(_w_1211),.q(_w_1212));
  or_bb g221(.a(n217_0),.b(n220_0),.q(n221));
  bfr _b_1421(.a(_w_1842),.q(_w_1843));
  bfr _b_1164(.a(_w_1585),.q(G5_5));
  bfr _b_718(.a(_w_1139),.q(_w_1140));
  or_bb g229(.a(n227),.b(n228),.q(n229));
  spl2 g298_s_1(.a(n298_1),.q0(n298_2),.q1(_w_1428));
  and_bi g223(.a(n221),.b(n222),.q(n223));
  bfr _b_829(.a(_w_1250),.q(_w_1251));
  bfr _b_1061(.a(_w_1482),.q(_w_1483));
  or_bb g277(.a(n229_3),.b(n78_3),.q(n277));
  bfr _b_885(.a(_w_1306),.q(_w_1307));
  spl3L G7_s_0(.a(G7),.q0(G7_0),.q1(G7_1),.q2(G7_2));
  and_bb g224(.a(n214_0),.b(n223_0),.q(n224));
  bfr _b_1155(.a(_w_1576),.q(_w_1577));
  and_bi g192(.a(n172_0),.b(n191_0),.q(n192));
  bfr _b_1100(.a(_w_1521),.q(_w_1522));
  and_bi g227(.a(n226_0),.b(n205_0),.q(n227));
  and_bi g247(.a(n246_0),.b(n234_0),.q(n247));
  bfr _b_874(.a(_w_1295),.q(_w_1296));
  spl2 g48_s_0(.a(n48),.q0(n48_0),.q1(n48_1));
  and_bi g259(.a(G4_1),.b(G12_1),.q(n259));
  or_bi g344(.a(n343),.b(n342),.q(G1337));
  spl3L G11_s_0(.a(G11),.q0(G11_0),.q1(G11_1),.q2(G11_2));
  or_bb g238(.a(G3_0),.b(G7_0),.q(n238));
  and_bi g212(.a(n211_0),.b(n208_0),.q(n212));
  spl2 g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1));
  and_bb g231(.a(_w_1985),.b(G41_1),.q(_w_1424));
  spl3L G29_s_1(.a(G29_2),.q0(G29_3),.q1(G29_4),.q2(_w_1463));
  bfr _b_697(.a(_w_1118),.q(_w_1119));
  bfr _b_1024(.a(_w_1445),.q(_w_1446));
  bfr _b_781(.a(_w_1202),.q(_w_1203));
  bfr _b_1067(.a(_w_1488),.q(_w_1489));
  and_bi g232(.a(n51_2),.b(n231_0),.q(n232));
  and_bi g233(.a(n231_1),.b(n51_3),.q(n233));
  spl2 G17_s_2(.a(G17_5),.q0(G17_6),.q1(G17_7));
  and_bb g304(.a(n229_6),.b(n299_1),.q(n304));
  bfr _b_1018(.a(_w_1439),.q(_w_1440));
  and_bi g243(.a(n241),.b(n242),.q(n243));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(n179_1));
  and_bi g177(.a(G26_3),.b(G18_3),.q(n177));
  and_ii g422(.a(n420),.b(n421),.q(_w_1774));
  bfr _b_959(.a(_w_1380),.q(_w_1381));
  spl2 g331_s_0(.a(n331),.q0(n331_0),.q1(n331_1));
  and_bi g410(.a(G28_6),.b(n409_0),.q(n410));
  bfr _b_807(.a(_w_1228),.q(G10_5));
  or_bb g101(.a(G19_3),.b(G23_3),.q(n101));
  or_bb g260(.a(n258),.b(n259),.q(n260));
  and_bb g419(.a(n191_8),.b(n414_1),.q(n419));
  and_bi g120(.a(G5_4),.b(G6_4),.q(n120));
  and_bb g262(.a(G16_1),.b(G8_1),.q(n262));
  or_bb g97(.a(n95),.b(n96),.q(n97));
  bfr _b_656(.a(_w_1077),.q(_w_1078));
  and_bi g236(.a(G15_1),.b(G11_1),.q(n236));
  bfr _b_1527(.a(_w_1948),.q(_w_1949));
  bfr _b_1518(.a(_w_1939),.q(_w_1940));
  and_bb g282(.a(n281_0),.b(n78_5),.q(n282));
  spl3L G31_s_1(.a(G31_2),.q0(G31_3),.q1(G31_4),.q2(_w_1401));
  bfr _b_971(.a(_w_1392),.q(G22_5));
  or_bb g205(.a(n203),.b(n204),.q(n205));
  bfr _b_966(.a(_w_1387),.q(_w_1388));
  or_bb g60(.a(n58),.b(n59),.q(n60));
  and_bb g267(.a(n202_2),.b(n266_0),.q(n267));
  spl4L g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1),.q2(n379_2),.q3(n379_3));
  bfr _b_1508(.a(_w_1929),.q(_w_1930));
  bfr _b_871(.a(_w_1292),.q(_w_1293));
  and_bi g109(.a(n107),.b(n108),.q(n109));
  and_bi g275(.a(n272_2),.b(n249_4),.q(n275));
  bfr _b_1299(.a(_w_1720),.q(G1340));
  bfr _b_1262(.a(_w_1683),.q(G28_5));
  spl2 g153_s_1(.a(n153_1),.q0(n153_2),.q1(_w_1400));
  and_bi g104(.a(G27_3),.b(G31_3),.q(n104));
  bfr _b_646(.a(_w_1067),.q(_w_1068));
  or_bb g276(.a(n274_0),.b(n275),.q(n276));
  and_bi g278(.a(n276),.b(n277),.q(n278));
  spl2 g205_s_0(.a(n205),.q0(n205_0),.q1(n205_1));
  bfr _b_1093(.a(_w_1514),.q(_w_1515));
  and_bb g280(.a(n192_1),.b(n279_0),.q(n280));
  spl2 g191_s_1(.a(n191_2),.q0(n191_3),.q1(_w_1393));
  bfr _b_812(.a(_w_1233),.q(_w_1234));
  or_bb g69(.a(n67),.b(n68),.q(n69));
  and_bb g286(.a(n229_5),.b(n281_1),.q(n286));
  spl2 g298_s_0(.a(n298),.q0(n298_0),.q1(_w_1883));
  and_bb g80(.a(G3_4),.b(G4_4),.q(n80));
  and_bi g295(.a(G4_6),.b(n294_0),.q(n295));
  spl2 g91_s_0(.a(n91),.q0(n91_0),.q1(n91_1));
  bfr _b_1071(.a(_w_1492),.q(_w_1493));
  and_bi g114(.a(n91_1),.b(n112_1),.q(n114));
  spl2 g341_s_0(.a(n341),.q0(n341_0),.q1(n341_1));
  spl4L g202_s_0(.a(n202),.q0(n202_0),.q1(n202_1),.q2(n202_2),.q3(n202_3));
  bfr _b_1352(.a(_w_1773),.q(G11_5));
  spl2 G29_s_2(.a(G29_5),.q0(G29_6),.q1(G29_7));
  spl2 g254_s_0(.a(n254),.q0(n254_0),.q1(n254_1));
  spl2 g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1));
  spl3L G22_s_1(.a(G22_2),.q0(G22_3),.q1(G22_4),.q2(_w_1370));
  bfr _b_916(.a(_w_1337),.q(_w_1338));
  bfr _b_1146(.a(_w_1567),.q(_w_1568));
  spl2 G22_s_2(.a(G22_5),.q0(G22_6),.q1(G22_7));
  spl3L G21_s_1(.a(G21_2),.q0(G21_3),.q1(G21_4),.q2(_w_1347));
  spl2 G21_s_2(.a(G21_5),.q0(G21_6),.q1(G21_7));
  spl3L G20_s_1(.a(G20_2),.q0(G20_3),.q1(G20_4),.q2(_w_1324));
  spl2 G20_s_2(.a(G20_5),.q0(G20_6),.q1(G20_7));
  bfr _b_777(.a(_w_1198),.q(_w_1199));
  spl3L G2_s_0(.a(G2),.q0(G2_0),.q1(G2_1),.q2(G2_2));
  bfr _b_1195(.a(_w_1616),.q(n193));
  and_bi g316(.a(n191_1),.b(n172_1),.q(n316));
  spl3L G2_s_1(.a(G2_2),.q0(G2_3),.q1(G2_4),.q2(_w_1300));
  spl2 g401_s_0(.a(n401),.q0(n401_0),.q1(n401_1));
  bfr _b_694(.a(_w_1115),.q(_w_1116));
  bfr _b_1442(.a(_w_1863),.q(_w_1864));
  spl3L G18_s_0(.a(G18),.q0(G18_0),.q1(G18_1),.q2(G18_2));
  bfr _b_1217(.a(_w_1638),.q(_w_1639));
  and_bb g361(.a(n251_1),.b(n360_0),.q(n361));
  spl2 G18_s_2(.a(G18_5),.q0(G18_6),.q1(G18_7));
  bfr _b_1570(.a(_w_1991),.q(_w_1990));
  bfr _b_1060(.a(_w_1481),.q(_w_1482));
  spl3L G17_s_0(.a(G17),.q0(G17_0),.q1(G17_1),.q2(G17_2));
  spl3L G17_s_1(.a(G17_2),.q0(G17_3),.q1(G17_4),.q2(_w_1277));
  spl3L G16_s_0(.a(G16),.q0(G16_0),.q1(G16_1),.q2(G16_2));
  bfr _b_739(.a(_w_1160),.q(_w_1161));
  spl3L g272_s_3(.a(n272_5),.q0(n272_6),.q1(n272_7),.q2(_w_1807));
  spl3L G16_s_1(.a(G16_2),.q0(G16_3),.q1(G16_4),.q2(_w_1253));
  spl3L G9_s_0(.a(G9),.q0(G9_0),.q1(G9_1),.q2(G9_2));
  spl4L g214_s_0(.a(n214),.q0(n214_0),.q1(n214_1),.q2(n214_2),.q3(n214_3));
  bfr _b_1394(.a(_w_1815),.q(_w_1816));
  spl3L G9_s_1(.a(G9_2),.q0(G9_3),.q1(G9_4),.q2(_w_1229));
  spl2 G9_s_2(.a(G9_5),.q0(G9_6),.q1(G9_7));
  bfr _b_776(.a(_w_1197),.q(_w_1198));
  bfr _b_1016(.a(_w_1437),.q(_w_1438));
  bfr _b_842(.a(_w_1263),.q(_w_1264));
  spl2 g97_s_0(.a(n97),.q0(n97_0),.q1(n97_1));
  spl2 G1_s_2(.a(G1_5),.q0(G1_6),.q1(G1_7));
  spl3L G10_s_0(.a(G10),.q0(G10_0),.q1(G10_1),.q2(G10_2));
  bfr _b_782(.a(_w_1203),.q(_w_1204));
  spl3L G10_s_1(.a(G10_2),.q0(G10_3),.q1(G10_4),.q2(_w_1205));
  bfr _b_951(.a(_w_1372),.q(_w_1373));
  spl2 G10_s_2(.a(G10_5),.q0(G10_6),.q1(G10_7));
  or_bb g268(.a(n202_3),.b(n266_1),.q(n268));
  spl3L G1_s_1(.a(G1_2),.q0(G1_3),.q1(G1_4),.q2(_w_1181));
  spl2 g106_s_0(.a(n106),.q0(n106_0),.q1(n106_1));
  spl2 g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1));
  spl2 g427_s_0(.a(n427),.q0(n427_0),.q1(n427_1));
  spl2 g42_s_0(.a(n42),.q0(n42_0),.q1(n42_1));
  spl2 g154_s_0(.a(n154),.q0(n154_0),.q1(n154_1));
  spl3L G4_s_0(.a(G4),.q0(G4_0),.q1(G4_1),.q2(G4_2));
  and_bi g355(.a(n353),.b(n354),.q(n355));
  spl3L G4_s_1(.a(G4_2),.q0(G4_3),.q1(G4_4),.q2(_w_1157));
  bfr _b_1437(.a(_w_1858),.q(n191_2));
  spl3L g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1),.q2(_w_1156));
  bfr _b_864(.a(_w_1285),.q(_w_1286));
  spl3L G6_s_0(.a(G6),.q0(G6_0),.q1(G6_1),.q2(G6_2));
  bfr _b_693(.a(_w_1114),.q(_w_1115));
  bfr _b_1069(.a(_w_1490),.q(_w_1491));
  spl2 g196_s_0(.a(n196),.q0(n196_0),.q1(n196_1));
  spl2 g131_s_0(.a(n131),.q0(n131_0),.q1(n131_1));
  spl2 g290_s_0(.a(n290),.q0(n290_0),.q1(n290_1));
  bfr _b_824(.a(_w_1245),.q(_w_1246));
  bfr _b_1485(.a(_w_1906),.q(_w_1907));
  spl2 g134_s_0(.a(n134),.q0(n134_0),.q1(n134_1));
  bfr _b_1368(.a(_w_1789),.q(_w_1790));
  bfr _b_658(.a(_w_1079),.q(_w_1080));
  or_bb g211(.a(n209),.b(n210),.q(n211));
  spl3L G13_s_1(.a(G13_2),.q0(G13_3),.q1(G13_4),.q2(_w_1132));
  bfr _b_648(.a(_w_1069),.q(_w_1070));
  or_bb g79(.a(G3_3),.b(G4_3),.q(n79));
  bfr _b_768(.a(_w_1189),.q(_w_1190));
  spl3L G14_s_1(.a(G14_2),.q0(G14_3),.q1(G14_4),.q2(_w_1108));
  bfr _b_995(.a(_w_1416),.q(_w_1417));
  spl2 G14_s_2(.a(G14_5),.q0(G14_6),.q1(G14_7));
  bfr _b_982(.a(_w_1403),.q(_w_1404));
  spl2 g419_s_0(.a(n419),.q0(n419_0),.q1(n419_1));
  spl2 g152_s_1(.a(n152_2),.q0(n152_3),.q1(_w_1101));
  and_bb g388(.a(n115_6),.b(n379_2),.q(n388));
  spl4L g152_s_2(.a(n152_4),.q0(n152_5),.q1(n152_6),.q2(n152_7),.q3(n152_8));
  spl3L G12_s_0(.a(G12),.q0(G12_0),.q1(G12_1),.q2(G12_2));
  spl3L G12_s_1(.a(G12_2),.q0(G12_3),.q1(G12_4),.q2(_w_1077));
  spl2 G4_s_2(.a(G4_5),.q0(G4_6),.q1(G4_7));
  spl2 G12_s_2(.a(G12_5),.q0(G12_6),.q1(G12_7));
  and_bb g71(.a(n66_1),.b(n69_1),.q(n71));
  spl4L g396_s_0(.a(n396),.q0(n396_0),.q1(n396_1),.q2(n396_2),.q3(n396_3));
  bfr _b_1205(.a(_w_1626),.q(_w_1627));
  spl2 g415_s_0(.a(n415),.q0(n415_0),.q1(n415_1));
  bfr _b_1208(.a(_w_1629),.q(_w_1630));
  and_bb g351(.a(G16_7),.b(n349_1),.q(n351));
  bfr _b_835(.a(_w_1256),.q(_w_1257));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  bfr _b_1075(.a(_w_1496),.q(_w_1497));
  spl2 g163_s_0(.a(n163),.q0(n163_0),.q1(n163_1));
  spl2 g192_s_0(.a(n192),.q0(n192_0),.q1(_w_1072));
  spl4L g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1),.q2(n63_2),.q3(n63_3));
  spl2 g115_s_1(.a(n115_2),.q0(n115_3),.q1(_w_1065));
  spl2 g409_s_0(.a(n409),.q0(n409_0),.q1(n409_1));
  and_bi g386(.a(n384_1),.b(G22_7),.q(n386));
  bfr _b_798(.a(_w_1219),.q(_w_1220));
  spl4L g115_s_2(.a(n115_4),.q0(n115_5),.q1(n115_6),.q2(n115_7),.q3(n115_8));
  spl2 g208_s_0(.a(n208),.q0(n208_0),.q1(n208_1));
  spl2 g220_s_0(.a(n220),.q0(n220_0),.q1(n220_1));
  spl2 g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1));
  bfr _b_644(.a(_w_1065),.q(_w_1066));
  bfr _b_1066(.a(_w_1487),.q(_w_1488));
  or_bb g257(.a(n255),.b(n256),.q(n257));
  bfr _b_650(.a(_w_1071),.q(n115_4));
  bfr _b_651(.a(_w_1072),.q(_w_1073));
  bfr _b_653(.a(_w_1074),.q(_w_1075));
  bfr _b_654(.a(_w_1075),.q(_w_1076));
  bfr _b_1477(.a(_w_1898),.q(_w_1899));
  bfr _b_1385(.a(_w_1806),.q(n272_3));
  bfr _b_659(.a(_w_1080),.q(_w_1081));
  bfr _b_662(.a(_w_1083),.q(_w_1084));
  bfr _b_663(.a(_w_1084),.q(_w_1085));
  bfr _b_1446(.a(_w_1867),.q(_w_1868));
  spl4L g272_s_4(.a(n272_8),.q0(n272_9),.q1(n272_10),.q2(n272_11),.q3(n272_12));
  bfr _b_664(.a(_w_1085),.q(_w_1086));
  bfr _b_686(.a(_w_1107),.q(n152_4));
  bfr _b_979(.a(_w_1400),.q(n153_3));
  bfr _b_886(.a(_w_1307),.q(_w_1308));
  bfr _b_1225(.a(_w_1646),.q(_w_1647));
  bfr _b_669(.a(_w_1090),.q(_w_1091));
  bfr _b_1096(.a(_w_1517),.q(_w_1518));
  bfr _b_670(.a(_w_1091),.q(_w_1092));
  bfr _b_1400(.a(_w_1821),.q(n249_5));
  bfr _b_891(.a(_w_1312),.q(_w_1313));
  bfr _b_671(.a(_w_1092),.q(_w_1093));
  bfr _b_729(.a(_w_1150),.q(_w_1151));
  bfr _b_1202(.a(_w_1623),.q(_w_1624));
  or_bb g124(.a(n122),.b(n123),.q(n124));
  bfr _b_672(.a(_w_1093),.q(_w_1094));
  bfr _b_673(.a(_w_1094),.q(_w_1095));
  bfr _b_839(.a(_w_1260),.q(_w_1261));
  bfr _b_675(.a(_w_1096),.q(_w_1097));
  bfr _b_661(.a(_w_1082),.q(_w_1083));
  bfr _b_676(.a(_w_1097),.q(_w_1098));
  bfr _b_678(.a(_w_1099),.q(_w_1100));
  bfr _b_679(.a(_w_1100),.q(G12_5));
  bfr _b_1019(.a(_w_1440),.q(_w_1441));
  or_bb g172(.a(n170),.b(n171),.q(n172));
  or_bb g48(.a(n46),.b(n47),.q(n48));
  bfr _b_938(.a(_w_1359),.q(_w_1360));
  bfr _b_682(.a(_w_1103),.q(_w_1104));
  bfr _b_683(.a(_w_1104),.q(_w_1105));
  bfr _b_1365(.a(_w_1786),.q(_w_1787));
  bfr _b_685(.a(_w_1106),.q(_w_1107));
  bfr _b_1448(.a(_w_1869),.q(_w_1870));
  spl2 g66_s_0(.a(n66),.q0(n66_0),.q1(n66_1));
  bfr _b_766(.a(_w_1187),.q(_w_1188));
  bfr _b_896(.a(_w_1317),.q(_w_1318));
  bfr _b_689(.a(_w_1110),.q(_w_1111));
  bfr _b_699(.a(_w_1120),.q(_w_1121));
  bfr _b_1436(.a(_w_1857),.q(n249));
  and_bi g385(.a(G22_6),.b(n384_0),.q(n385));
  bfr _b_701(.a(_w_1122),.q(_w_1123));
  bfr _b_784(.a(_w_1205),.q(_w_1206));
  bfr _b_702(.a(_w_1123),.q(_w_1124));
  bfr _b_1367(.a(_w_1788),.q(_w_1789));
  bfr _b_704(.a(_w_1125),.q(_w_1126));
  bfr _b_1326(.a(_w_1747),.q(_w_1748));
  bfr _b_1005(.a(_w_1426),.q(_w_1427));
  bfr _b_708(.a(_w_1129),.q(_w_1130));
  bfr _b_893(.a(_w_1314),.q(_w_1315));
  and_ii g303(.a(n301),.b(n302),.q(G1328));
  bfr _b_709(.a(_w_1130),.q(_w_1131));
  bfr _b_710(.a(_w_1131),.q(G14_5));
  bfr _b_711(.a(_w_1132),.q(_w_1133));
  bfr _b_1488(.a(_w_1909),.q(_w_1910));
  bfr _b_1333(.a(_w_1754),.q(_w_1755));
  bfr _b_712(.a(_w_1133),.q(_w_1134));
  bfr _b_715(.a(_w_1136),.q(_w_1137));
  bfr _b_919(.a(_w_1340),.q(_w_1341));
  bfr _b_716(.a(_w_1137),.q(_w_1138));
  or_bb g148(.a(n137_1),.b(n146_1),.q(n148));
  bfr _b_720(.a(_w_1141),.q(_w_1142));
  spl4L g336_s_0(.a(n336),.q0(n336_0),.q1(n336_1),.q2(n336_2),.q3(n336_3));
  bfr _b_721(.a(_w_1142),.q(_w_1143));
  bfr _b_1049(.a(_w_1470),.q(_w_1471));
  bfr _b_1008(.a(_w_1429),.q(n298_3));
  bfr _b_723(.a(_w_1144),.q(_w_1145));
  bfr _b_724(.a(_w_1145),.q(_w_1146));
  bfr _b_1054(.a(_w_1475),.q(_w_1476));
  and_bi g159(.a(G25_4),.b(G21_4),.q(n159));
  bfr _b_1022(.a(_w_1443),.q(_w_1444));
  bfr _b_725(.a(_w_1146),.q(_w_1147));
  bfr _b_1494(.a(_w_1915),.q(_w_1916));
  bfr _b_1238(.a(_w_1659),.q(n172_4));
  bfr _b_727(.a(_w_1148),.q(_w_1149));
  bfr _b_1390(.a(_w_1811),.q(_w_1812));
  bfr _b_728(.a(_w_1149),.q(_w_1150));
  bfr _b_734(.a(_w_1155),.q(G13_5));
  bfr _b_884(.a(_w_1305),.q(_w_1306));
  and_bi g189(.a(n188_0),.b(n176_0),.q(n189));
  bfr _b_677(.a(_w_1098),.q(_w_1099));
  bfr _b_735(.a(_w_1156),.q(n152_2));
  bfr _b_740(.a(_w_1161),.q(_w_1162));
  bfr _b_1097(.a(_w_1518),.q(_w_1519));
  bfr _b_783(.a(_w_1204),.q(G1_5));
  bfr _b_732(.a(_w_1153),.q(_w_1154));
  bfr _b_743(.a(_w_1164),.q(_w_1165));
  and_bi g136(.a(n131_1),.b(n134_1),.q(n136));
  bfr _b_808(.a(_w_1229),.q(_w_1230));
  bfr _b_745(.a(_w_1166),.q(_w_1167));
  bfr _b_746(.a(_w_1167),.q(_w_1168));
  bfr _b_1569(.a(G38),.q(_w_1991));
  bfr _b_747(.a(_w_1168),.q(_w_1169));
  and_ii g348(.a(n346),.b(n347),.q(G1338));
  and_bi g153(.a(n115_0),.b(n152_0),.q(n153));
  bfr _b_876(.a(_w_1297),.q(_w_1298));
  bfr _b_748(.a(_w_1169),.q(_w_1170));
  bfr _b_749(.a(_w_1170),.q(_w_1171));
  bfr _b_939(.a(_w_1360),.q(_w_1361));
  bfr _b_750(.a(_w_1171),.q(_w_1172));
  and_bi g146(.a(n144),.b(n145),.q(n146));
  bfr _b_751(.a(_w_1172),.q(_w_1173));
  bfr _b_785(.a(_w_1206),.q(_w_1207));
  spl4L g100_s_0(.a(n100),.q0(n100_0),.q1(n100_1),.q2(n100_2),.q3(n100_3));
  bfr _b_815(.a(_w_1236),.q(_w_1237));
  bfr _b_1055(.a(_w_1476),.q(_w_1477));
  bfr _b_752(.a(_w_1173),.q(_w_1174));
  bfr _b_753(.a(_w_1174),.q(_w_1175));
  bfr _b_779(.a(_w_1200),.q(_w_1201));
  spl2 g223_s_0(.a(n223),.q0(n223_0),.q1(n223_1));
  bfr _b_754(.a(_w_1175),.q(_w_1176));
  bfr _b_755(.a(_w_1176),.q(_w_1177));
  bfr _b_756(.a(_w_1177),.q(_w_1178));
  bfr _b_757(.a(_w_1178),.q(_w_1179));
  bfr _b_927(.a(_w_1348),.q(_w_1349));
  bfr _b_758(.a(_w_1179),.q(_w_1180));
  or_bb g357(.a(n172_3),.b(n191_3),.q(n357));
  bfr _b_759(.a(_w_1180),.q(G4_5));
  spl2 g54_s_0(.a(n54),.q0(n54_0),.q1(n54_1));
  bfr _b_762(.a(_w_1183),.q(_w_1184));
  bfr _b_763(.a(_w_1184),.q(_w_1185));
  and_bi g142(.a(G28_4),.b(G32_4),.q(n142));
  bfr _b_764(.a(_w_1185),.q(_w_1186));
  bfr _b_792(.a(_w_1213),.q(_w_1214));
  bfr _b_771(.a(_w_1192),.q(_w_1193));
  bfr _b_1102(.a(_w_1523),.q(n42));
  bfr _b_773(.a(_w_1194),.q(_w_1195));
  bfr _b_817(.a(_w_1238),.q(_w_1239));
  bfr _b_1009(.a(_w_1430),.q(_w_1431));
  and_bb g145(.a(n140_1),.b(n143_1),.q(n145));
  bfr _b_774(.a(_w_1195),.q(_w_1196));
  bfr _b_775(.a(_w_1196),.q(_w_1197));
  bfr _b_852(.a(_w_1273),.q(_w_1274));
  bfr _b_1547(.a(_w_1968),.q(_w_1969));
  bfr _b_778(.a(_w_1199),.q(_w_1200));
  and_bi g403(.a(n401_1),.b(G26_7),.q(n403));
  bfr _b_789(.a(_w_1210),.q(_w_1211));
  bfr _b_791(.a(_w_1212),.q(_w_1213));
  bfr _b_793(.a(_w_1214),.q(_w_1215));
  bfr _b_796(.a(_w_1217),.q(_w_1218));
  bfr _b_799(.a(_w_1220),.q(_w_1221));
  bfr _b_1505(.a(_w_1926),.q(_w_1927));
  bfr _b_947(.a(_w_1368),.q(_w_1369));
  bfr _b_977(.a(_w_1398),.q(_w_1399));
  bfr _b_801(.a(_w_1222),.q(_w_1223));
  bfr _b_802(.a(_w_1223),.q(_w_1224));
  bfr _b_952(.a(_w_1373),.q(_w_1374));
  bfr _b_803(.a(_w_1224),.q(_w_1225));
  bfr _b_804(.a(_w_1225),.q(_w_1226));
  bfr _b_806(.a(_w_1227),.q(_w_1228));
  bfr _b_809(.a(_w_1230),.q(_w_1231));
  bfr _b_1308(.a(_w_1729),.q(_w_1730));
  bfr _b_810(.a(_w_1231),.q(_w_1232));
  bfr _b_811(.a(_w_1232),.q(_w_1233));
  bfr _b_826(.a(_w_1247),.q(_w_1248));
  bfr _b_830(.a(_w_1251),.q(_w_1252));
  bfr _b_953(.a(_w_1374),.q(_w_1375));
  bfr _b_1511(.a(_w_1932),.q(_w_1933));
  bfr _b_816(.a(_w_1237),.q(_w_1238));
  bfr _b_900(.a(_w_1321),.q(_w_1322));
  bfr _b_1095(.a(_w_1516),.q(_w_1517));
  bfr _b_819(.a(_w_1240),.q(_w_1241));
  bfr _b_823(.a(_w_1244),.q(_w_1245));
  and_bi g411(.a(n409_1),.b(G28_7),.q(n411));
  bfr _b_825(.a(_w_1246),.q(_w_1247));
  bfr _b_827(.a(_w_1248),.q(_w_1249));
  bfr _b_649(.a(_w_1070),.q(_w_1071));
  spl2 g234_s_0(.a(n234),.q0(n234_0),.q1(n234_1));
  and_bi g98(.a(n97_0),.b(n94_0),.q(n98));
  bfr _b_828(.a(_w_1249),.q(_w_1250));
  bfr _b_674(.a(_w_1095),.q(_w_1096));
  bfr _b_834(.a(_w_1255),.q(_w_1256));
  bfr _b_836(.a(_w_1257),.q(_w_1258));
  bfr _b_837(.a(_w_1258),.q(_w_1259));
  bfr _b_846(.a(_w_1267),.q(_w_1268));
  bfr _b_968(.a(_w_1389),.q(_w_1390));
  bfr _b_991(.a(_w_1412),.q(_w_1413));
  bfr _b_840(.a(_w_1261),.q(_w_1262));
  bfr _b_841(.a(_w_1262),.q(_w_1263));
  bfr _b_1411(.a(_w_1832),.q(_w_1833));
  bfr _b_843(.a(_w_1264),.q(_w_1265));
  bfr _b_845(.a(_w_1266),.q(_w_1267));
  and_bb g181(.a(G22_4),.b(G30_4),.q(n181));
  bfr _b_645(.a(_w_1066),.q(_w_1067));
  bfr _b_667(.a(_w_1088),.q(_w_1089));
  bfr _b_847(.a(_w_1268),.q(_w_1269));
  bfr _b_850(.a(_w_1271),.q(_w_1272));
  spl3L G1_s_0(.a(G1),.q0(G1_0),.q1(G1_1),.q2(G1_2));
  bfr _b_851(.a(_w_1272),.q(_w_1273));
  bfr _b_1041(.a(_w_1462),.q(n173));
  bfr _b_854(.a(_w_1275),.q(_w_1276));
  and_bi g68(.a(G9_1),.b(G1_1),.q(n68));
  bfr _b_855(.a(_w_1276),.q(G16_5));
  bfr _b_849(.a(_w_1270),.q(_w_1271));
  bfr _b_856(.a(_w_1277),.q(_w_1278));
  bfr _b_1029(.a(_w_1450),.q(_w_1451));
  bfr _b_857(.a(_w_1278),.q(_w_1279));
  bfr _b_862(.a(_w_1283),.q(_w_1284));
  bfr _b_865(.a(_w_1286),.q(_w_1287));
  bfr _b_866(.a(_w_1287),.q(_w_1288));
  bfr _b_1538(.a(_w_1959),.q(_w_1960));
  bfr _b_868(.a(_w_1289),.q(_w_1290));
  and_ii g293(.a(n291),.b(n292),.q(G1326));
  or_bb g51(.a(n49),.b(n50),.q(n51));
  bfr _b_869(.a(_w_1290),.q(_w_1291));
  bfr _b_870(.a(_w_1291),.q(_w_1292));
  bfr _b_1261(.a(_w_1682),.q(_w_1683));
  bfr _b_872(.a(_w_1293),.q(_w_1294));
  bfr _b_1478(.a(_w_1899),.q(_w_1900));
  bfr _b_877(.a(_w_1298),.q(_w_1299));
  bfr _b_719(.a(_w_1140),.q(_w_1141));
  bfr _b_878(.a(_w_1299),.q(G17_5));
  bfr _b_879(.a(_w_1300),.q(_w_1301));
  bfr _b_883(.a(_w_1304),.q(_w_1305));
  bfr _b_887(.a(_w_1308),.q(_w_1309));
  bfr _b_888(.a(_w_1309),.q(_w_1310));
  bfr _b_1031(.a(_w_1452),.q(G32_5));
  bfr _b_909(.a(_w_1330),.q(_w_1331));
  bfr _b_889(.a(_w_1310),.q(_w_1311));
  bfr _b_1383(.a(_w_1804),.q(_w_1805));
  or_bb g416(.a(G29_6),.b(n415_0),.q(n416));
  spl3L G5_s_1(.a(G5_2),.q0(G5_3),.q1(G5_4),.q2(_w_1562));
  or_bb g87(.a(n85),.b(n86),.q(n87));
  bfr _b_892(.a(_w_1313),.q(_w_1314));
  bfr _b_925(.a(_w_1346),.q(G20_5));
  bfr _b_1003(.a(_w_1424),.q(_w_1425));
  bfr _b_894(.a(_w_1315),.q(_w_1316));
  bfr _b_1469(.a(_w_1890),.q(_w_1891));
  bfr _b_705(.a(_w_1126),.q(_w_1127));
  bfr _b_895(.a(_w_1316),.q(_w_1317));
  bfr _b_897(.a(_w_1318),.q(_w_1319));
  bfr _b_901(.a(_w_1322),.q(_w_1323));
  bfr _b_1315(.a(_w_1736),.q(_w_1737));
  bfr _b_902(.a(_w_1323),.q(G2_5));
  and_bi g81(.a(n79),.b(n80),.q(n81));
  bfr _b_903(.a(_w_1324),.q(_w_1325));
  bfr _b_904(.a(_w_1325),.q(_w_1326));
  bfr _b_905(.a(_w_1326),.q(_w_1327));
  bfr _b_1346(.a(_w_1767),.q(_w_1768));
  bfr _b_906(.a(_w_1327),.q(_w_1328));
  spl2 g193_s_0(.a(n193),.q0(n193_0),.q1(n193_1));
  spl2 g60_s_0(.a(n60),.q0(n60_0),.q1(n60_1));
  spl2 g349_s_0(.a(n349),.q0(n349_0),.q1(n349_1));
  bfr _b_907(.a(_w_1328),.q(_w_1329));
  spl4L g281_s_0(.a(n281),.q0(n281_0),.q1(n281_1),.q2(n281_2),.q3(n281_3));
  bfr _b_972(.a(_w_1393),.q(_w_1394));
  bfr _b_741(.a(_w_1162),.q(_w_1163));
  bfr _b_910(.a(_w_1331),.q(_w_1332));
  bfr _b_911(.a(_w_1332),.q(_w_1333));
  and_bi g266(.a(n264),.b(n265),.q(n266));
  bfr _b_913(.a(_w_1334),.q(_w_1335));
  bfr _b_917(.a(_w_1338),.q(_w_1339));
  bfr _b_918(.a(_w_1339),.q(_w_1340));
  bfr _b_920(.a(_w_1341),.q(_w_1342));
  bfr _b_923(.a(_w_1344),.q(_w_1345));
  bfr _b_1182(.a(_w_1603),.q(_w_1604));
  bfr _b_929(.a(_w_1350),.q(_w_1351));
  bfr _b_717(.a(_w_1138),.q(_w_1139));
  bfr _b_930(.a(_w_1351),.q(_w_1352));
  bfr _b_1492(.a(_w_1913),.q(_w_1914));
  bfr _b_1392(.a(_w_1813),.q(n252_1));
  and_bb g323(.a(n229_7),.b(n318_1),.q(n323));
  bfr _b_931(.a(_w_1352),.q(_w_1353));
  bfr _b_932(.a(_w_1353),.q(_w_1354));
  bfr _b_933(.a(_w_1354),.q(_w_1355));
  and_bi g94(.a(n92),.b(n93),.q(n94));
  bfr _b_848(.a(_w_1269),.q(_w_1270));
  bfr _b_1006(.a(_w_1427),.q(n231));
  bfr _b_934(.a(_w_1355),.q(_w_1356));
  bfr _b_937(.a(_w_1358),.q(_w_1359));
  bfr _b_941(.a(_w_1362),.q(_w_1363));
  bfr _b_945(.a(_w_1366),.q(_w_1367));
  bfr _b_1382(.a(_w_1803),.q(_w_1804));
  bfr _b_948(.a(_w_1369),.q(G21_5));
  bfr _b_949(.a(_w_1370),.q(_w_1371));
  bfr _b_950(.a(_w_1371),.q(_w_1372));
  bfr _b_973(.a(_w_1394),.q(_w_1395));
  bfr _b_955(.a(_w_1376),.q(_w_1377));
  bfr _b_761(.a(_w_1182),.q(_w_1183));
  bfr _b_975(.a(_w_1396),.q(_w_1397));
  bfr _b_1015(.a(_w_1436),.q(_w_1437));
  bfr _b_956(.a(_w_1377),.q(_w_1378));
  bfr _b_1209(.a(_w_1630),.q(_w_1631));
  bfr _b_960(.a(_w_1381),.q(_w_1382));
  bfr _b_961(.a(_w_1382),.q(_w_1383));
  bfr _b_1353(.a(_w_1774),.q(G1353));
  bfr _b_962(.a(_w_1383),.q(_w_1384));
  bfr _b_963(.a(_w_1384),.q(_w_1385));
  spl2 g374_s_0(.a(n374),.q0(n374_0),.q1(n374_1));
  bfr _b_969(.a(_w_1390),.q(_w_1391));
  bfr _b_1284(.a(_w_1705),.q(_w_1706));
  bfr _b_1252(.a(_w_1673),.q(_w_1674));
  bfr _b_974(.a(_w_1395),.q(_w_1396));
  bfr _b_976(.a(_w_1397),.q(_w_1398));
  bfr _b_980(.a(_w_1401),.q(_w_1402));
  bfr _b_983(.a(_w_1404),.q(_w_1405));
  bfr _b_736(.a(_w_1157),.q(_w_1158));
  bfr _b_987(.a(_w_1408),.q(_w_1409));
  bfr _b_988(.a(_w_1409),.q(_w_1410));
  bfr _b_989(.a(_w_1410),.q(_w_1411));
  bfr _b_992(.a(_w_1413),.q(_w_1414));
  bfr _b_1001(.a(_w_1422),.q(_w_1423));
  bfr _b_994(.a(_w_1415),.q(_w_1416));
  bfr _b_997(.a(_w_1418),.q(_w_1419));
  and_bb g44(.a(G17_1),.b(G19_1),.q(n44));
  bfr _b_998(.a(_w_1419),.q(_w_1420));
  spl2 g316_s_1(.a(n316_1),.q0(n316_2),.q1(_w_1692));
  bfr _b_1002(.a(_w_1423),.q(G31_5));
  bfr _b_1004(.a(_w_1425),.q(_w_1426));
  bfr _b_1007(.a(_w_1428),.q(_w_1429));
  bfr _b_1010(.a(_w_1431),.q(_w_1432));
  bfr _b_986(.a(_w_1407),.q(_w_1408));
  bfr _b_1011(.a(_w_1432),.q(_w_1433));
  bfr _b_1487(.a(_w_1908),.q(_w_1909));
  bfr _b_1012(.a(_w_1433),.q(_w_1434));
  bfr _b_1013(.a(_w_1434),.q(_w_1435));
  bfr _b_1331(.a(_w_1752),.q(_w_1753));
  and_bb g239(.a(G3_1),.b(G7_1),.q(n239));
  bfr _b_946(.a(_w_1367),.q(_w_1368));
  bfr _b_1017(.a(_w_1438),.q(_w_1439));
  bfr _b_1020(.a(_w_1441),.q(_w_1442));
  bfr _b_1021(.a(_w_1442),.q(_w_1443));
  bfr _b_800(.a(_w_1221),.q(_w_1222));
  bfr _b_1026(.a(_w_1447),.q(_w_1448));
  bfr _b_1030(.a(_w_1451),.q(_w_1452));
  and_bi g284(.a(n282_1),.b(G1_7),.q(n284));
  bfr _b_1032(.a(_w_1453),.q(_w_1454));
  bfr _b_1034(.a(_w_1455),.q(_w_1456));
  bfr _b_1036(.a(_w_1457),.q(n153_1));
  bfr _b_1037(.a(_w_1458),.q(G1354));
  bfr _b_1285(.a(_w_1706),.q(_w_1707));
  bfr _b_687(.a(_w_1108),.q(_w_1109));
  bfr _b_1038(.a(_w_1459),.q(_w_1460));
  bfr _b_680(.a(_w_1101),.q(_w_1102));
  bfr _b_1046(.a(_w_1467),.q(_w_1468));
  bfr _b_822(.a(_w_1243),.q(_w_1244));
  bfr _b_1050(.a(_w_1471),.q(_w_1472));
  bfr _b_1452(.a(_w_1873),.q(_w_1874));
  bfr _b_1051(.a(_w_1472),.q(_w_1473));
  and_bb g139(.a(G20_4),.b(G24_4),.q(n139));
  bfr _b_954(.a(_w_1375),.q(_w_1376));
  bfr _b_936(.a(_w_1357),.q(_w_1358));
  bfr _b_1053(.a(_w_1474),.q(_w_1475));
  bfr _b_1185(.a(_w_1606),.q(_w_1607));
  bfr _b_1059(.a(_w_1480),.q(_w_1481));
  bfr _b_1223(.a(_w_1644),.q(G15_5));
  bfr _b_1062(.a(_w_1483),.q(_w_1484));
  bfr _b_1064(.a(_w_1485),.q(G29_5));
  bfr _b_1065(.a(_w_1486),.q(_w_1487));
  bfr _b_978(.a(_w_1399),.q(n191_4));
  bfr _b_1107(.a(_w_1528),.q(_w_1529));
  bfr _b_1070(.a(_w_1491),.q(_w_1492));
  bfr _b_1072(.a(_w_1493),.q(_w_1494));
  bfr _b_1184(.a(_w_1605),.q(_w_1606));
  bfr _b_1074(.a(_w_1495),.q(_w_1496));
  bfr _b_1076(.a(_w_1497),.q(_w_1498));
  bfr _b_1438(.a(_w_1859),.q(_w_1860));
  bfr _b_1078(.a(_w_1499),.q(_w_1500));
  bfr _b_881(.a(_w_1302),.q(_w_1303));
  bfr _b_1080(.a(_w_1501),.q(_w_1502));
  bfr _b_1084(.a(_w_1505),.q(_w_1506));
  spl2 g231_s_0(.a(n231),.q0(n231_0),.q1(n231_1));
  bfr _b_1088(.a(_w_1509),.q(G1349));
  bfr _b_805(.a(_w_1226),.q(_w_1227));
  bfr _b_1089(.a(_w_1510),.q(_w_1511));
  bfr _b_1090(.a(_w_1511),.q(_w_1512));
  bfr _b_1094(.a(_w_1515),.q(_w_1516));
  bfr _b_1099(.a(_w_1520),.q(_w_1521));
  bfr _b_1101(.a(_w_1522),.q(_w_1523));
  bfr _b_1104(.a(_w_1525),.q(_w_1526));
  bfr _b_1558(.a(_w_1979),.q(_w_1980));
  bfr _b_1108(.a(_w_1529),.q(_w_1530));
endmodule
