module c3540 (G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G6,G7,G8,G9,G3519,G3520,G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540);
  input G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G6,G7,G8,G9;
  output G3519,G3520,G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540;
  wire _w_3570,_w_3567,_w_3566,_w_3565,_w_3563,_w_3557,_w_3556,_w_3555,_w_3554,_w_3553,_w_3552,_w_3551,_w_3549,_w_3548,_w_3547,_w_3546,_w_3545,_w_3543,_w_3541,_w_3540,_w_3539,_w_3537,_w_3533,_w_3526,_w_3525,_w_3523,_w_3521,_w_3518,_w_3516,_w_3515,_w_3514,_w_3509,_w_3508,_w_3507,_w_3506,_w_3504,_w_3502,_w_3501,_w_3498,_w_3497,_w_3494,_w_3491,_w_3490,_w_3486,_w_3485,_w_3483,_w_3482,_w_3480,_w_3479,_w_3478,_w_3476,_w_3475,_w_3474,_w_3472,_w_3471,_w_3465,_w_3462,_w_3564,_w_3461,_w_3460,_w_3459,_w_3454,_w_3453,_w_3451,_w_3449,_w_3448,_w_3447,_w_3446,_w_3445,_w_3444,_w_3442,_w_3439,_w_3438,_w_3437,_w_3436,_w_3435,_w_3434,_w_3432,_w_3431,_w_3427,_w_3426,_w_3423,_w_3422,_w_3421,_w_3419,_w_3414,_w_3413,_w_3410,_w_3409,_w_3408,_w_3466,_w_3407,_w_3404,_w_3402,_w_3401,_w_3394,_w_3391,_w_3389,_w_3385,_w_3384,_w_3380,_w_3560,_w_3371,_w_3369,_w_3367,_w_3364,_w_3361,_w_3359,_w_3357,_w_3355,_w_3354,_w_3353,_w_3350,_w_3348,_w_3347,_w_3346,_w_3343,_w_3340,_w_3337,_w_3335,_w_3334,_w_3333,_w_3332,_w_3331,_w_3329,_w_3328,_w_3327,_w_3324,_w_3318,_w_3316,_w_3313,_w_3310,_w_3309,_w_3308,_w_3307,_w_3306,_w_3305,_w_3416,_w_3304,_w_3301,_w_3300,_w_3358,_w_3299,_w_3298,_w_3297,_w_3296,_w_3294,_w_3293,_w_3292,_w_3290,_w_3289,_w_3288,_w_3286,_w_3285,_w_3283,_w_3279,_w_3278,_w_3277,_w_3276,_w_3275,_w_3272,_w_3271,_w_3269,_w_3268,_w_3265,_w_3263,_w_3262,_w_3261,_w_3260,_w_3259,_w_3257,_w_3255,_w_3253,_w_3252,_w_3249,_w_3248,_w_3246,_w_3243,_w_3241,_w_3239,_w_3238,_w_3233,_w_3231,_w_3230,_w_3229,_w_3228,_w_3223,_w_3222,_w_3251,_w_3221,_w_3219,_w_3217,_w_3216,_w_3215,_w_3212,_w_3211,_w_3208,_w_3206,_w_3205,_w_3204,_w_3203,_w_3199,_w_3382,_w_3198,_w_3197,_w_3196,_w_3194,_w_3189,_w_3188,_w_3182,_w_3178,_w_3175,_w_3172,_w_3171,_w_3169,_w_3168,_w_3192,_w_3166,_w_3164,_w_3163,_w_3161,_w_3160,_w_3159,_w_3157,_w_3234,_w_3156,_w_3155,_w_3152,_w_3150,_w_3147,_w_3146,_w_3145,_w_3137,_w_3134,_w_3133,_w_3132,_w_3131,_w_3128,_w_3126,_w_3123,_w_3121,_w_3120,_w_3464,_w_3117,_w_3116,_w_3114,_w_3112,_w_3107,_w_3106,_w_3105,_w_3496,_w_3104,_w_3452,_w_3102,_w_3097,_w_3094,_w_3088,_w_3086,_w_3077,_w_3074,_w_3073,_w_3065,_w_3064,_w_3455,_w_3062,_w_3061,_w_3060,_w_3059,_w_3057,_w_3056,_w_3054,_w_3173,_w_3053,_w_3051,_w_3048,_w_3046,_w_3045,_w_3041,_w_3037,_w_3035,_w_3034,_w_3033,_w_3030,_w_3028,_w_3026,_w_3025,_w_3023,_w_3022,_w_3020,_w_3018,_w_3345,_w_3017,_w_3016,_w_3015,_w_3013,_w_3010,_w_3411,_w_3009,_w_3008,_w_3005,_w_3004,_w_2999,_w_2998,_w_2997,_w_2996,_w_2995,_w_3519,_w_2993,_w_3174,_w_2992,_w_2991,_w_2990,_w_2984,_w_2980,_w_2979,_w_2977,_w_2976,_w_2975,_w_2974,_w_2972,_w_2971,_w_2968,_w_2966,_w_2965,_w_2964,_w_2963,_w_2962,_w_2960,_w_3542,_w_3024,_w_2956,_w_2955,_w_2951,_w_2949,_w_2947,_w_2970,_w_2945,_w_2942,_w_3363,_w_2941,_w_2939,_w_2936,_w_2933,_w_2932,_w_2931,_w_2929,_w_2928,_w_2926,_w_2924,_w_2917,_w_2915,_w_2914,_w_2912,_w_2911,_w_2910,_w_2909,_w_2908,_w_2907,_w_3374,_w_2906,_w_2905,_w_2904,_w_2903,_w_2900,_w_2899,_w_2898,_w_2934,_w_2897,_w_2895,_w_2892,_w_2890,_w_2888,_w_2886,_w_2887,_w_2885,_w_2883,_w_2881,_w_2879,_w_2877,_w_2875,_w_2873,_w_2872,_w_2870,_w_2864,_w_3395,_w_2863,_w_2862,_w_2861,_w_2860,_w_2859,_w_2858,_w_2855,_w_2854,_w_2852,_w_2851,_w_2849,_w_2848,_w_2847,_w_2845,_w_2844,_w_2843,_w_2840,_w_2839,_w_3532,_w_2836,_w_2834,_w_2833,_w_2988,_w_2831,_w_2830,_w_2829,_w_2827,_w_2824,_w_2819,_w_2818,_w_2817,_w_3295,_w_2809,_w_2807,_w_2805,_w_2804,_w_2803,_w_2802,_w_2800,_w_2799,_w_2797,_w_2793,_w_2790,_w_2788,_w_2787,_w_2786,_w_2784,_w_3084,_w_2783,_w_3377,_w_2782,_w_2780,_w_3398,_w_2779,_w_2776,_w_2774,_w_2773,_w_2772,_w_2882,_w_2770,_w_2769,_w_2767,_w_2766,_w_2763,_w_2761,_w_2760,_w_2759,_w_2758,_w_2756,_w_2753,_w_2752,_w_2751,_w_2749,_w_2748,_w_2747,_w_2930,_w_2746,_w_2745,_w_2744,_w_2742,_w_2740,_w_2739,_w_2738,_w_2737,_w_3038,_w_2735,_w_2734,_w_2733,_w_2732,_w_2731,_w_2730,_w_2729,_w_2725,_w_2724,_w_2723,_w_2720,_w_2717,_w_2716,_w_2714,_w_2712,_w_2711,_w_2709,_w_2706,_w_3456,_w_2705,_w_2704,_w_2703,_w_2822,_w_2702,_w_2700,_w_2698,_w_2697,_w_2696,_w_2695,_w_3287,_w_2694,_w_2693,_w_2691,_w_2690,_w_2687,_w_2684,_w_2681,_w_2680,_w_2678,_w_2677,_w_2676,_w_3534,_w_2953,_w_2675,_w_2674,_w_2673,_w_2671,_w_3090,_w_2669,_w_2666,_w_2665,_w_2664,_w_2663,_w_2662,_w_2660,_w_2655,_w_2653,_w_2652,_w_3050,_w_2650,_w_2649,_w_2648,_w_2647,_w_3181,_w_2646,_w_2645,_w_2643,_w_2642,_w_2641,_w_2640,_w_2639,_w_2708,_w_2638,_w_2636,_w_2896,_w_2632,_w_2627,_w_2626,_w_2667,_w_2623,_w_2622,_w_2978,_w_2620,_w_3527,_w_2619,_w_3561,_w_2618,_w_2617,_w_2614,_w_2612,_w_2610,_w_2609,_w_2605,_w_2604,_w_2603,_w_2601,_w_2599,_w_2598,_w_2595,_w_2594,_w_2593,_w_3220,_w_2592,_w_2591,_w_3063,_w_2590,_w_2589,_w_2587,_w_3495,_w_2586,_w_2585,_w_2994,_w_2584,_w_2583,_w_2582,_w_2581,_w_2579,_w_2578,_w_2657,_w_2577,_w_2575,_w_2573,_w_2571,_w_2944,_w_2569,_w_3517,_w_2568,_w_2567,_w_2566,_w_2564,_w_2562,_w_2561,_w_2560,_w_2565,_w_2559,_w_2557,_w_2555,_w_2554,_w_2551,_w_3100,_w_2935,_w_2550,_w_2549,_w_2546,_w_2544,_w_2543,_w_2542,_w_3122,_w_2541,_w_2539,_w_2536,_w_2534,_w_2533,_w_2532,_w_2528,_w_2527,_w_2524,_w_2523,_w_3176,_w_2522,_w_2519,_w_2517,_w_2516,_w_2515,_w_2514,_w_2512,_w_2511,_w_2810,_w_2510,_w_2868,_w_2506,_w_2505,_w_2821,_w_2503,_w_3368,_w_2501,_w_2499,_w_2497,_w_2496,_w_2492,_w_3424,_w_3320,_w_2490,_w_2489,_w_2487,_w_2718,_w_2486,_w_3085,_w_2713,_w_2485,_w_2483,_w_2482,_w_2481,_w_2480,_w_2478,_w_3058,_w_2572,_w_2477,_w_2472,_w_2468,_w_2467,_w_2466,_w_2465,_w_2464,_w_2507,_w_2462,_w_2461,_w_2459,_w_2458,_w_2457,_w_3405,_w_2456,_w_3226,_w_2455,_w_2454,_w_2453,_w_2451,_w_2850,_w_2450,_w_2449,_w_2446,_w_2445,_w_2443,_w_2442,_w_2440,_w_2438,_w_2437,_w_2435,_w_3467,_w_3415,_w_2434,_w_2432,_w_2428,_w_2427,_w_2811,_w_2425,_w_2424,_w_2422,_w_2421,_w_3111,_w_2420,_w_3477,_w_2419,_w_2418,_w_2417,_w_2414,_w_2412,_w_2410,_w_2408,_w_2406,_w_2405,_w_2404,_w_2403,_w_2741,_w_2402,_w_2401,_w_2399,_w_2398,_w_2397,_w_2396,_w_2395,_w_2894,_w_2394,_w_2393,_w_3512,_w_3096,_w_3021,_w_2710,_w_2392,_w_2390,_w_2389,_w_2388,_w_2391,_w_2386,_w_2385,_w_2384,_w_2615,_w_2383,_w_2382,_w_3473,_w_2381,_w_2631,_w_2380,_w_2379,_w_2377,_w_2375,_w_2373,_w_2488,_w_2372,_w_2371,_w_3069,_w_2368,_w_2366,_w_2365,_w_2362,_w_2361,_w_2360,_w_2358,_w_2357,_w_3109,n630,n127,n581_0,n135_4,n559_0,n372_5,_w_2644,n135_0,n372_10,n553_3,n137_4,n536,n751,_w_2247,n137_1,n137_0,n240_3,G37_1,_w_2433,n129_8,_w_2144,n572_1,n572_0,n148_1,G3535_2,G11_15,G3535_1,n149_3,n361_14,n374_6,n149_1,n123_6,n123_5,n151_7,n151_3,n151_2,_w_3323,n533_5,n363,n250_0,_w_2178,_w_2426,n151_1,_w_3378,n455_1,n107,n455_0,G12_15,n659,G12_12,_w_2283,_w_3195,G12_11,G12_10,G12_7,G12_6,n145_5,n582,G12_3,n185_0,n495_1,n214_2,n214_1,n593,_w_3388,n214_0,n388,_w_2218,n162_8,G7_3,n162_5,G19_1,_w_3284,n401_24,n162_3,_w_3280,n533,_w_3530,n372_7,n74_0,_w_2954,n162_10,n392_14,n392_11,n568,n392_10,_w_2113,n392_3,n287,n437_0,n216_1,n171_0,n831,G47_5,_w_3529,_w_3191,n130_3,G47_4,n830,G3531_0,G47_1,_w_3470,G8_12,_w_3218,_w_2206,n537_0,G3535_0,n201_0,_w_3186,n134,n105_0,G7_8,n88_1,n398_13,n295_1,n746,n235_0,n627_0,n533_7,n124,n385_14,_w_3400,_w_2969,n533_4,n533_1,n372_1,n534_1,_w_3082,_w_2823,n540_2,n540_0,n254_0,_w_2553,n629_1,_w_3052,n130,n549_1,_w_2470,G10_3,_w_3071,n554_1,n566_1,n54_0,n654_0,n315,_w_2880,n224_1,n521,n553_1,_w_2545,_w_2314,n832_1,_w_3154,n381_9,n765_1,n224_2,n523,n683_2,G4_44,n688_3,G11_12,G20_3,n688_0,G4_14,n696_0,n384,n554_2,n813_1,n320,n701_1,G13_2,n201_1,_w_2125,n457,_w_2143,n812_1,G43_3,n130_0,n829_0,n688_1,n836,n829,n822_1,n828,n827,_w_2987,n825,_w_2239,n824,G9_19,_w_3245,n823,_w_3488,_w_2448,n422,n385_20,n821,n130_1,n701_0,_w_2866,_w_2679,n819,_w_2529,G30_5,_w_2563,n604_1,n302,_w_2348,n813,n441,_w_3468,n812_0,n372_6,n808,n807,n806,n804,n159_1,n802,n495_0,n801,n190_1,n795,_w_2370,n792,_w_2224,n542_0,n419_0,n791,n758,n176_3,n790,G17_2,n788,n546_2,n553_0,_w_3190,_w_2891,_w_2670,n670,n775,_w_3099,_w_3031,G7_16,n812,_w_3379,G9_1,n773,n143_9,n143_11,_w_2701,G24_6,_w_2495,n770,n761,n367,n320_2,_w_2973,n756,_w_2474,n822,n755,n754,n753,n752,n601,n334,n768,n634,n742,_w_3522,G35_2,n737,n734,n381_1,n730,_w_2537,n395_0,n729,n112,n398_10,_w_2791,n725,G37_3,n560,n338_1,_w_2835,n748,G39_1,n724,G7_13,n723,n261,n395_10,_w_3425,G7_20,n135_2,n75_0,_w_3118,n719,n718,n490_6,_w_2814,n99,_w_2513,n715,n713,n119,n710,_w_3342,n738,_w_2867,_w_2400,n709,n484_0,n707,n94_0,G20_6,n706,n295,G11_8,n705,n410,n401,G17_1,n696,_w_2508,n590,_w_3012,n690,n176_2,n687,n459,G4_32,n490_4,n151_9,n162_9,n826,n392_7,G4_31,_w_3319,n126_0,_w_3042,n151_6,n129_4,_w_2430,n84,n240_6,n129_1,G20_5,_w_2248,n676,n240_0,n674,_w_2538,n765,_w_2305,n176_0,n361_17,n673,n672,n144,n667,_w_2806,n665,_w_2270,n217,n826_0,_w_2837,n662,n656,n444,_w_3387,n560_1,n616,n627_1,n558,n640,n551_0,_w_2334,n805,n639,G21_9,n563_0,n164_0,n628,n327,_w_2407,n800,_w_3430,n627,G24_7,n661,G14_12,n622,G12_5,_w_3336,_w_2961,n143_0,_w_2838,n613,n620,n619,_w_2137,n618,n306_0,n617,G42_1,n615,n610,_w_2260,G4_33,G14_17,n700,n607,n605,n149,G3_14,G8_6,n411_1,n602,G21_0,_w_3544,n600,_w_2278,n599,n212,G10_13,n202,G40_5,_w_2525,G1_1,n382_0,_w_2423,n201_3,_w_3079,G47_0,n272,n648,n597,_w_2755,n654,n578,n293_0,n595,G3_8,G3_24,n589,n587_1,n588,n587,n542,n586,n535_0,_w_3536,n585,n626,n584,n684_1,n361_11,n712,n191_1,n666,G39_4,G47_3,n72,n575,n377_2,n306,_w_2479,n293_1,n570,n567,_w_2801,n566,n733,n581,G11_13,_w_3339,n835,_w_3127,_w_2878,n436_0,n565,n129_2,n379_2,_w_2637,n561,n344_0,n769,n556,n171_1,n554,n587_0,n669,n552,_w_2460,_w_2298,n551,n54,n408_0,n223,n549,n77_0,n392_1,n398_9,_w_3183,n545,n385_18,_w_2921,_w_2796,n544,G36_2,n708,n541,n368,n540,n537,n579,n149_2,n534,n74_1,G11_2,n832_0,n771,n532,n632,_w_3119,n505_0,n402,n811_2,_w_2376,n228,n162_0,n505_1,_w_3571,n843,n361_13,_w_2221,n342,n235,n232,G12_18,_w_2820,n392_13,n475,n732_0,n230,n401_19,n220,G3_21,_w_2181,_w_2313,n162_6,n686,n338_2,n635,G4_13,_w_3214,n219,n162_7,n213,_w_2194,_w_2600,n353,_w_3266,n741,_w_2531,n778,n477,_w_2919,n824_1,G11_11,n115,_w_2439,G9_14,n66,_w_3341,n362_0,n97,_w_3356,n314,_w_2686,_w_2204,n766,n813_0,n737_0,n216,_w_3338,n728,n201,G9_17,G3526_3,n373,n147_7,_w_2633,n123_8,n785,_w_3412,_w_2986,n247,G14_0,_w_3101,_w_2794,n320_1,n500_0,_w_2198,n229,_w_2699,G3531_3,_w_2668,n657,G18_2,_w_2359,n254_1,n695_2,n309,G41_2,n188,n183,n307,_w_2494,n171,n354,_w_3254,G47_2,G19_3,n524,n165,_w_2940,n392,_w_3075,n88,n143_2,_w_3193,n194,n517,_w_2596,n789,n480_1,n162,n62,G30_2,_w_3151,n678,n299_0,n496_0,n668,_w_2901,n458,G20_2,n214,G3_3,n554_0,_w_2750,n123_7,_w_3141,_w_2726,n495,n236,n727,n138,n638,n443,n75_1,n147_10,_w_3153,n193,n658,n663,n184,n123_3,_w_3177,n772_0,n157,n462,n361_20,n155,_w_3072,_w_3007,n180,n621,n77_1,_w_2127,_w_2179,n548_0,n833,n152,G11_4,n162_2,n560_0,n696_2,n250_3,n110,n74,n624,_w_3067,_w_2411,n150,n374_5,n123,n105_1,_w_2608,_w_2558,G14_4,n735_2,_w_3568,_w_2621,n694,n137_2,n162_4,n350,n566_0,n419,G4_11,n141,n505,n612,n572,_w_3201,n398_7,G24_2,_w_3311,_w_2884,G6_0,n596,_w_2160,n104,_w_2958,G27_3,_w_2902,n669_1,_w_2229,n684,n699,n240,n580,n288,n139,n137,n484,G18_1,_w_3235,n553,n681,n198,n454,_w_2727,n629,n204,n693,_w_3383,n430,n137_5,n168,_w_2841,G3_1,n136,n235_1,_w_2692,n118,n231,_w_3092,n85_1,_w_2216,_w_2227,n604,_w_3170,n135,n548,n461,n290,G35_8,_w_2228,G3528_0,n372_9,n123_4,n685,n135_1,n571,n129,n517_0,_w_2364,n826_1,n493,G3532_3,n392_6,G5_2,n256,_w_3140,G33_4,G10_8,_w_2441,n451,n784,n352,_w_3247,n385_19,n757,G22_8,_w_3403,_w_2205,n120,_w_3076,G1_12,n781,n722,G12_17,n221,n732_1,n206,_w_2656,n321_0,n361_4,n187,n803,n497_0,_w_2736,n669_0,n815,n125,n101,_w_2981,n604_0,n551_1,n559,G22_2,n655,_w_2243,n178,n154,n645,n170,n401_21,G23_0,n161_1,n501,n192,_w_3047,_w_2498,G3_12,n423,G40_0,n838_0,n215_0,n406,_w_3362,n384_1,n146,_w_2447,n762,G12_1,_w_2625,n128,n321,n249,n189_0,n166,n392_4,n467,_w_3349,_w_3044,_w_2688,G34_5,_w_2871,n301,n623,_w_3237,n133,G31_2,n341,_w_2242,n839,G4_5,n298_1,n111,G9_16,G14_2,n280,n322,_w_3429,n205,n598,n520,n286,n267_1,_w_3242,n428,n90,G3534_1,n196,_w_2126,n737_1,G3_20,n420_0,G11_3,n143_5,n636,n175,G1_3,n176,_w_2946,G1_5,G21_4,n653,n57,n77,n162_1,_w_3029,n496_2,_w_2154,n191,n98,n537_1,n591,n73_0,G12_16,_w_3558,_w_2324,n395_8,n250_2,_w_3326,_w_2281,n482,n117,n94,_w_3210,n408_1,n197,n543_0,n325,n692,n375,n745,_w_2580,n81,n543,n160,G7_19,n780,n564,n52_1,_w_2607,n740,_w_2171,n557,n190_0,n395,G34_6,n400,n306_3,_w_3489,n842,n73_3,G36_6,n106,_w_2869,n145_6,n447,n413,n339,_w_3520,G2_6,n343_2,_w_3162,n153,_w_2150,n398,n569,_w_3487,n772_1,n417,_w_2431,n123_2,n121,n275_0,n606,_w_2889,n546_3,n174,_w_3006,_w_2344,n200,_w_2927,_w_2658,_w_2186,_w_3500,_w_3184,n735_3,_w_2322,_w_2502,n744,G4_26,_w_2225,n535,n125_0,n539,_w_3225,_w_2826,n71,_w_3240,_w_2754,n651,_w_2349,n390,n164_1,n191_0,n201_2,n649,n116,n487,_w_2982,n392_8,n303,_w_2363,n234,G4_50,n438,n225,n540_1,n507_0,_w_3321,_w_2920,n332,_w_3428,n445,n703,_w_2325,n630_1,n716,n764,n559_1,G3536_0,_w_2957,G3529_2,n503,n61,n449,n553_2,n73,n743,_w_3036,n395_1,n56,G22_1,n75,n58,G4_43,n389,_w_3569,n392_12,n59,n60,_w_3511,_w_2781,n480,_w_2413,G4_8,_w_3492,n129_5,n483,G4_40,G9_10,n691,n227,_w_3270,n720,n316,_w_3572,n494_3,_w_2219,n404,G33_3,n485,_w_3538,_w_2191,n145,G22_9,_w_3366,n147,n664,n361,n64,_w_3344,_w_2147,_w_2266,n275,G25_0,_w_3080,_w_3032,_w_2570,n300,n542_1,n497,_w_2416,n401_18,n68,n711,_w_2597,n270,G18_0,n76,_w_2816,n277,G20_1,_w_3207,n436_3,n509,n427,n347,n51_2,n195,_w_3165,_w_2249,_w_2846,n637,n527,n305,n392_9,n96,_w_3440,n73_1,n543_1,n156,n293,n533_6,n464,n629_2,n52,_w_2634,n83,n79,n395_2,_w_2948,n502,_w_3312,n181,n85,n547,G8_14,_w_3373,_w_3142,n549_0,n87,G3_4,n163,n507_2,n105,_w_2683,n243,n238,_w_2916,n372_4,G3535_3,n378,n714,n697,n246,n440,n291,_w_2473,n86,n250_1,_w_2813,n250,G13_12,G39_7,n530,n838_1,n834,n428_0,n403,_w_2211,G1_0,_w_2287,n481,_w_2950,n611,n108,n528,n258,n365_0,n259,n385_21,n262,n143_6,_w_3103,_w_3014,G19_2,n500_4,G14_1,n255,n277_1,n392_5,n330,n317,n396,n767,_w_2330,_w_2355,n265,_w_2521,n421,_w_2415,n695_0,_w_2874,n574,n298,_w_3510,G12_2,n315_1,n109,n414,n269,n313,n534_0,G3536_2,n51_0,n123_10,n273,_w_2778,n274,n364,n344,_w_2484,n276,n609,n182,G3_17,n437_4,n279,G12_13,_w_2651,_w_2475,n281,G3_11,n362,_w_2174,n351,n455,n702,n282,n446,n407_2,n283,n499,_w_2574,n284,n293_3,n452,_w_3232,n285,G44_0,n365,_w_3535,_w_2163,n294,n501_0,n137_6,G48_1,n296,_w_2196,n399_1,n735_1,n372,n233,n52_2,n299_1,_w_2262,n70,n381_0,n297,_w_3291,n88_0,n736,n211,n299,G35_9,G7_5,_w_3418,_w_3365,n510,G29_0,G37_2,_w_2795,n199,_w_2547,_w_2369,n308,G22_5,n646,n239,_w_2246,n491,_w_2792,_w_2188,n395_15,n604_2,_w_3458,n358,_w_3244,n478,n165_2,n260,_w_2185,_w_2552,n91,n783,n787,n772,n260_3,n340_3,n208,n519,n328,n329,G11_5,_w_3493,_w_2444,n186,_w_3273,n526,n173,n335,n382_3,_w_2320,n338,n555,n420,n386_0,n135_3,n759,_w_2317,n340,n130_2,n511_0,_w_3202,n343,_w_3513,G40_3,n369,G14_7,n401_9,n840,_w_2267,n92,n348,n179_0,G3534_2,_w_2310,_w_3000,n357,n91_1,n210,G40_7,n424,n814,n360,n366,n237_1,n407,n418,_w_2387,n407_13,n592,_w_2985,n496_1,n515,n78,n264,n379,n240_4,_w_3450,n145_4,n324,n614,n411,n165_1,n110_1,_w_3443,n177,_w_2251,_w_2210,n383,n385,n321_1,n625,n386,n318,_w_3503,n387,_w_2471,G24_0,n508,n797,n513,n362_1,n242,n399,_w_2263,_w_2264,n129_9,_w_3393,n405,_w_2853,n381_8,n514,n546,n379_3,n491_1,G14_9,n837,G3526_1,n474,n829_1,n190,n89,n426,n240_2,n407_7,_w_3267,n652,n494_1,n409,n429,_w_2233,n433,_w_2159,n486,n562,n434,_w_2255,n501_2,n129_6,n563,n224_0,_w_2757,n490_0,n149_0,n114,_w_3322,_w_2122,_w_2832,n435,n436,n832_3,G4_17,n439,_w_3095,G4_7,_w_3282,n304,n216_0,n514_3,n129_3,n442,n56_1,n629_0,n533_3,G32_6,_w_2319,n51,_w_2765,G10_0,_w_3250,n472,_w_2296,G4_45,_w_2197,n224,n450,G24_5,n453,_w_2156,n793,n317_2,n148,G4_49,_w_2124,_w_3314,G24_1,n463,G13_15,n151_0,n774,n241,n654_1,G22_0,_w_2309,n93,n496,n573,n476,n469,n189,G13_8,n511,n747,n393,n100,n516,n125_1,n473,G12_0,n314_0,n358_0,n644,n267,n107_0,n479,_w_3390,G10_5,G7_17,_w_3528,n311,_w_2452,n548_1,n361_15,n697_0,n763,n395_9,n492,n298_0,G33_7,n683_0,n695,n129_0,n647,n798,n538,n237,n498,n143,n349,n360_0,_w_3138,n533_8,n500,n169,n63,_w_2409,n504,G32_0,n507,n704,n750,_w_2199,_w_3149,G13_6,n630_0,n518,n428_1,_w_3167,n643,n151_5,n215,_w_2943,G4_10,n265_4,n415,n525,n671,n529,n394_0,_w_3469,n240_5,G8_10,G12_4,n394_1,n653_0,n653_1,_w_2938,G1_8,G14_6,n123_9,n377_0,n377_1,n51_1,n377_3,n814_0,G33_0,G11_1,G33_1,G7_15,n94_1,G33_2,n796,G33_6,_w_2530,G11_0,n816,G32_1,_w_2768,G11_6,_w_3236,_w_2893,G3534_3,G11_9,G11_14,G11_16,G11_17,_w_3143,n361_2,G4_0,n696_1,G4_1,G4_38,_w_3352,G4_2,n67,n437_1,G24_4,G4_3,G4_4,G4_6,n381,G4_9,n395_3,n167,n511_1,n814_1,G4_12,G4_18,n91_0,_w_2220,G4_19,G4_20,_w_2292,_w_3125,n809,n832,G4_21,G4_22,G4_24,G4_27,G4_29,G4_30,G4_35,n292,G5_5,n113,G4_37,_w_3406,G4_39,G4_41,n721,n147_8,G4_42,G22_4,_w_3019,n123_0,G4_46,G4_47,G4_48,n159,G4_15,G3_13,_w_3093,G4_51,_w_2952,n97_0,_w_3531,n97_1,_w_2654,G44_2,G16_0,n130_4,n233_1,G16_1,G3533_0,G17_0,G17_3,_w_2200,n428_2,n398_16,G42_2,G9_0,G9_6,G9_2,n185,G9_3,n717,G9_4,G9_7,_w_3524,n401_16,G9_8,G41_8,n295_2,_w_2336,n490,G9_9,G14_11,G9_12,G9_13,n385_3,_w_2172,G9_15,n146_0,G32_2,n251,n146_1,G20_0,n726,n437_3,_w_2548,G20_4,_w_3264,n689_0,n398_12,_w_2328,n689_1,G29_1,_w_2842,G3536_1,G23_1,G50_1,G14_3,n132,G14_5,G14_8,n142_0,_w_2865,G14_10,n533_0,n148_0,n490_5,_w_2611,G14_13,G14_14,G3537_0,G14_16,_w_2812,n361_18,n338_0,G14_18,n401_4,G40_1,n431,G3_22,G40_2,n56_2,n331,G40_4,n448,n395_12,n374_2,_w_2771,G40_6,G40_8,n265_0,_w_3187,G40_9,G3_7,G8_7,n491_0,_w_2540,n786,n210_1,n298_2,n456,n176_1,n77_2,n501_1,n401_13,n683,G26_1,_w_3224,_w_3091,G26_2,n105_3,G26_3,_w_2798,n675,n399_0,n319,G27_0,G27_1,G27_2,n425,n314_1,G35_0,G35_1,_w_2661,_w_2476,G35_3,_w_3375,_w_2276,G35_5,n95,n361_7,G35_7,_w_2815,G3_0,n581_1,n688_2,n73_2,G33_5,n346,_w_2351,G3_2,n164,G3_5,G11_18,n306_1,G3_6,_w_2707,n822_0,_w_3087,G3_9,n392_2,G3_10,G3_15,_w_2300,_w_2504,G3_16,G3_18,_w_2722,_w_2526,G3_19,G3_25,G3_27,n407_1,G31_0,_w_2775,n436_1,_w_2288,n172,G31_1,_w_3376,_w_2491,G31_3,n401_12,n514_0,_w_2764,n509_1,G31_5,n56_0,_w_2187,G31_6,_w_3399,G3528_2,G31_7,n374_8,G14_19,G3529_0,n832_2,n533_2,G3529_1,G3529_3,n679,n680,G3532_2,n179_1,G42_0,n692_1,G36_0,G36_1,G36_4,_w_3396,G36_5,n145_0,G36_7,_w_2128,n385_11,G38_0,G38_1,G34_0,_w_2576,G34_1,n401_20,_w_2306,n631,G34_4,G34_7,G43_0,G35_4,_w_2331,G34_8,G9_18,n401_6,G3533_1,G4_36,G3533_2,G37_0,G3533_3,n506,n107_1,G39_0,G1_4,G8_8,_w_3070,G39_2,G39_5,G39_6,G39_8,G39_9,n563_1,G39_10,_w_3115,G39_11,_w_3001,n190_2,G6_2,G19_4,n494_0,n310,n494_4,n395_6,n395_7,n395_11,_w_3463,n207,n395_13,n395_14,n329_2,n395_18,n374_7,_w_3110,_w_2602,n395_19,G41_0,G41_1,n358_1,n179,G41_3,G9_11,n383_0,n361_10,G41_5,_w_2290,G41_6,_w_3136,G41_7,n126_1,n126_3,G5_0,G5_1,G34_2,G5_3,G5_6,n460,_w_2327,_w_2918,n623_0,_w_3397,n379_7,n623_1,n490_1,_w_3213,n145_2,_w_2202,n490_2,n490_3,_w_2743,n732,G1_2,n252,G1_6,_w_2165,G1_7,G1_9,_w_2913,G8_4,G9_5,_w_2114,G1_10,G1_11,n113_0,n517_1,n385_4,n113_1,G50_0,_w_3144,n153_0,_w_2518,n381_6,_w_2989,n392_0,n395_5,n153_1,_w_2762,G3532_0,_w_3420,n398_4,G3532_1,n315_0,_w_2193,G10_1,n397,G10_2,G10_4,n398_2,G10_6,_w_3180,G10_7,_w_3158,n65,G10_9,n735,G10_10,G10_11,n407_6,G10_12,_w_3317,n312,G10_14,n116_1,n395_4,G3528_1,G44_1,G3528_3,G3531_1,_w_3185,n385_8,G3531_2,n379_5,G11_7,n284_0,G32_3,_w_3148,G32_4,G32_5,n356,n692_0,G30_0,_w_3303,G30_1,G30_3,n633,n407_9,_w_2280,n468,n253,G30_4,_w_3011,G30_6,G31_4,G21_1,n401_1,n799,G13_0,G21_2,_w_3066,_w_2192,G21_3,G21_5,n100_1,n522,G21_6,G21_7,G8_5,n240_1,G21_8,G25_1,_w_2630,n481_0,G3537_1,_w_2268,n73_4,n73_5,G43_1,G18_3,n161,G43_2,G13_13,G2_0,n140,n142,G2_1,n379_10,_w_3499,G2_2,n283_1,G2_3,n433_1,_w_2183,G2_4,n385_5,G2_5,_w_2613,n480_0,G2_8,n370,G3526_0,n227_0,n227_1,n145_1,_w_2157,n145_3,_w_2469,n147_1,n398_21,n677,n382_2,n147_4,n147_5,n147_6,n147_9,n147_11,n361_1,n642,n394,n361_3,G3526_2,n361_5,n257,n361_6,n361_8,n701,n361_9,n361_12,_w_3351,_w_3281,n361_16,G4_23,n361_19,_w_3256,n385_12,n377,n275_1,_w_3370,n270_0,n577,n315_3,n270_1,n381_5,_w_3315,_w_3108,n382_1,n594,_w_2299,_w_3083,G2_7,n509_0,n54_1,n263,n238_1,n54_2,_w_3130,n69,G13_9,n293_2,_w_2333,n52_0,G12_8,n161_0,n85_0,_w_2721,n147_2,n105_2,_w_2340,n116_0,n105_4,_w_3179,n105_5,_w_2606,n238_0,n268,n238_2,n185_1,G3534_0,n697_1,n834_1,_w_2155,n834_2,n834_3,n834_4,_w_2367,n550,n147_0,n834_5,n481_1,n254_2,_w_3417,n433_0,n215_3,n563_2,n385_10,n563_3,_w_2689,n333,G8_9,n317_0,_w_2158,_w_3274,n317_1,_w_2346,G12_9,n102,n317_3,_w_3129,n660,n265_1,n265_2,n265_3,_w_3550,n151_8,n269_0,n269_1,n344_1,_w_2212,n779,G7_7,_w_2207,_w_2304,_w_2520,n407_3,n407_4,_w_2463,n407_5,n129_7,n244,n407_10,G7_14,n407_11,_w_2509,n158,n407_12,n237_2,n407_14,n277_2,n283_0,_w_2177,n189_1,n282_1,n385_16,_w_2857,n282_2,_w_2685,n271,n218,n282_3,n380,n283_2,n283_3,n284_1,_w_2825,n284_2,G7_1,G7_2,G7_9,_w_3003,n379_6,G7_10,G7_11,G7_12,_w_2876,_w_2232,G7_18,_w_3372,n372_0,n372_2,G4_25,n372_3,_w_3258,_w_3068,n372_8,n159_0,n323,_w_2245,n372_11,G4_52,_w_2214,n277_0,_w_2341,n226,_w_2293,n372_12,n512_0,n192_0,n192_1,n282_0,n192_2,G48_0,n192_3,n137_3,n329_0,_w_2983,n470,_w_2231,G22_3,G22_6,n289,_w_2269,G22_7,n398_0,n398_1,G24_3,n398_3,n398_5,n398_6,n351_0,n398_8,n398_14,_w_2777,_w_2715,n398_17,_w_2789,n123_1,n760,n379_1,n398_19,n484_1,G39_3,n398_20,G3_23,G8_17,_w_3227,_w_2289,n142_1,n142_2,n260_0,n260_1,n260_2,_w_2429,n460_0,n320_3,n222,_w_2190,n838,n749,n320_4,G7_4,n343_0,n329_1,n329_3,G8_0,G32_7,G8_1,G8_3,G8_11,n337_0,n366_0,_w_2356,n398_11,G8_15,G10_15,G8_16,_w_2354,G8_18,n337_1,n420_1,n834_0,n340_0,n340_1,n735_0,n209,n343_1,n369_0,_w_2923,n248,n369_1,_w_2728,_w_2672,n369_2,n369_3,G5_4,G19_5,_w_3481,n391,n351_1,n407_8,n811_0,n270_2,n379_8,n811_1,n360_1,n365_1,_w_3484,n365_2,G7_0,n466,n265_5,_w_2273,n151,n366_1,n100_0,n374_0,n126,n374_1,_w_3330,n698,n374_4,n374_3,n374_9,n374_10,n379_0,n320_0,n428_3,n379_4,n379_9,n379_11,_w_3505,n379_12,n237_0,_w_3457,_w_3089,n237_3,n381_2,n650,n126_2,_w_2323,n381_3,n381_4,n381_7,n383_1,n385_1,n337,n385_2,n385_6,G11_10,n385_7,n385_9,n385_13,_w_3113,n684_0,n416,n385_17,n386_1,_w_2659,G13_20,n401_0,_w_3049,n401_2,n401_3,_w_2629,_w_2535,n401_5,n315_2,n401_7,n401_8,n401_10,_w_3200,n739,n401_11,_w_2335,n395_17,n401_14,_w_2588,_w_2175,_w_2374,G36_3,n401_15,n401_17,_w_3360,n401_22,n583,n278,n401_23,n131,n437_2,_w_3027,n576,n336,n409_0,n409_1,n411_0,_w_3392,n546_0,n165_0,n546_1,_w_2343,_w_3078,n266,n535_1,n436_2,_w_2164,n465,n436_4,_w_2235,n436_5,_w_2112,n51_4,n51_5,_w_2436,n460_1,_w_3135,n189_2,n119_1,n340_2,n267_0,n482_0,G3536_3,n306_2,n482_1,G3_26,G42_3,G42_4,n695_1,G42_5,n494_2,G13_1,n245,_w_2123,G7_6,G13_3,n608,G13_4,n385_0,_w_2222,G13_5,G13_7,_w_3043,G1_13,n488,G13_10,G41_4,G13_14,G13_16,_w_3139,G13_17,G13_18,G13_19,G14_15,G13_21,_w_2237,n688,n497_1,G13_11,n143_1,_w_2616,n143_3,n77_3,n398_15,_w_2140,n143_4,n776,n143_7,G4_16,n143_8,n143_10,G26_0,n500_1,n295_0,n500_2,n500_3,n500_5,n507_1,n512_1,n514_1,n412,n514_2,n514_4,n631_0,n631_1,n215_1,n215_2,n521_0,n151_4,G35_6,n521_1,G6_1,_w_2111,n80,_w_2115,n419_1,_w_2116,_w_2635,n203,n765_0,_w_2117,G34_3,_w_2118,G19_0,_w_2119,_w_2134,_w_2350,_w_2120,_w_2121,_w_2129,n210_0,_w_2130,n437,_w_2347,_w_2131,_w_2922,n824_0,_w_2132,n384_0,_w_2133,_w_2253,_w_2135,G12_14,n51_3,_w_2139,_w_2141,_w_2142,_w_2959,n385_15,_w_2145,_w_2146,_w_2148,_w_2151,n395_16,_w_2152,_w_2153,_w_2161,_w_2162,_w_2500,n374,_w_2166,n233_0,_w_2167,_w_2168,n782,n254,n494,_w_2169,_w_2937,_w_2856,_w_2170,_w_2378,_w_2315,_w_2173,G4_34,_w_2332,_w_2176,n407_0,_w_2136,_w_2180,_w_2182,_w_3302,_w_2719,_w_2184,_w_2189,_w_2195,n147_3,G8_2,_w_2149,n683_1,n119_0,_w_2201,_w_2785,n398_18,_w_2203,_w_2208,_w_3433,_w_2209,_w_3441,_w_2213,_w_3562,_w_2215,_w_3381,_w_2808,_w_2624,_w_2217,_w_2628,_w_2223,_w_3039,_w_2226,G4_28,_w_2342,_w_2230,_w_2234,_w_3081,_w_2236,n355,_w_2238,_w_3559,_w_3386,G8_13,_w_2240,_w_2241,_w_2244,n811,_w_2250,_w_2252,_w_2254,_w_2256,n382,_w_2257,_w_2258,_w_3040,_w_2259,_w_2261,_w_3209,_w_2265,_w_3124,_w_2682,n110_0,_w_2271,_w_3098,_w_2272,_w_2274,n818,_w_2275,_w_2277,_w_2279,n326,_w_2282,_w_2284,_w_2493,n794,n471,_w_2285,_w_3325,_w_2828,_w_2286,_w_2291,_w_2294,_w_2967,_w_2295,_w_2297,_w_2301,_w_2302,_w_2303,_w_2307,n361_0,_w_2308,n689,_w_2311,_w_3002,_w_2312,_w_3055,_w_2316,_w_2318,_w_2321,_w_2326,n408,_w_2329,_w_2556,_w_2337,_w_2925,_w_2338,_w_2138,_w_2339,_w_2345,_w_2352,n512,_w_2353;

  bfr _b_2756(.a(G9),.q(_w_3572));
  bfr _b_2754(.a(G7),.q(_w_3570));
  bfr _b_2753(.a(_w_3569),.q(_w_3525));
  bfr _b_2750(.a(_w_3566),.q(_w_3567));
  bfr _b_2749(.a(_w_3565),.q(_w_3566));
  bfr _b_2748(.a(_w_3564),.q(_w_3565));
  bfr _b_2746(.a(_w_3562),.q(_w_3563));
  bfr _b_2745(.a(_w_3561),.q(_w_3562));
  bfr _b_2744(.a(_w_3560),.q(_w_3561));
  bfr _b_2743(.a(_w_3559),.q(_w_3560));
  bfr _b_2742(.a(_w_3558),.q(_w_3559));
  bfr _b_2741(.a(_w_3557),.q(_w_3558));
  bfr _b_2739(.a(_w_3555),.q(_w_3556));
  bfr _b_2738(.a(_w_3554),.q(_w_3555));
  bfr _b_2735(.a(_w_3551),.q(_w_3552));
  bfr _b_2733(.a(_w_3549),.q(_w_3550));
  bfr _b_2730(.a(_w_3546),.q(_w_3547));
  bfr _b_2729(.a(_w_3545),.q(_w_3546));
  bfr _b_2727(.a(_w_3543),.q(_w_3544));
  bfr _b_2726(.a(_w_3542),.q(_w_3543));
  bfr _b_2724(.a(_w_3540),.q(_w_3541));
  bfr _b_2722(.a(_w_3538),.q(_w_3539));
  bfr _b_2721(.a(_w_3537),.q(_w_3538));
  bfr _b_2720(.a(_w_3536),.q(_w_3537));
  bfr _b_2719(.a(_w_3535),.q(_w_3536));
  bfr _b_2718(.a(_w_3534),.q(_w_3535));
  bfr _b_2717(.a(_w_3533),.q(_w_3534));
  bfr _b_2715(.a(_w_3531),.q(_w_3532));
  bfr _b_2714(.a(_w_3530),.q(_w_3531));
  bfr _b_2713(.a(_w_3529),.q(_w_3530));
  bfr _b_2712(.a(_w_3528),.q(_w_3529));
  bfr _b_2711(.a(_w_3527),.q(_w_3528));
  bfr _b_2705(.a(_w_3521),.q(_w_3522));
  bfr _b_2704(.a(_w_3520),.q(_w_3521));
  bfr _b_2703(.a(_w_3519),.q(_w_3520));
  bfr _b_2701(.a(_w_3517),.q(_w_3518));
  bfr _b_2699(.a(G48),.q(_w_3516));
  bfr _b_2697(.a(_w_3513),.q(_w_3514));
  bfr _b_2696(.a(_w_3512),.q(_w_3513));
  bfr _b_2695(.a(_w_3511),.q(_w_3512));
  bfr _b_2693(.a(_w_3509),.q(_w_3510));
  bfr _b_2692(.a(_w_3508),.q(_w_3509));
  bfr _b_2690(.a(_w_3506),.q(_w_3507));
  bfr _b_2689(.a(_w_3505),.q(_w_3506));
  bfr _b_2688(.a(_w_3504),.q(_w_3505));
  bfr _b_2687(.a(_w_3503),.q(_w_3504));
  bfr _b_2686(.a(_w_3502),.q(_w_3503));
  bfr _b_2685(.a(_w_3501),.q(_w_3502));
  bfr _b_2684(.a(_w_3500),.q(_w_3501));
  bfr _b_2682(.a(_w_3498),.q(_w_3499));
  bfr _b_2681(.a(_w_3497),.q(_w_3498));
  bfr _b_2679(.a(G47),.q(_w_3496));
  bfr _b_2674(.a(_w_3490),.q(_w_3491));
  bfr _b_2672(.a(_w_3488),.q(_w_3489));
  bfr _b_2671(.a(G44),.q(_w_3488));
  bfr _b_2670(.a(_w_3486),.q(_w_3482));
  bfr _b_2669(.a(_w_3485),.q(_w_3486));
  bfr _b_2666(.a(G43),.q(_w_3483));
  bfr _b_2665(.a(_w_3481),.q(_w_3480));
  bfr _b_2755(.a(G8),.q(_w_3571));
  bfr _b_2663(.a(_w_3479),.q(_w_3478));
  bfr _b_2662(.a(G39),.q(_w_3479));
  bfr _b_2660(.a(G38),.q(_w_3477));
  bfr _b_2659(.a(G37),.q(_w_3475));
  bfr _b_2658(.a(G36),.q(_w_3474));
  bfr _b_2657(.a(G35),.q(_w_3473));
  bfr _b_2652(.a(G30),.q(_w_3468));
  bfr _b_2648(.a(G28),.q(_w_3465));
  bfr _b_2647(.a(_w_3463),.q(_w_3455));
  bfr _b_2752(.a(_w_3568),.q(_w_3569));
  bfr _b_2645(.a(_w_3461),.q(_w_3462));
  bfr _b_2643(.a(_w_3459),.q(_w_3460));
  bfr _b_2636(.a(_w_3452),.q(_w_3446));
  bfr _b_2635(.a(_w_3451),.q(_w_3452));
  bfr _b_2634(.a(_w_3450),.q(_w_3451));
  bfr _b_2633(.a(_w_3449),.q(_w_3450));
  bfr _b_2626(.a(_w_3442),.q(_w_3438));
  bfr _b_2678(.a(G46),.q(_w_3494));
  bfr _b_2625(.a(_w_3441),.q(_w_3442));
  bfr _b_2624(.a(_w_3440),.q(_w_3441));
  bfr _b_2623(.a(_w_3439),.q(_w_3440));
  bfr _b_2620(.a(_w_3436),.q(_w_3437));
  bfr _b_2619(.a(_w_3435),.q(_w_3436));
  bfr _b_2613(.a(_w_3429),.q(_w_3430));
  bfr _b_2611(.a(G18),.q(_w_3428));
  bfr _b_2610(.a(_w_3426),.q(_w_3421));
  bfr _b_2606(.a(_w_3422),.q(_w_3423));
  bfr _b_2605(.a(G17),.q(_w_3422));
  bfr _b_2602(.a(_w_3418),.q(_w_3419));
  bfr _b_2600(.a(_w_3416),.q(_w_3417));
  bfr _b_2599(.a(_w_3415),.q(_w_3416));
  bfr _b_2598(.a(_w_3414),.q(_w_3415));
  bfr _b_2596(.a(G15),.q(_w_3412));
  bfr _b_2593(.a(G12),.q(_w_3409));
  bfr _b_2592(.a(G11),.q(_w_3408));
  bfr _b_2591(.a(G10),.q(_w_3407));
  bfr _b_2589(.a(_w_3405),.q(_w_3406));
  bfr _b_2588(.a(_w_3404),.q(_w_3405));
  bfr _b_2584(.a(_w_3400),.q(_w_3401));
  bfr _b_2583(.a(_w_3399),.q(n275_1));
  bfr _b_2579(.a(_w_3395),.q(n361_16));
  bfr _b_2577(.a(_w_3393),.q(n472));
  bfr _b_2573(.a(_w_3389),.q(_w_3390));
  bfr _b_2568(.a(_w_3384),.q(_w_3385));
  bfr _b_2567(.a(_w_3383),.q(_w_3384));
  bfr _b_2563(.a(_w_3379),.q(_w_3380));
  bfr _b_2561(.a(_w_3377),.q(_w_3378));
  bfr _b_2560(.a(_w_3376),.q(_w_3377));
  bfr _b_2558(.a(_w_3374),.q(_w_3375));
  bfr _b_2557(.a(_w_3373),.q(_w_3374));
  bfr _b_2555(.a(_w_3371),.q(_w_3372));
  bfr _b_2554(.a(_w_3370),.q(_w_3371));
  bfr _b_2553(.a(_w_3369),.q(_w_3370));
  bfr _b_2552(.a(_w_3368),.q(_w_3369));
  bfr _b_2550(.a(_w_3366),.q(G43_1));
  bfr _b_2547(.a(_w_3363),.q(_w_3364));
  bfr _b_2580(.a(_w_3396),.q(_w_3397));
  bfr _b_2546(.a(_w_3362),.q(_w_3363));
  bfr _b_2543(.a(_w_3359),.q(G21_9));
  bfr _b_2542(.a(_w_3358),.q(G3528));
  bfr _b_2541(.a(_w_3357),.q(_w_3358));
  bfr _b_2539(.a(_w_3355),.q(_w_3356));
  bfr _b_2537(.a(_w_3353),.q(_w_3354));
  bfr _b_2536(.a(_w_3352),.q(_w_3353));
  bfr _b_2535(.a(_w_3351),.q(_w_3352));
  bfr _b_2534(.a(_w_3350),.q(_w_3351));
  bfr _b_2531(.a(_w_3347),.q(G10_2));
  bfr _b_2529(.a(_w_3345),.q(_w_3346));
  bfr _b_2525(.a(_w_3341),.q(G2_2));
  bfr _b_2522(.a(_w_3338),.q(_w_3339));
  bfr _b_2521(.a(_w_3337),.q(_w_3338));
  bfr _b_2520(.a(_w_3336),.q(_w_3337));
  bfr _b_2518(.a(_w_3334),.q(_w_3335));
  bfr _b_2513(.a(_w_3329),.q(G1_11));
  bfr _b_2511(.a(_w_3327),.q(G1_6));
  bfr _b_2510(.a(_w_3326),.q(G32_7));
  bfr _b_2509(.a(_w_3325),.q(_w_3326));
  bfr _b_2508(.a(_w_3324),.q(_w_3325));
  bfr _b_2507(.a(_w_3323),.q(G5_2));
  bfr _b_2506(.a(_w_3322),.q(G48_1));
  bfr _b_2504(.a(_w_3320),.q(_w_3321));
  bfr _b_2503(.a(_w_3319),.q(_w_3320));
  bfr _b_2501(.a(_w_3317),.q(_w_3318));
  bfr _b_2500(.a(_w_3316),.q(_w_3317));
  bfr _b_2499(.a(_w_3315),.q(_w_3316));
  bfr _b_2497(.a(_w_3313),.q(_w_3314));
  bfr _b_2494(.a(_w_3310),.q(_w_3311));
  bfr _b_2649(.a(_w_3465),.q(_w_3466));
  bfr _b_2493(.a(_w_3309),.q(_w_3310));
  bfr _b_2492(.a(_w_3308),.q(_w_3309));
  bfr _b_2489(.a(_w_3305),.q(_w_3306));
  bfr _b_2488(.a(_w_3304),.q(_w_3305));
  bfr _b_2486(.a(_w_3302),.q(_w_3303));
  bfr _b_2485(.a(_w_3301),.q(_w_3302));
  bfr _b_2484(.a(_w_3300),.q(_w_3301));
  bfr _b_2483(.a(_w_3299),.q(_w_3300));
  bfr _b_2480(.a(_w_3296),.q(_w_3297));
  bfr _b_2478(.a(_w_3294),.q(_w_3295));
  bfr _b_2477(.a(_w_3293),.q(_w_3294));
  bfr _b_2475(.a(_w_3291),.q(_w_3292));
  bfr _b_2471(.a(_w_3287),.q(_w_3288));
  bfr _b_2470(.a(_w_3286),.q(G41_3));
  bfr _b_2468(.a(_w_3284),.q(_w_3285));
  bfr _b_2462(.a(_w_3278),.q(G3533));
  bfr _b_2461(.a(_w_3277),.q(_w_3278));
  bfr _b_2559(.a(_w_3375),.q(_w_3376));
  bfr _b_2459(.a(_w_3275),.q(_w_3276));
  bfr _b_2458(.a(_w_3274),.q(_w_3275));
  bfr _b_2457(.a(_w_3273),.q(_w_3274));
  bfr _b_2453(.a(_w_3269),.q(_w_3270));
  bfr _b_2452(.a(_w_3268),.q(_w_3269));
  bfr _b_2451(.a(_w_3267),.q(G34_8));
  bfr _b_2449(.a(_w_3265),.q(G36_5));
  bfr _b_2448(.a(_w_3264),.q(n240));
  bfr _b_2447(.a(_w_3263),.q(_w_3264));
  bfr _b_2444(.a(_w_3260),.q(_w_3261));
  bfr _b_2443(.a(_w_3259),.q(G31_5));
  bfr _b_2442(.a(_w_3258),.q(G3_6));
  bfr _b_2440(.a(_w_3256),.q(n176_3));
  bfr _b_2439(.a(_w_3255),.q(n75_1));
  bfr _b_2438(.a(_w_3254),.q(_w_3255));
  bfr _b_2437(.a(_w_3253),.q(_w_3254));
  bfr _b_2436(.a(_w_3252),.q(_w_3253));
  bfr _b_2429(.a(_w_3245),.q(_w_3246));
  bfr _b_2426(.a(_w_3242),.q(_w_3243));
  bfr _b_2424(.a(_w_3240),.q(_w_3241));
  bfr _b_2422(.a(_w_3238),.q(_w_3239));
  bfr _b_2421(.a(_w_3237),.q(_w_3238));
  bfr _b_2419(.a(_w_3235),.q(_w_3236));
  bfr _b_2425(.a(_w_3241),.q(_w_3242));
  bfr _b_2418(.a(_w_3234),.q(_w_3235));
  bfr _b_2416(.a(_w_3232),.q(_w_3233));
  bfr _b_2415(.a(_w_3231),.q(G14_19));
  bfr _b_2413(.a(_w_3229),.q(_w_3230));
  bfr _b_2412(.a(_w_3228),.q(_w_3229));
  bfr _b_2408(.a(_w_3224),.q(n581_1));
  bfr _b_2407(.a(_w_3223),.q(G17_3));
  bfr _b_2405(.a(_w_3221),.q(G16_1));
  bfr _b_2403(.a(_w_3219),.q(_w_3220));
  bfr _b_2533(.a(_w_3349),.q(_w_3350));
  bfr _b_2402(.a(_w_3218),.q(G1_9));
  bfr _b_2540(.a(_w_3356),.q(_w_3357));
  bfr _b_2399(.a(_w_3215),.q(G4_35));
  bfr _b_2395(.a(_w_3211),.q(G4_6));
  bfr _b_2394(.a(_w_3210),.q(G4_5));
  bfr _b_2393(.a(_w_3209),.q(G3529_0));
  bfr _b_2392(.a(_w_3208),.q(_w_3209));
  bfr _b_2391(.a(_w_3207),.q(_w_3208));
  bfr _b_2389(.a(_w_3205),.q(_w_3206));
  bfr _b_2388(.a(_w_3204),.q(_w_3205));
  bfr _b_2571(.a(_w_3387),.q(_w_3388));
  bfr _b_2387(.a(_w_3203),.q(_w_3204));
  bfr _b_2386(.a(_w_3202),.q(n129_3));
  bfr _b_2384(.a(_w_3200),.q(_w_3201));
  bfr _b_2383(.a(_w_3199),.q(n542_1));
  bfr _b_2382(.a(_w_3198),.q(_w_3199));
  bfr _b_2381(.a(_w_3197),.q(_w_3198));
  bfr _b_2380(.a(_w_3196),.q(n137_6));
  bfr _b_2379(.a(_w_3195),.q(_w_3196));
  bfr _b_2378(.a(_w_3194),.q(_w_3195));
  bfr _b_2374(.a(_w_3190),.q(G3536_2));
  bfr _b_2372(.a(_w_3188),.q(n263));
  bfr _b_2371(.a(_w_3187),.q(n240_1));
  bfr _b_2370(.a(_w_3186),.q(G37_3));
  bfr _b_2367(.a(_w_3183),.q(n501_2));
  bfr _b_2365(.a(_w_3181),.q(_w_3182));
  bfr _b_2364(.a(_w_3180),.q(_w_3181));
  bfr _b_2362(.a(_w_3178),.q(_w_3179));
  bfr _b_2360(.a(_w_3176),.q(_w_3177));
  bfr _b_2411(.a(_w_3227),.q(G23_1));
  bfr _b_2359(.a(_w_3175),.q(_w_3176));
  bfr _b_2357(.a(_w_3173),.q(n123_10));
  and_bi g500(.a(n498),.b(n499),.q(n500));
  bfr _b_1398(.a(_w_2214),.q(_w_2215));
  bfr _b_1865(.a(_w_2681),.q(_w_2682));
  bfr _b_2396(.a(_w_3212),.q(_w_3213));
  spl2 g361_s_5(.a(n361_14),.q0(n361_15),.q1(_w_3395));
  bfr _b_2210(.a(_w_3026),.q(_w_3027));
  spl2 g361_s_4(.a(n361_12),.q0(n361_13),.q1(n361_14));
  spl2 g145_s_2(.a(n145_4),.q0(n145_5),.q1(n145_6));
  spl3L g145_s_0(.a(n145),.q0(n145_0),.q1(n145_1),.q2(n145_2));
  spl2 g371_s_1(.a(G3526_2),.q0(G3526_3),.q1(_w_3368));
  bfr _b_1710(.a(_w_2526),.q(n580));
  spl2 G2_s_3(.a(G2_6),.q0(G2_7),.q1(G2_8));
  and_bb g655(.a(G22_7),.b(n395_10),.q(n655));
  spl2 G2_s_1(.a(G2_2),.q0(G2_3),.q1(G2_4));
  and_bi g316(.a(n162_10),.b(n315_2),.q(n316));
  spl2 G39_s_3(.a(G39_7),.q0(G39_8),.q1(G39_9));
  spl2 G43_s_0(.a(_w_3482),.q0(G43_0),.q1(_w_3366));
  spl2 G21_s_3(.a(G21_7),.q0(G21_8),.q1(_w_3359));
  bfr _b_1536(.a(_w_2352),.q(_w_2353));
  spl2 g603_s_0(.a(G3531_0),.q0(G3531_1),.q1(G3531_2));
  spl4L G10_s_2(.a(G10_4),.q0(G10_5),.q1(G10_6),.q2(G10_7),.q3(G10_8));
  spl2 g315_s_0(.a(n315),.q0(n315_0),.q1(n315_1));
  spl2 g641_s_0(.a(G3532_0),.q0(G3532_1),.q1(G3532_2));
  spl2 g321_s_0(.a(n321),.q0(n321_0),.q1(n321_1));
  bfr _b_2548(.a(_w_3364),.q(_w_3365));
  bfr _b_2187(.a(_w_3003),.q(_w_3004));
  spl2 g113_s_0(.a(n113),.q0(n113_0),.q1(n113_1));
  spl3L G2_s_0(.a(G2),.q0(G2_0),.q1(G2_1),.q2(_w_3334));
  spl4L g369_s_0(.a(n369),.q0(n369_0),.q1(n369_1),.q2(n369_2),.q3(_w_3330));
  bfr _b_1739(.a(_w_2555),.q(_w_2556));
  spl3L G1_s_1(.a(G1_3),.q0(G1_4),.q1(G1_5),.q2(_w_3327));
  and_bi g268(.a(n143_3),.b(n265_5),.q(n268));
  spl2 g490_s_2(.a(n490_4),.q0(n490_5),.q1(n490_6));
  spl2 G32_s_2(.a(G32_5),.q0(G32_6),.q1(_w_3324));
  spl3L G5_s_0(.a(G5),.q0(G5_0),.q1(G5_1),.q2(_w_3323));
  spl4L g398_s_3(.a(n398_7),.q0(n398_12),.q1(n398_13),.q2(n398_14),.q3(n398_15));
  spl2 G48_s_0(.a(_w_3515),.q0(G48_0),.q1(_w_3289));
  bfr _b_2630(.a(G23),.q(_w_3447));
  and_bi g138(.a(n137_0),.b(G8_6),.q(n138));
  bfr _b_2291(.a(_w_3107),.q(n604_2));
  spl2 g126_s_1(.a(n126_1),.q0(n126_2),.q1(_w_3287));
  bfr _b_1535(.a(_w_2351),.q(_w_2352));
  spl2 g623_s_0(.a(n623),.q0(n623_0),.q1(_w_3283));
  bfr _b_2127(.a(_w_2943),.q(_w_2944));
  spl4L g395_s_2(.a(n395_6),.q0(n395_8),.q1(n395_9),.q2(n395_10),.q3(n395_11));
  bfr _b_1400(.a(_w_2216),.q(_w_2217));
  spl3L g190_s_0(.a(n190),.q0(n190_0),.q1(n190_1),.q2(n190_2));
  bfr _b_2487(.a(_w_3303),.q(_w_3304));
  and_bb g660(.a(G42_4),.b(n395_5),.q(n660));
  and_bi g324(.a(n123_9),.b(G14_8),.q(n324));
  spl2 G39_s_4(.a(G39_9),.q0(G39_10),.q1(G39_11));
  bfr _b_1659(.a(_w_2475),.q(_w_2476));
  spl2 g107_s_0(.a(n107),.q0(n107_0),.q1(n107_1));
  bfr _b_2204(.a(_w_3020),.q(_w_3021));
  spl3L G41_s_2(.a(G41_3),.q0(G41_4),.q1(G41_5),.q2(_w_3279));
  and_bb g497(.a(n176_3),.b(n496_0),.q(n497));
  spl2 G34_s_2(.a(G34_6),.q0(G34_7),.q1(_w_3266));
  spl2 G36_s_1(.a(G36_3),.q0(G36_4),.q1(_w_3265));
  and_bb g240(.a(n191_0),.b(n239),.q(_w_3262));
  spl2 g692_s_0(.a(n692),.q0(n692_0),.q1(n692_1));
  bfr _b_2377(.a(_w_3193),.q(_w_3194));
  bfr _b_2347(.a(_w_3163),.q(n214_2));
  spl2 g489_s_0(.a(G3529_0),.q0(G3529_1),.q1(_w_3260));
  spl2 G31_s_1(.a(G31_3),.q0(G31_4),.q1(_w_3259));
  bfr _b_2463(.a(_w_3279),.q(_w_3280));
  bfr _b_2076(.a(_w_2892),.q(n513));
  spl4L G3_s_5(.a(G3_13),.q0(G3_14),.q1(G3_15),.q2(G3_16),.q3(G3_17));
  and_bi g80(.a(n79),.b(n77_0),.q(n80));
  bfr _b_2015(.a(_w_2831),.q(_w_2832));
  spl4L g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1),.q2(n361_2),.q3(n361_3));
  spl4L G3_s_2(.a(G3_3),.q0(G3_4),.q1(G3_5),.q2(_w_3258),.q3(G3_7));
  spl2 G3_s_1(.a(G3_1),.q0(G3_2),.q1(G3_3));
  bfr _b_1666(.a(_w_2482),.q(_w_2483));
  and_bb g131(.a(G7_8),.b(n130_0),.q(n131));
  bfr _b_2297(.a(_w_3113),.q(n775));
  spl2 G26_s_0(.a(_w_3454),.q0(G26_0),.q1(G26_1));
  and_bb g783(.a(G10_7),.b(G14_10),.q(n783));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(_w_3232));
  bfr _b_2193(.a(_w_3009),.q(_w_3010));
  bfr _b_1787(.a(_w_2603),.q(_w_2604));
  or_bb g315(.a(n284_1),.b(n314_0),.q(n315));
  spl2 g91_s_0(.a(n91),.q0(n91_0),.q1(n91_1));
  and_bb g295(.a(n282_0),.b(n294),.q(n295));
  spl2 G20_s_2(.a(G20_4),.q0(G20_5),.q1(_w_3226));
  bfr _b_1736(.a(_w_2552),.q(_w_2553));
  spl4L G32_s_0(.a(_w_3470),.q0(G32_0),.q1(G32_1),.q2(G32_2),.q3(G32_3));
  bfr _b_2616(.a(G20),.q(_w_3433));
  spl2 G20_s_0(.a(_w_3432),.q0(G20_0),.q1(G20_1));
  bfr _b_1952(.a(_w_2768),.q(_w_2769));
  spl4L G9_s_4(.a(G9_8),.q0(G9_9),.q1(G9_10),.q2(G9_11),.q3(G9_12));
  spl2 g824_s_0(.a(n824),.q0(n824_0),.q1(n824_1));
  bfr _b_1381(.a(_w_2197),.q(_w_2198));
  spl2 G9_s_2(.a(G9_3),.q0(G9_4),.q1(_w_3225));
  spl2 g428_s_1(.a(n428_1),.q0(n428_2),.q1(n428_3));
  spl2 g581_s_0(.a(n581),.q0(n581_0),.q1(_w_3224));
  and_bi g211(.a(n143_10),.b(n210_1),.q(n211));
  spl2 g546_s_1(.a(n546_1),.q0(n546_2),.q1(n546_3));
  spl2 G13_s_1(.a(G13_1),.q0(G13_2),.q1(G13_3));
  and_bb g474(.a(G24_7),.b(n265_2),.q(n474));
  and_bb g501(.a(n495_0),.b(n500_5),.q(n501));
  bfr _b_1595(.a(_w_2411),.q(G3525));
  spl3L G1_s_2(.a(G1_6),.q0(G1_7),.q1(G1_8),.q2(_w_3216));
  spl4L G4_s_13(.a(G4_42),.q0(G4_45),.q1(G4_46),.q2(G4_47),.q3(G4_48));
  spl4L G4_s_9(.a(G4_31),.q0(G4_32),.q1(G4_33),.q2(G4_34),.q3(_w_3215));
  spl2 g654_s_0(.a(n654),.q0(n654_0),.q1(n654_1));
  spl4L G4_s_7(.a(G4_22),.q0(G4_25),.q1(G4_26),.q2(G4_27),.q3(G4_28));
  bfr _b_2198(.a(_w_3014),.q(_w_3015));
  spl4L G4_s_1(.a(G4_2),.q0(G4_4),.q1(_w_3210),.q2(_w_3211),.q3(G4_7));
  bfr _b_2590(.a(_w_3406),.q(n509_1));
  and_bb g355(.a(n191_1),.b(n354),.q(n355));
  bfr _b_2257(.a(_w_3073),.q(_w_3074));
  and_bb g612(.a(G43_2),.b(n395_4),.q(n612));
  spl2 G11_s_5(.a(G11_12),.q0(G11_13),.q1(G11_14));
  or_bb g489(.a(n468),.b(n488),.q(_w_3203));
  bfr _b_2629(.a(_w_3445),.q(_w_3443));
  bfr _b_2132(.a(_w_2948),.q(_w_2949));
  spl2 G33_s_1(.a(G33_3),.q0(G33_4),.q1(G33_5));
  bfr _b_2465(.a(_w_3281),.q(_w_3282));
  or_bb g698(.a(n372_10),.b(n697_0),.q(n698));
  bfr _b_1777(.a(_w_2593),.q(_w_2594));
  and_bi g781(.a(G40_6),.b(n398_12),.q(n781));
  spl4L G14_s_4(.a(G14_7),.q0(G14_8),.q1(G14_9),.q2(G14_10),.q3(G14_11));
  bfr _b_1708(.a(_w_2524),.q(n381));
  bfr _b_1738(.a(_w_2554),.q(_w_2555));
  spl2 g814_s_0(.a(n814),.q0(n814_0),.q1(n814_1));
  bfr _b_1422(.a(_w_2238),.q(G3534));
  spl2 g394_s_0(.a(n394),.q0(n394_0),.q1(n394_1));
  spl4L g129_s_0(.a(n129),.q0(n129_0),.q1(n129_1),.q2(n129_2),.q3(_w_3202));
  spl2 G13_s_0(.a(_w_3410),.q0(G13_0),.q1(G13_1));
  and_bi g153(.a(G10_1),.b(G4_4),.q(n153));
  and_bb g348(.a(n269_1),.b(n295_1),.q(n348));
  bfr _b_2680(.a(_w_3496),.q(_w_3497));
  bfr _b_1731(.a(_w_2547),.q(_w_2548));
  spl2 g542_s_0(.a(n542),.q0(n542_0),.q1(_w_3197));
  spl2 g553_s_1(.a(n553_1),.q0(n553_2),.q1(n553_3));
  and_bi g270(.a(n269_0),.b(n267_0),.q(n270));
  spl2 g337_s_0(.a(n337),.q0(n337_0),.q1(n337_1));
  spl2 g110_s_0(.a(n110),.q0(n110_0),.q1(n110_1));
  spl2 g240_s_1(.a(n240_1),.q0(n240_2),.q1(_w_3191));
  spl4L g147_s_2(.a(n147_5),.q0(n147_6),.q1(n147_7),.q2(n147_8),.q3(n147_9));
  spl2 g810_s_0(.a(G3536_0),.q0(G3536_1),.q1(_w_3189));
  bfr _b_1481(.a(_w_2297),.q(_w_2298));
  spl4L G37_s_0(.a(_w_3475),.q0(G37_0),.q1(G37_1),.q2(G37_2),.q3(_w_3184));
  spl2 g419_s_0(.a(n419),.q0(n419_0),.q1(n419_1));
  bfr _b_2473(.a(_w_3289),.q(_w_3290));
  bfr _b_1800(.a(_w_2616),.q(_w_2617));
  spl3L g501_s_0(.a(n501),.q0(n501_0),.q1(n501_1),.q2(_w_3183));
  bfr _b_2068(.a(_w_2884),.q(_w_2885));
  spl2 g777_s_1(.a(G3535_2),.q0(G3535_3),.q1(_w_3174));
  spl2 g777_s_0(.a(G3535_0),.q0(G3535_1),.q1(G3535_2));
  bfr _b_1493(.a(_w_2309),.q(_w_2310));
  spl4L g123_s_3(.a(n123_3),.q0(n123_7),.q1(n123_8),.q2(n123_9),.q3(_w_3173));
  bfr _b_2045(.a(_w_2861),.q(_w_2862));
  and_bi g428(.a(G47_0),.b(n369_1),.q(n428));
  or_bb g471(.a(n469),.b(n470),.q(n471));
  spl3L G12_s_5(.a(G12_12),.q0(G12_13),.q1(G12_14),.q2(G12_15));
  spl2 G31_s_2(.a(G31_5),.q0(G31_6),.q1(_w_3172));
  spl2 G12_s_3(.a(G12_6),.q0(G12_7),.q1(_w_3170));
  spl2 G12_s_2(.a(G12_4),.q0(G12_5),.q1(G12_6));
  spl4L G4_s_2(.a(G4_3),.q0(_w_3169),.q1(G4_9),.q2(G4_10),.q3(G4_11));
  bfr _b_1848(.a(_w_2664),.q(_w_2665));
  spl2 G36_s_2(.a(G36_5),.q0(G36_6),.q1(G36_7));
  spl2 G1_s_3(.a(G1_9),.q0(G1_10),.q1(_w_3328));
  spl4L g129_s_2(.a(n129_5),.q0(n129_6),.q1(n129_7),.q2(n129_8),.q3(n129_9));
  spl2 G9_s_0(.a(_w_3572),.q0(G9_0),.q1(G9_1));
  spl2 g361_s_7(.a(n361_18),.q0(n361_19),.q1(n361_20));
  spl2 G35_s_1(.a(G35_3),.q0(G35_4),.q1(G35_5));
  spl3L g343_s_0(.a(n343),.q0(n343_0),.q1(n343_1),.q2(_w_3164));
  spl3L g214_s_0(.a(n214),.q0(n214_0),.q1(n214_1),.q2(_w_3161));
  spl3L g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1),.q2(n165_2));
  spl2 g171_s_0(.a(n171),.q0(n171_0),.q1(_w_3157));
  spl2 G14_s_0(.a(_w_3411),.q0(G14_0),.q1(G14_1));
  spl3L G47_s_1(.a(G47_2),.q0(G47_3),.q1(G47_4),.q2(G47_5));
  spl3L G47_s_0(.a(_w_3495),.q0(G47_0),.q1(G47_1),.q2(_w_3154));
  bfr _b_2184(.a(_w_3000),.q(_w_3001));
  spl2 g201_s_0(.a(n201),.q0(n201_0),.q1(n201_1));
  spl3L g554_s_0(.a(n554),.q0(n554_0),.q1(n554_1),.q2(n554_2));
  spl2 g505_s_0(.a(n505),.q0(n505_0),.q1(n505_1));
  and_bi g371(.a(n370),.b(n365_2),.q(G3526_0));
  spl2 g533_s_0(.a(n533),.q0(n533_0),.q1(_w_3151));
  spl2 g534_s_0(.a(n534),.q0(n534_0),.q1(n534_1));
  bfr _b_1679(.a(_w_2495),.q(_w_2496));
  bfr _b_1793(.a(_w_2609),.q(n51_3));
  bfr _b_1849(.a(_w_2665),.q(_w_2666));
  bfr _b_2476(.a(_w_3292),.q(_w_3293));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(n235_1));
  spl2 g329_s_1(.a(n329_1),.q0(n329_2),.q1(_w_3149));
  spl3L g629_s_0(.a(n629),.q0(n629_0),.q1(n629_1),.q2(n629_2));
  spl2 g484_s_0(.a(n484),.q0(n484_0),.q1(n484_1));
  and_bi g822(.a(n812_1),.b(n821),.q(n822));
  spl2 g533_s_3(.a(n533_6),.q0(n533_7),.q1(n533_8));
  spl4L g361_s_1(.a(n361_3),.q0(n361_4),.q1(n361_5),.q2(n361_6),.q3(n361_7));
  spl2 g559_s_0(.a(n559),.q0(n559_0),.q1(n559_1));
  spl2 g495_s_0(.a(n495),.q0(n495_0),.q1(_w_3147));
  bfr _b_2549(.a(_w_3365),.q(G3537));
  bfr _b_2307(.a(_w_3123),.q(_w_3124));
  spl2 g735_s_1(.a(n735_1),.q0(n735_2),.q1(n735_3));
  spl2 g735_s_0(.a(n735),.q0(n735_0),.q1(_w_3140));
  spl4L g832_s_0(.a(n832),.q0(n832_0),.q1(n832_1),.q2(n832_2),.q3(n832_3));
  and_bi g749(.a(n748),.b(n741),.q(n749));
  bfr _b_2516(.a(_w_3332),.q(_w_3333));
  bfr _b_2135(.a(_w_2951),.q(_w_2952));
  spl3L G9_s_6(.a(G9_14),.q0(G9_15),.q1(G9_16),.q2(G9_17));
  spl4L G4_s_11(.a(G4_38),.q0(G4_39),.q1(G4_40),.q2(G4_41),.q3(G4_42));
  spl2 g627_s_0(.a(n627),.q0(n627_0),.q1(n627_1));
  spl2 g688_s_0(.a(n688),.q0(n688_0),.q1(_w_3137));
  bfr _b_1650(.a(_w_2466),.q(_w_2467));
  spl2 g838_s_0(.a(n838),.q0(n838_0),.q1(n838_1));
  bfr _b_2526(.a(_w_3342),.q(_w_3343));
  spl2 g737_s_0(.a(n737),.q0(n737_0),.q1(_w_3134));
  and_bi g132(.a(n124),.b(n131),.q(n132));
  bfr _b_1581(.a(_w_2397),.q(_w_2398));
  bfr _b_2094(.a(_w_2910),.q(_w_2911));
  spl2 g829_s_0(.a(n829),.q0(n829_0),.q1(n829_1));
  and_bi g844(.a(n842),.b(n843),.q(G3540));
  bfr _b_1671(.a(_w_2487),.q(_w_2488));
  bfr _b_2240(.a(_w_3056),.q(_w_3057));
  and_bb g843(.a(n832_3),.b(n834_5),.q(n843));
  bfr _b_1504(.a(_w_2320),.q(n546));
  or_bb g842(.a(n832_2),.b(n834_4),.q(n842));
  or_bb g113(.a(n111),.b(n112),.q(n113));
  and_bi g838(.a(n837),.b(n835),.q(n838));
  and_bi g505(.a(n490_5),.b(n504),.q(n505));
  bfr _b_1431(.a(_w_2247),.q(_w_2248));
  bfr _b_1585(.a(_w_2401),.q(_w_2402));
  and_bb g102(.a(n100_1),.b(n91_1),.q(n102));
  and_bi g245(.a(n243),.b(n244),.q(n245));
  and_bi g837(.a(n836),.b(n360_1),.q(n837));
  and_bb g833(.a(G3534_3),.b(G3535_3),.q(n833));
  spl2 G8_s_2(.a(G8_3),.q0(G8_4),.q1(_w_3132));
  and_bi g826(.a(n813_0),.b(n825),.q(n826));
  bfr _b_2532(.a(_w_3348),.q(_w_3349));
  bfr _b_2157(.a(_w_2973),.q(G3527));
  and_bb g825(.a(G3531_3),.b(G3533_3),.q(n825));
  or_bb g787(.a(G12_18),.b(n407_10),.q(n787));
  and_bb g821(.a(G3529_3),.b(G3536_3),.q(n821));
  and_bi g199(.a(n129_7),.b(n198),.q(n199));
  spl3L g162_s_3(.a(n162_7),.q0(n162_8),.q1(n162_9),.q2(n162_10));
  or_bi g820(.a(n818),.b(n819),.q(_w_3128));
  bfr _b_2650(.a(_w_3466),.q(_w_3464));
  and_bi g228(.a(G4_29),.b(G31_6),.q(n228));
  spl2 g566_s_0(.a(n566),.q0(n566_0),.q1(n566_1));
  and_bi g819(.a(G27_3),.b(G3537_1),.q(n819));
  bfr _b_1894(.a(_w_2710),.q(_w_2711));
  or_bi g817(.a(n811_0),.b(n816),.q(G3537_0));
  or_bb g810(.a(n778),.b(n809),.q(G3536_0));
  and_bi g807(.a(n806),.b(n779),.q(_w_3115));
  or_bb g804(.a(n791),.b(n803),.q(n804));
  and_bi g803(.a(n802),.b(n795),.q(n803));
  and_bb g828(.a(n824_1),.b(n826_1),.q(n828));
  or_bb g259(.a(n255),.b(n258),.q(n259));
  or_bb g797(.a(n171_1),.b(n796),.q(n797));
  spl3L G21_s_1(.a(G21_1),.q0(G21_2),.q1(G21_3),.q2(G21_4));
  and_bi g796(.a(n737_0),.b(n398_4),.q(n796));
  bfr _b_2084(.a(_w_2900),.q(_w_2901));
  or_bb g795(.a(n792),.b(n794),.q(n795));
  or_bb g794(.a(n631_1),.b(n793),.q(n794));
  and_bi g792(.a(G17_3),.b(n401_21),.q(n792));
  or_bb g470(.a(G24_6),.b(n265_0),.q(n470));
  spl2 G8_s_3(.a(G8_5),.q0(G8_6),.q1(G8_7));
  and_bb g790(.a(n787),.b(n789),.q(n790));
  bfr _b_1537(.a(_w_2353),.q(_w_2354));
  bfr _b_1690(.a(_w_2506),.q(n209));
  or_bb g788(.a(n401_12),.b(n669_1),.q(n788));
  and_bi g786(.a(n785),.b(n782),.q(n786));
  bfr _b_2247(.a(_w_3063),.q(_w_3064));
  and_bi g785(.a(n784),.b(n630_1),.q(n785));
  or_bb g782(.a(n780),.b(n781),.q(n782));
  and_bb g830(.a(n822_0),.b(n829_0),.q(n830));
  spl3L G4_s_8(.a(G4_28),.q0(G4_29),.q1(G4_30),.q2(G4_31));
  and_bb g780(.a(G39_8),.b(n395_12),.q(n780));
  and_bb g779(.a(n437_4),.b(n494_1),.q(n779));
  bfr _b_2345(.a(_w_3161),.q(_w_3162));
  and_bi g776(.a(n775),.b(n769),.q(n776));
  bfr _b_2466(.a(_w_3282),.q(G39_1));
  or_bb g772(.a(n770),.b(n771),.q(n772));
  bfr _b_2165(.a(_w_2981),.q(_w_2982));
  spl3L G34_s_1(.a(G34_3),.q0(G34_4),.q1(G34_5),.q2(G34_6));
  and_bi g771(.a(n735_3),.b(n514_1),.q(n771));
  spl2 g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1));
  and_bi g770(.a(n514_0),.b(n735_2),.q(n770));
  spl4L G11_s_4(.a(G11_8),.q0(G11_9),.q1(G11_10),.q2(G11_11),.q3(G11_12));
  and_bi g766(.a(n696_2),.b(n688_0),.q(n766));
  spl3L g604_s_0(.a(n604),.q0(n604_0),.q1(n604_1),.q2(_w_3107));
  bfr _b_2329(.a(_w_3145),.q(_w_3146));
  spl3L G11_s_3(.a(G11_5),.q0(G11_6),.q1(_w_3106),.q2(G11_8));
  and_bb g765(.a(n695_1),.b(n696_1),.q(n765));
  and_bi g764(.a(n763),.b(n736),.q(_w_3088));
  and_bb g759(.a(n756),.b(n758),.q(n759));
  bfr _b_1579(.a(_w_2395),.q(_w_2396));
  and_bb g758(.a(n629_1),.b(n757),.q(n758));
  and_bi g755(.a(n623_0),.b(n754),.q(n755));
  bfr _b_2183(.a(_w_2999),.q(n673));
  and_bi g753(.a(n752),.b(n581_0),.q(n753));
  spl2 G4_s_6(.a(G4_21),.q0(G4_23),.q1(G4_24));
  bfr _b_2482(.a(_w_3298),.q(_w_3299));
  or_bb g752(.a(G14_13),.b(n398_11),.q(n752));
  and_bb g475(.a(n293_2),.b(n474),.q(n475));
  and_bi g747(.a(n146_1),.b(n746),.q(n747));
  and_bi g818(.a(G48_1),.b(n811_2),.q(_w_3084));
  and_bi g744(.a(n743),.b(n401_1),.q(n744));
  bfr _b_1647(.a(_w_2463),.q(_w_2464));
  and_bi g740(.a(G20_5),.b(n407_1),.q(n740));
  bfr _b_1601(.a(_w_2417),.q(n354));
  spl2 g201_s_1(.a(n201_1),.q0(n201_2),.q1(_w_3078));
  and_bi g735(.a(n733),.b(n734),.q(n735));
  and_bb g734(.a(n165_2),.b(n732_1),.q(n734));
  bfr _b_1298(.a(_w_2114),.q(_w_2115));
  bfr _b_1818(.a(_w_2634),.q(n358_1));
  or_bb g733(.a(n165_1),.b(n732_0),.q(n733));
  and_bb g732(.a(n142_2),.b(n496_1),.q(n732));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  and_bi g719(.a(G21_8),.b(n407_0),.q(_w_3077));
  bfr _b_2569(.a(_w_3385),.q(_w_3386));
  bfr _b_1295(.a(_w_2111),.q(_w_2112));
  or_bb g726(.a(n713),.b(n725),.q(n726));
  or_bb g641(.a(n605),.b(n640),.q(_w_3070));
  bfr _b_2433(.a(_w_3249),.q(_w_3250));
  and_bi g725(.a(n724),.b(n718),.q(n725));
  and_bb g720(.a(G18_2),.b(n395_8),.q(n720));
  and_bb g716(.a(G22_8),.b(n392_13),.q(n716));
  spl2 G25_s_0(.a(_w_3453),.q0(G25_0),.q1(_w_3069));
  spl2 g399_s_0(.a(n399),.q0(n399_0),.q1(_w_3068));
  or_bb g737(.a(G18_0),.b(G22_2),.q(n737));
  bfr _b_2640(.a(_w_3456),.q(_w_3457));
  and_bb g115(.a(G12_17),.b(G14_16),.q(n115));
  and_bb g106(.a(G10_13),.b(G7_16),.q(n106));
  and_bi g707(.a(n411_1),.b(n654_1),.q(n707));
  and_bi g605(.a(n604_0),.b(n542_0),.q(n605));
  spl2 G41_s_3(.a(G41_6),.q0(G41_7),.q1(G41_8));
  bfr _b_2661(.a(_w_3477),.q(_w_3476));
  spl2 g151_s_2(.a(n151_7),.q0(n151_8),.q1(n151_9));
  bfr _b_1496(.a(_w_2312),.q(_w_2313));
  bfr _b_2274(.a(_w_3090),.q(_w_3091));
  spl2 G9_s_1(.a(G9_1),.q0(G9_2),.q1(G9_3));
  bfr _b_1394(.a(_w_2210),.q(G22_1));
  or_bb g704(.a(n401_24),.b(n587_1),.q(n704));
  bfr _b_2020(.a(_w_2836),.q(_w_2837));
  and_bb g703(.a(n437_0),.b(n500_0),.q(n703));
  and_bi g702(.a(n701_0),.b(n688_3),.q(n702));
  spl4L G3_s_3(.a(G3_7),.q0(G3_8),.q1(G3_9),.q2(G3_10),.q3(G3_11));
  spl2 g817_s_0(.a(G3537_0),.q0(G3537_1),.q1(_w_3360));
  and_bi g339(.a(n162_6),.b(n338_0),.q(n339));
  bfr _b_1425(.a(_w_2241),.q(_w_2242));
  bfr _b_2008(.a(_w_2824),.q(_w_2825));
  and_bi g700(.a(n688_2),.b(n699),.q(_w_3067));
  spl3L g374_s_0(.a(n374),.q0(n374_0),.q1(n374_1),.q2(n374_2));
  and_bi g699(.a(n698),.b(n533_7),.q(n699));
  bfr _b_1351(.a(_w_2167),.q(_w_2168));
  bfr _b_2346(.a(_w_3162),.q(_w_3163));
  and_bi g695(.a(n693),.b(n694),.q(n695));
  or_bb g693(.a(n689_0),.b(n692_0),.q(n693));
  and_bb g647(.a(G11_13),.b(G7_13),.q(n647));
  or_bb g691(.a(n494_4),.b(n690),.q(n691));
  or_bb g689(.a(n482_1),.b(n509_1),.q(_w_3065));
  spl2 g563_s_0(.a(n563),.q0(n563_0),.q1(_w_3058));
  spl2 g361_s_6(.a(n361_16),.q0(n361_17),.q1(n361_18));
  and_bi g686(.a(n685),.b(n512_1),.q(_w_3055));
  bfr _b_1670(.a(_w_2486),.q(_w_2487));
  bfr _b_1874(.a(_w_2690),.q(_w_2691));
  spl2 g548_s_0(.a(n548),.q0(n548_0),.q1(n548_1));
  and_bb g684(.a(n490_0),.b(n495_1),.q(n684));
  bfr _b_2115(.a(_w_2931),.q(n409_1));
  and_bb g683(.a(n490_3),.b(n501_2),.q(n683));
  bfr _b_2328(.a(_w_3144),.q(_w_3145));
  or_bb g681(.a(n677),.b(n680),.q(n681));
  and_bi g773(.a(n683_1),.b(n772_0),.q(n773));
  and_bi g680(.a(n554_1),.b(n679),.q(n680));
  and_bb g596(.a(n593),.b(n595),.q(n596));
  spl2 g688_s_1(.a(n688_1),.q0(n688_2),.q1(n688_3));
  and_bb g128(.a(G4_20),.b(n127),.q(n128));
  bfr _b_1617(.a(_w_2433),.q(_w_2434));
  bfr _b_1837(.a(_w_2653),.q(_w_2654));
  and_bi g677(.a(n676),.b(n644),.q(_w_3040));
  and_ii g53(.a(n51_5),.b(n52_2),.q(_w_3000));
  and_bi g673(.a(n672),.b(n667),.q(_w_2999));
  or_bb g670(.a(n385_14),.b(n669_0),.q(n670));
  or_bb g667(.a(n663),.b(n666),.q(_w_2998));
  or_bb g666(.a(n664),.b(n665),.q(n666));
  and_bi g665(.a(n392_8),.b(G14_9),.q(n665));
  and_bi g664(.a(G43_3),.b(n398_5),.q(n664));
  or_bb g663(.a(n660),.b(n662),.q(n663));
  and_bi g662(.a(n661),.b(n401_6),.q(n662));
  and_bi g814(.a(G3528_1),.b(G3532_1),.q(n814));
  bfr _b_2104(.a(_w_2920),.q(_w_2921));
  and_bi g708(.a(n707),.b(n706),.q(n708));
  or_bb g333(.a(n331),.b(n332),.q(n333));
  and_bi g658(.a(n651),.b(n657),.q(n658));
  spl3L G20_s_1(.a(G20_1),.q0(G20_2),.q1(G20_3),.q2(G20_4));
  bfr _b_2628(.a(_w_3444),.q(_w_3445));
  and_bi g652(.a(G20_2),.b(n401_8),.q(n652));
  and_bb g543(.a(n282_3),.b(n361_1),.q(n543));
  or_bb g653(.a(G4_39),.b(n652),.q(n653));
  and_bi g645(.a(G21_9),.b(n398_21),.q(_w_2997));
  and_bi g643(.a(n642),.b(n554_2),.q(_w_2996));
  spl2 G35_s_2(.a(G35_5),.q0(G35_6),.q1(G35_7));
  and_bi g639(.a(n638),.b(n607),.q(_w_2987));
  bfr _b_2530(.a(_w_3346),.q(_w_3347));
  bfr _b_1944(.a(_w_2760),.q(_w_2761));
  or_bb g636(.a(n619),.b(n635),.q(n636));
  and_bi g557(.a(n556),.b(n533_4),.q(n557));
  bfr _b_2253(.a(_w_3069),.q(G25_1));
  spl4L g162_s_2(.a(n162_1),.q0(n162_4),.q1(n162_5),.q2(n162_6),.q3(n162_7));
  spl2 g813_s_0(.a(n813),.q0(n813_0),.q1(n813_1));
  and_bb g635(.a(n626),.b(n634),.q(n635));
  and_bi g629(.a(n628),.b(G4_40),.q(n629));
  bfr _b_2512(.a(_w_3328),.q(_w_3329));
  or_bb g627(.a(G10_15),.b(n407_8),.q(n627));
  and_bi g805(.a(n804),.b(n381_0),.q(_w_2979));
  and_bi g723(.a(n722),.b(n719),.q(n723));
  and_bi g626(.a(n625),.b(n622),.q(n626));
  bfr _b_2700(.a(_w_3516),.q(_w_3517));
  bfr _b_2639(.a(G27),.q(_w_3456));
  bfr _b_2627(.a(G22),.q(_w_3444));
  and_bb g625(.a(n623_1),.b(n624),.q(n625));
  spl2 g572_s_0(.a(n572),.q0(n572_0),.q1(n572_1));
  bfr _b_2309(.a(_w_3125),.q(_w_3126));
  and_bi g829(.a(n827),.b(n828),.q(n829));
  spl4L g398_s_0(.a(n398),.q0(n398_0),.q1(n398_1),.q2(n398_2),.q3(n398_3));
  spl2 G4_s_14(.a(G4_48),.q0(G4_49),.q1(G4_50));
  and_bb g360(.a(G27_0),.b(G48_0),.q(n360));
  or_bb g622(.a(n620),.b(n621),.q(n622));
  and_bb g746(.a(G21_3),.b(n392_1),.q(n746));
  bfr _b_2551(.a(_w_3367),.q(n147_11));
  bfr _b_1990(.a(_w_2806),.q(_w_2807));
  and_bb g617(.a(G4_44),.b(n616),.q(n617));
  bfr _b_1305(.a(_w_2121),.q(n500_5));
  or_bb g767(.a(n372_8),.b(n766),.q(n767));
  or_bb g616(.a(n385_13),.b(n460_0),.q(n616));
  and_bi g615(.a(G40_9),.b(n407_7),.q(n615));
  bfr _b_2441(.a(_w_3257),.q(G27_1));
  or_bb g614(.a(n610),.b(n613),.q(n614));
  bfr _b_2544(.a(_w_3360),.q(_w_3361));
  or_bb g305(.a(n301),.b(n304),.q(_w_2977));
  bfr _b_1642(.a(_w_2458),.q(n478));
  bfr _b_1441(.a(_w_2257),.q(_w_2258));
  and_bb g607(.a(n365_1),.b(n377_3),.q(n607));
  bfr _b_2170(.a(_w_2986),.q(n637));
  bfr _b_1859(.a(_w_2675),.q(_w_2676));
  bfr _b_2223(.a(_w_3039),.q(G3519));
  or_bb g604(.a(n374_7),.b(n540_2),.q(n604));
  and_bi g160(.a(n143_2),.b(n159_0),.q(n160));
  bfr _b_1589(.a(_w_2405),.q(_w_2406));
  bfr _b_1760(.a(_w_2576),.q(_w_2577));
  or_bb g603(.a(n570),.b(n602),.q(_w_2974));
  bfr _b_2615(.a(_w_3431),.q(_w_3427));
  and_bi g602(.a(n601),.b(n571),.q(_w_2946));
  bfr _b_1421(.a(_w_2237),.q(_w_2238));
  bfr _b_2063(.a(_w_2879),.q(G6_2));
  and_bi g252(.a(n123_7),.b(G11_9),.q(n252));
  bfr _b_2078(.a(_w_2894),.q(n812_1));
  and_bi g676(.a(n379_0),.b(n675),.q(_w_3342));
  spl2 G17_s_1(.a(G17_1),.q0(G17_2),.q1(_w_3223));
  and_bi g601(.a(n379_6),.b(n600),.q(_w_2945));
  and_bb g331(.a(G36_4),.b(G4_18),.q(n331));
  and_bi g597(.a(n596),.b(n592),.q(n597));
  spl4L g395_s_1(.a(n395_3),.q0(n395_4),.q1(n395_5),.q2(n395_6),.q3(n395_7));
  bfr _b_1387(.a(_w_2203),.q(_w_2204));
  and_bi g594(.a(n392_12),.b(G13_15),.q(n594));
  or_bb g593(.a(G14_17),.b(n407_6),.q(n593));
  bfr _b_2401(.a(_w_3217),.q(_w_3218));
  or_bb g831(.a(n822_1),.b(n829_1),.q(n831));
  and_bb g839(.a(n832_0),.b(n838_0),.q(n839));
  and_bi g609(.a(G44_2),.b(n398_8),.q(n609));
  and_bi g294(.a(n162_5),.b(n293_0),.q(n294));
  bfr _b_1870(.a(_w_2686),.q(_w_2687));
  bfr _b_2296(.a(_w_3112),.q(_w_3113));
  bfr _b_2361(.a(_w_3177),.q(_w_3178));
  or_bb g592(.a(n590),.b(n591),.q(n592));
  spl2 G38_s_0(.a(_w_3476),.q0(G38_0),.q1(_w_2943));
  bfr _b_1753(.a(_w_2569),.q(_w_2570));
  spl2 G42_s_2(.a(G42_3),.q0(G42_4),.q1(_w_2941));
  spl2 g701_s_0(.a(n701),.q0(n701_0),.q1(n701_1));
  spl2 g560_s_0(.a(n560),.q0(n560_0),.q1(n560_1));
  or_bb g183(.a(n177),.b(n182),.q(n183));
  or_bb g777(.a(n764),.b(n776),.q(_w_2940));
  and_bb g280(.a(n277_0),.b(n279),.q(n280));
  spl3L g137_s_1(.a(n137_3),.q0(n137_4),.q1(n137_5),.q2(_w_3192));
  and_bb g276(.a(n192_1),.b(n275_0),.q(n276));
  or_bb g697(.a(n695_0),.b(n696_0),.q(n697));
  bfr _b_2751(.a(_w_3567),.q(_w_3568));
  and_bi g275(.a(n54_1),.b(n274),.q(n275));
  bfr _b_1743(.a(_w_2559),.q(_w_2560));
  and_bi g109(.a(n105_5),.b(n107_1),.q(n109));
  and_bi g526(.a(n525),.b(n524),.q(n526));
  bfr _b_2178(.a(_w_2994),.q(n640));
  and_bb g541(.a(n374_5),.b(n540_0),.q(n541));
  or_bb g494(.a(n492),.b(n493),.q(n494));
  spl4L g395_s_4(.a(n395_15),.q0(n395_16),.q1(n395_17),.q2(n395_18),.q3(n395_19));
  and_bb g267(.a(n254_0),.b(n266),.q(n267));
  spl2 g490_s_1(.a(n490_2),.q0(n490_3),.q1(n490_4));
  or_bb g386(.a(G39_3),.b(G43_0),.q(n386));
  spl2 g409_s_0(.a(n409),.q0(n409_0),.q1(_w_2930));
  bfr _b_1527(.a(_w_2343),.q(_w_2344));
  bfr _b_1955(.a(_w_2771),.q(_w_2772));
  and_bi g97(.a(n95),.b(n96),.q(n97));
  and_bi g262(.a(n260_1),.b(G34_4),.q(n262));
  and_bb g120(.a(n110_0),.b(n119_0),.q(n120));
  bfr _b_2460(.a(_w_3276),.q(_w_3277));
  spl2 g765_s_0(.a(n765),.q0(n765_0),.q1(_w_2928));
  or_bb g419(.a(G4_37),.b(n418),.q(n419));
  or_bb g260(.a(G1_2),.b(G6_1),.q(n260));
  or_bb g101(.a(n100_0),.b(n91_0),.q(n101));
  spl4L G1_s_0(.a(G1),.q0(G1_0),.q1(G1_1),.q2(G1_2),.q3(G1_3));
  and_bb g410(.a(n408_0),.b(n409_1),.q(n410));
  and_bi g654(.a(n392_7),.b(G10_6),.q(n654));
  bfr _b_2574(.a(_w_3390),.q(G3526));
  and_bi g177(.a(G31_7),.b(n145_3),.q(n177));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(_w_2927));
  bfr _b_1830(.a(_w_2646),.q(_w_2647));
  or_bb g119(.a(n117),.b(n118),.q(n119));
  or_bb g243(.a(G9_7),.b(n135_1),.q(n243));
  and_bi g286(.a(G33_7),.b(n151_4),.q(n286));
  spl3L G13_s_6(.a(G13_11),.q0(G13_12),.q1(G13_13),.q2(G13_14));
  bfr _b_2188(.a(_w_3004),.q(_w_3005));
  and_bi g530(.a(n527),.b(n529),.q(_w_2908));
  and_bi g454(.a(G41_7),.b(n398_17),.q(n454));
  spl2 g125_s_0(.a(n125),.q0(n125_0),.q1(n125_1));
  spl2 G42_s_0(.a(G42),.q0(G42_0),.q1(_w_2898));
  bfr _b_1709(.a(_w_2525),.q(_w_2526));
  and_bi g232(.a(n231),.b(n147_11),.q(n232));
  and_bi g551(.a(n549_0),.b(n550),.q(n551));
  spl2 g533_s_1(.a(n533_1),.q0(n533_2),.q1(_w_2896));
  and_bi g631(.a(G21_6),.b(n401_9),.q(n631));
  or_bb g542(.a(n372_2),.b(n541),.q(n542));
  spl3L g240_s_2(.a(n240_3),.q0(n240_4),.q1(n240_5),.q2(n240_6));
  bfr _b_2159(.a(_w_2975),.q(G3531_0));
  and_bi g748(.a(n747),.b(n745),.q(_w_2895));
  or_bb g231(.a(n225),.b(n230),.q(n231));
  or_bb g549(.a(n546_2),.b(n548_0),.q(n549));
  spl2 g282_s_0(.a(n282),.q0(n282_0),.q1(n282_1));
  and_bi g304(.a(n277_1),.b(n303),.q(n304));
  bfr _b_1607(.a(_w_2423),.q(n763));
  and_bi g449(.a(n448),.b(n419_1),.q(n449));
  bfr _b_2175(.a(_w_2991),.q(_w_2992));
  spl2 G39_s_0(.a(_w_3478),.q0(G39_0),.q1(_w_3281));
  and_bi g815(.a(n814_1),.b(n813_1),.q(n815));
  or_bb g648(.a(n385_18),.b(n647),.q(n648));
  bfr _b_1817(.a(_w_2633),.q(_w_2634));
  and_bi g513(.a(n189_2),.b(n496_2),.q(_w_2883));
  bfr _b_2618(.a(_w_3434),.q(_w_3435));
  spl2 g684_s_0(.a(n684),.q0(n684_0),.q1(n684_1));
  and_bi g238(.a(n235_0),.b(n237_0),.q(n238));
  spl2 G11_s_0(.a(_w_3408),.q0(G11_0),.q1(G11_1));
  and_bi g706(.a(n395_18),.b(G14_18),.q(n706));
  or_bb g306(.a(n300),.b(n305),.q(n306));
  bfr _b_2409(.a(_w_3225),.q(G9_5));
  and_bb g438(.a(n436_0),.b(n437_3),.q(n438));
  spl2 G14_s_1(.a(G14_1),.q0(G14_2),.q1(_w_3114));
  bfr _b_1327(.a(_w_2143),.q(_w_2144));
  and_bb g694(.a(n689_1),.b(n692_1),.q(n694));
  and_bi g247(.a(n129_9),.b(n246),.q(n247));
  or_bb g227(.a(G12_3),.b(G4_25),.q(n227));
  and_bi g466(.a(n465),.b(n381_4),.q(_w_2880));
  or_bb g62(.a(n60),.b(n61),.q(n62));
  or_bb g745(.a(n742),.b(n744),.q(n745));
  bfr _b_2450(.a(_w_3266),.q(_w_3267));
  spl4L g401_s_5(.a(n401_15),.q0(n401_19),.q1(n401_20),.q2(n401_21),.q3(n401_22));
  bfr _b_2320(.a(_w_3136),.q(n737_1));
  or_bb g224(.a(n217),.b(n223),.q(n224));
  and_bi g277(.a(n126_3),.b(G3_15),.q(n277));
  or_bb g223(.a(n221),.b(n222),.q(n223));
  and_bi g116(.a(n114),.b(n115),.q(n116));
  bfr _b_2167(.a(_w_2983),.q(n105_3));
  bfr _b_2293(.a(_w_3109),.q(_w_3110));
  spl2 g772_s_0(.a(n772),.q0(n772_0),.q1(n772_1));
  bfr _b_1960(.a(_w_2776),.q(_w_2777));
  spl3L G6_s_0(.a(G6),.q0(G6_0),.q1(G6_1),.q2(_w_2865));
  bfr _b_2031(.a(_w_2847),.q(_w_2848));
  and_bb g345(.a(n240_6),.b(n344_1),.q(_w_2841));
  spl4L G8_s_5(.a(G8_9),.q0(G8_10),.q1(G8_11),.q2(G8_12),.q3(G8_13));
  spl2 g460_s_0(.a(n460),.q0(n460_0),.q1(_w_2839));
  spl2 G1_s_4(.a(G1_11),.q0(G1_12),.q1(_w_2821));
  bfr _b_1636(.a(_w_2452),.q(n123_1));
  and_bb g274(.a(G12_5),.b(G13_6),.q(n274));
  spl4L G3_s_7(.a(G3_17),.q0(G3_20),.q1(G3_21),.q2(G3_22),.q3(G3_23));
  and_bi g225(.a(G32_7),.b(n145_6),.q(n225));
  or_bb g661(.a(G40_3),.b(G44_1),.q(n661));
  bfr _b_2609(.a(_w_3425),.q(_w_3426));
  and_bi g215(.a(n212),.b(n214_0),.q(n215));
  and_bi g384(.a(G26_2),.b(n383_0),.q(n384));
  bfr _b_1360(.a(_w_2176),.q(_w_2177));
  and_bb g214(.a(n201_0),.b(n213),.q(n214));
  and_bb g789(.a(G4_47),.b(n788),.q(n789));
  and_bi g722(.a(n721),.b(n720),.q(n722));
  or_bb g70(.a(n66),.b(n69),.q(n70));
  or_bb g717(.a(n715),.b(n716),.q(n717));
  bfr _b_1543(.a(_w_2359),.q(_w_2360));
  or_bb g212(.a(n201_2),.b(n211),.q(n212));
  spl2 G4_s_12(.a(G4_41),.q0(G4_43),.q1(G4_44));
  spl2 g653_s_0(.a(n653),.q0(n653_0),.q1(_w_2820));
  bfr _b_2694(.a(_w_3510),.q(_w_3511));
  spl2 g631_s_0(.a(n631),.q0(n631_0),.q1(n631_1));
  or_bb g253(.a(n251),.b(n252),.q(n253));
  bfr _b_2490(.a(_w_3306),.q(_w_3307));
  bfr _b_1816(.a(_w_2632),.q(n600));
  or_bb g210(.a(n149_2),.b(n209),.q(_w_2819));
  bfr _b_1567(.a(_w_2383),.q(_w_2384));
  and_bi g595(.a(G4_43),.b(n594),.q(n595));
  and_bi g74(.a(n73_2),.b(G3_26),.q(n74));
  spl2 g162_s_0(.a(n162),.q0(n162_0),.q1(n162_1));
  bfr _b_2087(.a(_w_2903),.q(_w_2904));
  or_bb g646(.a(G8_18),.b(n401_16),.q(n646));
  spl2 g497_s_0(.a(n497),.q0(n497_0),.q1(n497_1));
  or_bb g207(.a(n203),.b(n206),.q(n207));
  and_bi g265(.a(n264),.b(n147_4),.q(n265));
  spl2 g603_s_1(.a(G3531_2),.q0(G3531_3),.q1(_w_2805));
  spl2 g682_s_1(.a(G3533_2),.q0(G3533_3),.q1(_w_3268));
  and_bi g288(.a(G4_15),.b(G34_5),.q(n288));
  bfr _b_2576(.a(_w_3392),.q(n227_1));
  bfr _b_2446(.a(_w_3262),.q(_w_3263));
  spl2 G35_s_3(.a(G35_7),.q0(G35_8),.q1(G35_9));
  bfr _b_2342(.a(_w_3158),.q(_w_3159));
  and_bi g774(.a(n772_1),.b(n683_2),.q(n774));
  or_bb g71(.a(n63),.b(n70),.q(_w_2801));
  and_ii g82(.a(n72),.b(n81),.q(_w_2764));
  bfr _b_2434(.a(_w_3250),.q(_w_3251));
  bfr _b_1309(.a(_w_2125),.q(_w_2126));
  bfr _b_1464(.a(_w_2280),.q(_w_2281));
  or_bi g432(.a(n427),.b(n431),.q(_w_2750));
  bfr _b_1364(.a(_w_2180),.q(_w_2181));
  or_bb g827(.a(n824_0),.b(n826_0),.q(n827));
  bfr _b_1919(.a(_w_2735),.q(_w_2736));
  or_bb g544(.a(n298_1),.b(n543_0),.q(n544));
  and_bb g705(.a(n408_1),.b(n704),.q(n705));
  or_bb g204(.a(G13_2),.b(G4_8),.q(n204));
  bfr _b_2239(.a(_w_3055),.q(_w_3056));
  spl2 g362_s_0(.a(n362),.q0(n362_0),.q1(n362_1));
  bfr _b_1390(.a(_w_2206),.q(n142_2));
  bfr _b_1987(.a(_w_2803),.q(_w_2804));
  spl2 g689_s_0(.a(n689),.q0(n689_0),.q1(n689_1));
  and_bi g226(.a(G30_6),.b(n151_9),.q(_w_2745));
  and_bi g202(.a(G33_6),.b(n145_1),.q(n202));
  and_bi g832(.a(n831),.b(n830),.q(n832));
  and_bb g690(.a(n436_5),.b(n490_1),.q(n690));
  bfr _b_1424(.a(_w_2240),.q(G41_1));
  and_bi g401(.a(n382_3),.b(n394_1),.q(n401));
  and_bi g292(.a(n291),.b(n147_6),.q(_w_2744));
  spl2 G8_s_0(.a(_w_3571),.q0(G8_0),.q1(G8_1));
  or_bb g157(.a(n150),.b(n156),.q(n157));
  spl2 G14_s_2(.a(G14_3),.q0(G14_4),.q1(_w_2743));
  bfr _b_2725(.a(_w_3541),.q(_w_3542));
  spl2 g386_s_0(.a(n386),.q0(n386_0),.q1(_w_2740));
  bfr _b_1823(.a(_w_2639),.q(_w_2640));
  bfr _b_1467(.a(_w_2283),.q(_w_2284));
  and_bi g711(.a(n710),.b(n709),.q(n711));
  and_bi g273(.a(n271),.b(n272),.q(n273));
  and_bb g189(.a(n176_0),.b(n188),.q(n189));
  or_bb g241(.a(G11_4),.b(n54_0),.q(n241));
  bfr _b_1313(.a(_w_2129),.q(n267_1));
  bfr _b_1560(.a(_w_2376),.q(_w_2377));
  bfr _b_1652(.a(_w_2468),.q(_w_2469));
  and_bi g668(.a(G39_10),.b(n407_9),.q(n668));
  and_bb g634(.a(n627_0),.b(n633),.q(n634));
  bfr _b_2090(.a(_w_2906),.q(_w_2907));
  bfr _b_2603(.a(_w_3419),.q(_w_3420));
  or_bb g768(.a(n765_0),.b(n767),.q(n768));
  or_bb g185(.a(n149_1),.b(n184),.q(n185));
  and_bi g186(.a(n143_4),.b(n185_1),.q(_w_2738));
  and_bb g191(.a(n165_0),.b(n190_0),.q(n191));
  bfr _b_2369(.a(_w_3185),.q(_w_3186));
  bfr _b_1792(.a(_w_2608),.q(_w_2609));
  bfr _b_2218(.a(_w_3034),.q(_w_3035));
  and_bb g346(.a(n321_1),.b(n340_3),.q(n346));
  spl2 G3_s_9(.a(G3_25),.q0(G3_26),.q1(G3_27));
  bfr _b_1678(.a(_w_2494),.q(_w_2495));
  and_bb g545(.a(n298_2),.b(n543_1),.q(n545));
  bfr _b_1909(.a(_w_2725),.q(_w_2726));
  or_bb g216(.a(n123_6),.b(n192_0),.q(n216));
  and_bi g257(.a(G4_5),.b(G33_4),.q(n257));
  bfr _b_1344(.a(_w_2160),.q(_w_2161));
  bfr _b_2185(.a(_w_3001),.q(_w_3002));
  or_bb g179(.a(G11_2),.b(G4_13),.q(n179));
  and_bi g178(.a(G29_1),.b(n151_8),.q(n178));
  and_bb g285(.a(G35_8),.b(n283_0),.q(n285));
  or_bb g290(.a(n286),.b(n289),.q(n290));
  bfr _b_2033(.a(_w_2849),.q(_w_2850));
  or_bb g757(.a(n401_20),.b(n455_1),.q(n757));
  spl2 g161_s_0(.a(n161),.q0(n161_0),.q1(n161_1));
  spl2 g275_s_0(.a(n275),.q0(n275_0),.q1(_w_3396));
  and_bi g195(.a(n123_10),.b(G10_10),.q(n195));
  bfr _b_1316(.a(_w_2132),.q(n436_5));
  spl2 g511_s_0(.a(n511),.q0(n511_0),.q1(_w_2995));
  bfr _b_2092(.a(_w_2908),.q(_w_2909));
  spl2 G18_s_0(.a(_w_3427),.q0(G18_0),.q1(_w_2729));
  bfr _b_1442(.a(_w_2258),.q(_w_2259));
  bfr _b_2495(.a(_w_3311),.q(_w_3312));
  or_bb g566(.a(n564),.b(n565),.q(n566));
  bfr _b_1721(.a(_w_2537),.q(_w_2538));
  bfr _b_2517(.a(_w_3333),.q(n369_3));
  bfr _b_1602(.a(_w_2418),.q(n551_1));
  and_bi g108(.a(n107_0),.b(n105_4),.q(n108));
  and_bi g728(.a(n379_8),.b(n727),.q(n728));
  and_bb g407(.a(G3_18),.b(n398_0),.q(n407));
  bfr _b_2177(.a(_w_2993),.q(_w_2994));
  and_bi g213(.a(n162_8),.b(n210_0),.q(n213));
  spl2 G11_s_1(.a(G11_1),.q0(G11_2),.q1(_w_2725));
  or_bb g623(.a(G12_11),.b(n385_5),.q(n623));
  bfr _b_2582(.a(_w_3398),.q(_w_3399));
  bfr _b_1843(.a(_w_2659),.q(_w_2660));
  and_bb g99(.a(n94_1),.b(n97_1),.q(n99));
  or_bb g156(.a(n152),.b(n155),.q(n156));
  or_bb g313(.a(n307),.b(n312),.q(n313));
  bfr _b_1693(.a(_w_2509),.q(_w_2510));
  or_bb g56(.a(G1_10),.b(G3_24),.q(n56));
  and_bb g344(.a(n321_0),.b(n343_2),.q(n344));
  and_bi g337(.a(n336),.b(n147_8),.q(n337));
  bfr _b_2114(.a(_w_2930),.q(_w_2931));
  and_bi g455(.a(G11_10),.b(G39_5),.q(n455));
  bfr _b_1352(.a(_w_2168),.q(_w_2169));
  and_bi g729(.a(n728),.b(n703),.q(_w_2707));
  or_bb g88(.a(n86),.b(n87),.q(n88));
  or_bb g329(.a(n323),.b(n328),.q(n329));
  and_bi g559(.a(n549_1),.b(n558),.q(n559));
  and_bi g701(.a(n697_1),.b(n372_11),.q(n701));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  and_bb g72(.a(n56_0),.b(n71),.q(_w_2704));
  and_bi g100(.a(n98),.b(n99),.q(n100));
  and_bi g107(.a(n52_0),.b(n106),.q(n107));
  bfr _b_1384(.a(_w_2200),.q(_w_2201));
  and_bi g806(.a(n379_9),.b(n805),.q(_w_3171));
  spl2 g546_s_0(.a(n546),.q0(n546_0),.q1(_w_2659));
  and_bb g76(.a(n74_0),.b(n75_0),.q(n76));
  or_bb g363(.a(n320_0),.b(n362_0),.q(n363));
  or_bb g52(.a(G10_9),.b(G7_11),.q(n52));
  bfr _b_1484(.a(_w_2300),.q(_w_2301));
  or_bb g89(.a(n85_0),.b(n88_0),.q(n89));
  bfr _b_1845(.a(_w_2661),.q(n546_1));
  and_bb g134(.a(G3_22),.b(n133),.q(n134));
  and_bi g87(.a(G35_2),.b(G34_2),.q(n87));
  spl2 G5_s_1(.a(G5_2),.q0(G5_3),.q1(_w_2651));
  and_bi g416(.a(n414),.b(n415),.q(n416));
  and_bi g798(.a(n392_9),.b(G7_9),.q(n798));
  or_bb g59(.a(n57),.b(n58),.q(n59));
  and_bb g141(.a(n129_4),.b(n140),.q(n141));
  and_bi g618(.a(n617),.b(n615),.q(n618));
  and_bi g197(.a(n137_4),.b(G11_6),.q(n197));
  bfr _b_2710(.a(_w_3526),.q(_w_3527));
  bfr _b_1315(.a(_w_2131),.q(_w_2132));
  bfr _b_1889(.a(_w_2705),.q(_w_2706));
  and_bi g778(.a(n701_1),.b(n765_1),.q(n778));
  spl2 g146_s_0(.a(n146),.q0(n146_0),.q1(_w_2646));
  and_bb g383(.a(G24_0),.b(G3_0),.q(n383));
  spl2 g176_s_0(.a(n176),.q0(n176_0),.q1(n176_1));
  bfr _b_2350(.a(_w_3166),.q(_w_3167));
  bfr _b_2740(.a(_w_3556),.q(_w_3557));
  and_bi g266(.a(n162_4),.b(n265_4),.q(n266));
  spl2 g344_s_0(.a(n344),.q0(n344_0),.q1(_w_2641));
  or_bb g249(.a(n123_0),.b(n248),.q(n249));
  bfr _b_1498(.a(_w_2314),.q(_w_2315));
  bfr _b_2306(.a(_w_3122),.q(_w_3123));
  spl2 g428_s_0(.a(n428),.q0(n428_0),.q1(n428_1));
  and_bb g340(.a(n329_0),.b(n339),.q(n340));
  bfr _b_1529(.a(_w_2345),.q(_w_2346));
  or_bb g201(.a(n194),.b(n200),.q(n201));
  bfr _b_1759(.a(_w_2575),.q(n437));
  and_bi g457(.a(n456),.b(n454),.q(n457));
  and_bb g79(.a(G34_8),.b(n78),.q(_w_2636));
  or_bb g632(.a(n630_0),.b(n631_0),.q(n632));
  spl3L g407_s_3(.a(n407_11),.q0(n407_12),.q1(n407_13),.q2(n407_14));
  and_bb g164(.a(n142_1),.b(n163),.q(n164));
  bfr _b_1592(.a(_w_2408),.q(_w_2409));
  and_bi g696(.a(n490_6),.b(n507_2),.q(_w_3228));
  and_bi g303(.a(n179_1),.b(n302),.q(_w_2635));
  spl2 g358_s_0(.a(n358),.q0(n358_0),.q1(_w_2633));
  and_bb g356(.a(n161_1),.b(n189_1),.q(n356));
  bfr _b_2496(.a(_w_3312),.q(_w_3313));
  and_bb g237(.a(n224_1),.b(n236),.q(n237));
  spl4L g395_s_0(.a(n395),.q0(n395_0),.q1(n395_1),.q2(n395_2),.q3(n395_3));
  and_bi g93(.a(G31_2),.b(G30_2),.q(n93));
  or_bb g143(.a(G25_0),.b(G26_0),.q(n143));
  and_bi g600(.a(n599),.b(n381_5),.q(_w_2630));
  or_bb g554(.a(n552),.b(n553_0),.q(n554));
  and_bb g84(.a(G36_2),.b(G37_2),.q(n84));
  or_bb g674(.a(n659),.b(n673),.q(n674));
  and_bi g92(.a(G30_1),.b(G31_1),.q(n92));
  and_bb g585(.a(n580),.b(n584),.q(n585));
  and_bi g172(.a(n171_0),.b(G4_33),.q(n172));
  and_bb g299(.a(n270_0),.b(n298_0),.q(n299));
  spl2 g630_s_0(.a(n630),.q0(n630_0),.q1(n630_1));
  spl2 g94_s_0(.a(n94),.q0(n94_0),.q1(n94_1));
  or_bb g271(.a(G12_9),.b(n123_8),.q(n271));
  spl2 g143_s_0(.a(n143),.q0(n143_0),.q1(_w_2624));
  and_bi g379(.a(n372_0),.b(G6_2),.q(n379));
  spl2 G3_s_6(.a(G3_16),.q0(G3_18),.q1(G3_19));
  and_bi g581(.a(n392_4),.b(G9_11),.q(n581));
  spl3L G30_s_1(.a(G30_3),.q0(_w_2622),.q1(G30_5),.q2(_w_2623));
  and_bi g298(.a(n297),.b(n295_0),.q(n298));
  bfr _b_1857(.a(_w_2673),.q(_w_2674));
  and_bb g486(.a(n481_0),.b(n484_0),.q(n486));
  bfr _b_1486(.a(_w_2302),.q(_w_2303));
  or_bb g442(.a(n440),.b(n441),.q(n442));
  and_bb g308(.a(G35_4),.b(G4_16),.q(n308));
  bfr _b_1682(.a(_w_2498),.q(_w_2499));
  spl4L G34_s_0(.a(_w_3472),.q0(G34_0),.q1(G34_1),.q2(G34_2),.q3(G34_3));
  bfr _b_1373(.a(_w_2189),.q(G19_3));
  or_bb g233(.a(n149_3),.b(n232),.q(n233));
  and_bi g564(.a(n559_0),.b(n563_2),.q(n564));
  bfr _b_1522(.a(_w_2338),.q(_w_2339));
  bfr _b_1644(.a(_w_2460),.q(n361_9));
  and_bi g263(.a(n261),.b(n262),.q(_w_3188));
  and_bi g373(.a(n75_1),.b(n372_12),.q(n373));
  bfr _b_1882(.a(_w_2698),.q(_w_2699));
  spl2 G50_s_0(.a(_w_3525),.q0(G50_0),.q1(_w_2621));
  and_bb g175(.a(n129_6),.b(n174),.q(n175));
  and_bi g198(.a(n196),.b(n197),.q(n198));
  or_bb g688(.a(n683_0),.b(n687),.q(_w_3086));
  and_bb g562(.a(n270_2),.b(n560_1),.q(n562));
  or_bb g81(.a(n76),.b(n80),.q(n81));
  and_bb g169(.a(G3_21),.b(n105_0),.q(n169));
  spl2 g317_s_1(.a(n317_1),.q0(n317_2),.q1(_w_2619));
  or_bb g114(.a(G12_16),.b(G14_14),.q(n114));
  and_bi g467(.a(n379_5),.b(n466),.q(_w_2618));
  spl3L G39_s_1(.a(G39_1),.q0(G39_2),.q1(G39_3),.q2(_w_3133));
  spl3L g56_s_0(.a(n56),.q0(n56_0),.q1(n56_1),.q2(_w_2615));
  spl2 g216_s_0(.a(n216),.q0(n216_0),.q1(n216_1));
  and_bb g317(.a(n306_0),.b(n316),.q(n317));
  or_bb g351(.a(n346),.b(n350),.q(n351));
  and_bb g146(.a(G4_0),.b(G5_1),.q(n146));
  and_bb g149(.a(n145_5),.b(n148_0),.q(n149));
  or_bb g235(.a(n224_0),.b(n234),.q(n235));
  bfr _b_1340(.a(_w_2156),.q(_w_2157));
  bfr _b_1980(.a(_w_2796),.q(_w_2797));
  spl2 G18_s_1(.a(G18_1),.q0(G18_2),.q1(G18_3));
  bfr _b_2233(.a(_w_3049),.q(_w_3050));
  and_bi g136(.a(G21_0),.b(n135_0),.q(n136));
  and_bi g816(.a(n815),.b(n812_0),.q(n816));
  or_bb g287(.a(G39_0),.b(G4_14),.q(n287));
  bfr _b_2118(.a(_w_2934),.q(_w_2935));
  or_bb g269(.a(n254_1),.b(n268),.q(n269));
  spl3L g135_s_0(.a(n135),.q0(n135_0),.q1(n135_1),.q2(n135_2));
  and_bi g754(.a(n395_11),.b(G13_16),.q(n754));
  and_bb g90(.a(n85_1),.b(n88_1),.q(n90));
  or_bb g741(.a(n739),.b(n740),.q(n741));
  and_bb g393(.a(G40_2),.b(n392_0),.q(n393));
  bfr _b_1432(.a(_w_2248),.q(_w_2249));
  and_bb g396(.a(G44_0),.b(n395_0),.q(n396));
  bfr _b_2491(.a(_w_3307),.q(_w_3308));
  or_bb g208(.a(n202),.b(n207),.q(n208));
  spl4L G13_s_8(.a(G13_17),.q0(G13_18),.q1(G13_19),.q2(G13_20),.q3(_w_2610));
  bfr _b_1423(.a(_w_2239),.q(n293_3));
  and_bi g150(.a(G30_4),.b(n145_0),.q(n150));
  or_bb g63(.a(n59),.b(n62),.q(n63));
  bfr _b_1744(.a(_w_2560),.q(_w_2561));
  spl2 G3_s_0(.a(G3),.q0(G3_0),.q1(G3_1));
  spl2 g51_s_1(.a(n51_1),.q0(n51_2),.q1(_w_2607));
  or_bb g761(.a(n750),.b(n760),.q(n761));
  or_bb g279(.a(n153_1),.b(n278),.q(n279));
  and_bb g536(.a(n320_4),.b(n534_1),.q(_w_3391));
  and_bi g284(.a(n148_1),.b(n283_3),.q(n284));
  and_bi g91(.a(n89),.b(n90),.q(n91));
  and_bb g239(.a(n215_0),.b(n238_0),.q(n239));
  or_bb g521(.a(G1_12),.b(G2_5),.q(n521));
  and_bb g671(.a(G4_45),.b(n670),.q(n671));
  or_bb g220(.a(n218),.b(n219),.q(n220));
  or_bb g836(.a(G50_0),.b(n834_0),.q(n836));
  bfr _b_1622(.a(_w_2438),.q(n192_3));
  bfr _b_2124(.a(_w_2940),.q(G3535_0));
  and_bi g222(.a(G9_13),.b(n130_4),.q(n222));
  or_bb g408(.a(G11_17),.b(n407_4),.q(n408));
  spl2 g810_s_1(.a(G3536_2),.q0(G3536_3),.q1(_w_2599));
  bfr _b_2683(.a(_w_3499),.q(_w_3500));
  and_bi g206(.a(n204),.b(n205),.q(n206));
  spl2 g129_s_1(.a(n129_3),.q0(_w_2598),.q1(n129_5));
  and_bi g739(.a(G16_0),.b(n398_10),.q(n739));
  bfr _b_1301(.a(_w_2117),.q(_w_2118));
  bfr _b_2301(.a(_w_3117),.q(_w_3118));
  and_bi g64(.a(G34_0),.b(G11_0),.q(n64));
  or_bb g264(.a(n259),.b(n263),.q(n264));
  spl2 g210_s_0(.a(n210),.q0(n210_0),.q1(_w_2597));
  bfr _b_1416(.a(_w_2232),.q(_w_2233));
  bfr _b_2456(.a(_w_3272),.q(_w_3273));
  bfr _b_1643(.a(_w_2459),.q(n203));
  spl2 g480_s_0(.a(n480),.q0(n480_0),.q1(n480_1));
  bfr _b_1797(.a(_w_2613),.q(_w_2614));
  or_bb g66(.a(n64),.b(n65),.q(n66));
  or_bb g124(.a(G7_7),.b(n123_4),.q(n124));
  or_bb g77(.a(G2_3),.b(n56_1),.q(n77));
  spl2 G10_s_1(.a(G10_2),.q0(G10_3),.q1(G10_4));
  spl3L g514_s_0(.a(n514),.q0(n514_0),.q1(n514_1),.q2(n514_2));
  and_bi g468(.a(n467),.b(n438),.q(_w_2587));
  spl4L G11_s_6(.a(G11_14),.q0(G11_15),.q1(G11_16),.q2(G11_17),.q3(G11_18));
  bfr _b_1779(.a(_w_2595),.q(_w_2596));
  spl2 g641_s_1(.a(G3532_2),.q0(G3532_3),.q1(_w_2576));
  spl2 g51_s_0(.a(n51),.q0(n51_0),.q1(n51_1));
  and_bi g234(.a(n143_6),.b(n233_0),.q(n234));
  bfr _b_2344(.a(_w_3160),.q(n164_1));
  and_bi g540(.a(n538),.b(n539),.q(n540));
  or_bb g297(.a(n282_2),.b(n296),.q(n297));
  or_bb g447(.a(n385_11),.b(n446),.q(n447));
  or_bb g506(.a(n240_2),.b(n374_1),.q(n506));
  bfr _b_1474(.a(_w_2290),.q(_w_2291));
  bfr _b_2642(.a(_w_3458),.q(_w_3459));
  spl2 g455_s_0(.a(n455),.q0(n455_0),.q1(n455_1));
  or_bb g256(.a(G14_2),.b(G4_6),.q(n256));
  bfr _b_1318(.a(_w_2134),.q(_w_2135));
  or_bb g465(.a(n451),.b(n464),.q(n465));
  and_bb g574(.a(G21_2),.b(n395_1),.q(n574));
  bfr _b_1582(.a(_w_2398),.q(_w_2399));
  and_bi g445(.a(G18_3),.b(n401_13),.q(n445));
  bfr _b_1877(.a(_w_2693),.q(_w_2694));
  bfr _b_2728(.a(_w_3544),.q(_w_3545));
  spl3L G12_s_1(.a(G12_1),.q0(G12_2),.q1(G12_3),.q2(G12_4));
  spl2 g432_s_0(.a(G3528_0),.q0(G3528_1),.q1(G3528_2));
  or_bb g358(.a(n355),.b(n357),.q(_w_2732));
  and_bi g762(.a(n761),.b(n381_9),.q(_w_2569));
  and_bb g439(.a(G20_6),.b(n395_19),.q(_w_2568));
  bfr _b_1999(.a(_w_2815),.q(G3531));
  and_bb g166(.a(G8_10),.b(n130_1),.q(n166));
  or_bb g409(.a(G13_13),.b(n385_3),.q(n409));
  and_bi g672(.a(n671),.b(n668),.q(n672));
  bfr _b_2096(.a(_w_2912),.q(_w_2913));
  spl2 g372_s_3(.a(n372_5),.q0(n372_6),.q1(_w_2562));
  and_bi g122(.a(n121),.b(n120),.q(_w_2528));
  and_bi g86(.a(G34_1),.b(G35_1),.q(n86));
  bfr _b_1457(.a(_w_2273),.q(_w_2274));
  and_bi g738(.a(n737_1),.b(n385_21),.q(n738));
  bfr _b_1587(.a(_w_2403),.q(_w_2404));
  bfr _b_2398(.a(_w_3214),.q(n349));
  bfr _b_1773(.a(_w_2589),.q(_w_2590));
  and_bb g325(.a(G39_2),.b(G4_32),.q(n325));
  or_bb g610(.a(n608),.b(n609),.q(n610));
  and_bi g389(.a(G4_36),.b(n388),.q(n389));
  bfr _b_2137(.a(_w_2953),.q(_w_2954));
  or_bb g514(.a(n512_0),.b(n513),.q(n514));
  bfr _b_1623(.a(_w_2439),.q(_w_2440));
  spl4L g392_s_3(.a(n392_10),.q0(n392_11),.q1(n392_12),.q2(n392_13),.q3(_w_2527));
  spl4L G35_s_0(.a(_w_3473),.q0(G35_0),.q1(G35_1),.q2(G35_2),.q3(G35_3));
  and_bb g791(.a(n786),.b(n790),.q(n791));
  or_bb g167(.a(G8_11),.b(n123_5),.q(n167));
  and_bb g580(.a(n577),.b(n579),.q(_w_2525));
  spl2 g143_s_3(.a(n143_9),.q0(n143_10),.q1(n143_11));
  or_bb g812(.a(G3529_1),.b(G3536_1),.q(n812));
  and_bi g381(.a(n73_4),.b(n380),.q(_w_2523));
  bfr _b_1662(.a(_w_2478),.q(_w_2479));
  and_bi g606(.a(n533_0),.b(n540_1),.q(n606));
  bfr _b_2081(.a(_w_2897),.q(n533_3));
  and_bi g375(.a(n374_10),.b(G1_13),.q(_w_2512));
  bfr _b_1362(.a(_w_2178),.q(_w_2179));
  and_bb g126(.a(G1_1),.b(G2_1),.q(n126));
  and_bi g193(.a(n130_3),.b(n192_3),.q(n193));
  and_bi g296(.a(n143_7),.b(n293_3),.q(n296));
  bfr _b_2653(.a(G31),.q(_w_3469));
  and_bi g168(.a(n167),.b(n166),.q(n168));
  and_bi g388(.a(G41_4),.b(G3_19),.q(n388));
  bfr _b_1888(.a(_w_2704),.q(_w_2705));
  bfr _b_2305(.a(_w_3121),.q(_w_3122));
  or_bb g187(.a(n176_2),.b(n186),.q(n187));
  and_bb g793(.a(G19_4),.b(n395_13),.q(n793));
  and_bi g575(.a(G20_0),.b(n398_2),.q(n575));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(_w_2735));
  or_bb g129(.a(n126_2),.b(n128),.q(n129));
  bfr _b_2154(.a(_w_2970),.q(_w_2971));
  spl2 g374_s_4(.a(n374_8),.q0(_w_2509),.q1(n374_10));
  and_bi g300(.a(n216_1),.b(G13_20),.q(n300));
  bfr _b_1415(.a(_w_2231),.q(_w_2232));
  and_bi g426(.a(n379_4),.b(n425),.q(_w_2611));
  and_bi g589(.a(n588),.b(n586),.q(n589));
  bfr _b_2209(.a(_w_3025),.q(_w_3026));
  spl4L G36_s_0(.a(_w_3474),.q0(G36_0),.q1(G36_1),.q2(G36_2),.q3(G36_3));
  bfr _b_1553(.a(_w_2369),.q(n379_10));
  bfr _b_1841(.a(_w_2657),.q(_w_2658));
  spl2 g123_s_1(.a(n123_1),.q0(n123_2),.q1(n123_3));
  bfr _b_1917(.a(_w_2733),.q(_w_2734));
  or_bb g130(.a(n125_0),.b(n129_0),.q(n130));
  or_bb g254(.a(n247),.b(n253),.q(n254));
  or_bb g628(.a(G8_12),.b(n385_6),.q(n628));
  bfr _b_2527(.a(_w_3343),.q(n676));
  and_bi g547(.a(n317_3),.b(n361_15),.q(_w_2508));
  or_bb g135(.a(G3_8),.b(G4_23),.q(n135));
  bfr _b_1762(.a(_w_2578),.q(_w_2579));
  and_bi g441(.a(G19_5),.b(n398_19),.q(n441));
  or_bb g174(.a(n169),.b(n173),.q(n174));
  spl2 g116_s_0(.a(n116),.q0(n116_0),.q1(n116_1));
  spl4L G10_s_3(.a(G10_8),.q0(G10_9),.q1(G10_10),.q2(G10_11),.q3(G10_12));
  spl3L G40_s_2(.a(G40_4),.q0(G40_5),.q1(G40_6),.q2(G40_7));
  bfr _b_1879(.a(_w_2695),.q(_w_2696));
  and_bi g750(.a(n749),.b(n738),.q(_w_2507));
  or_bb g133(.a(G7_2),.b(n51_2),.q(n133));
  bfr _b_1435(.a(_w_2251),.q(_w_2252));
  spl3L g683_s_0(.a(n683),.q0(n683_0),.q1(n683_1),.q2(n683_2));
  or_bb g200(.a(n195),.b(n199),.q(n200));
  and_bb g154(.a(G29_0),.b(G4_7),.q(_w_2505));
  bfr _b_1932(.a(_w_2748),.q(G40_1));
  and_bi g137(.a(G4_27),.b(G3_9),.q(n137));
  bfr _b_2406(.a(_w_3222),.q(G17_1));
  spl4L g151_s_0(.a(n151),.q0(n151_0),.q1(n151_1),.q2(_w_2504),.q3(n151_3));
  bfr _b_2420(.a(_w_3236),.q(_w_3237));
  or_bb g250(.a(n129_2),.b(n249),.q(n250));
  bfr _b_1414(.a(_w_2230),.q(_w_2231));
  or_bb g651(.a(G9_19),.b(n407_14),.q(n651));
  bfr _b_1564(.a(_w_2380),.q(_w_2381));
  and_bi g565(.a(n563_3),.b(n559_1),.q(n565));
  and_bb g751(.a(G5_5),.b(n627_1),.q(n751));
  bfr _b_1730(.a(_w_2546),.q(_w_2547));
  or_bb g140(.a(n134),.b(n139),.q(n140));
  or_bb g144(.a(G5_0),.b(G6_0),.q(n144));
  and_bb g591(.a(G41_8),.b(n395_16),.q(n591));
  bfr _b_2054(.a(_w_2870),.q(_w_2871));
  and_bi g318(.a(n143_11),.b(n315_3),.q(n318));
  spl3L G9_s_3(.a(G9_5),.q0(G9_6),.q1(G9_7),.q2(_w_3394));
  or_bb g151(.a(G4_1),.b(_w_3524),.q(n151));
  spl2 g269_s_0(.a(n269),.q0(n269_0),.q1(n269_1));
  and_bi g509(.a(n214_2),.b(n361_10),.q(n509));
  and_bi g145(.a(n144),.b(G1_5),.q(_w_2502));
  and_bi g65(.a(G35_0),.b(G12_0),.q(n65));
  bfr _b_2464(.a(_w_3280),.q(G41_6));
  and_bi g163(.a(n162_2),.b(n159_1),.q(n163));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(n88_1));
  bfr _b_1445(.a(_w_2261),.q(_w_2262));
  and_bi g289(.a(n287),.b(n288),.q(n289));
  or_ii g55(.a(G11_18),.b(n54_2),.q(_w_2461));
  bfr _b_2098(.a(_w_2914),.q(_w_2915));
  and_bi g834(.a(n811_1),.b(n833),.q(n834));
  and_bi g638(.a(n379_7),.b(n637),.q(_w_2739));
  and_bi g517(.a(n516),.b(n515),.q(n517));
  and_bi g520(.a(n519),.b(n518),.q(n520));
  and_bi g584(.a(n583),.b(G4_51),.q(n584));
  and_bi g117(.a(n113_0),.b(n116_0),.q(n117));
  and_bb g392(.a(G3_12),.b(n391),.q(n392));
  and_bi g148(.a(G38_1),.b(n147_0),.q(n148));
  bfr _b_1653(.a(_w_2469),.q(_w_2470));
  spl2 g361_s_2(.a(n361_7),.q0(n361_8),.q1(_w_2460));
  spl2 g265_s_1(.a(n265_1),.q0(n265_2),.q1(n265_3));
  and_bb g463(.a(n459),.b(n462),.q(n463));
  or_bb g434(.a(n215_1),.b(n433_0),.q(n434));
  or_bb g139(.a(n136),.b(n138),.q(n139));
  or_bb g155(.a(n153_0),.b(n154),.q(n155));
  and_bb g423(.a(n410),.b(n422),.q(n423));
  spl2 g126_s_0(.a(n126),.q0(n126_0),.q1(n126_1));
  and_bi g125(.a(G3_6),.b(G1_7),.q(n125));
  bfr _b_1769(.a(_w_2585),.q(_w_2586));
  spl4L g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1),.q2(n137_2),.q3(n137_3));
  and_bi g105(.a(n51_0),.b(n104),.q(n105));
  and_bi g203(.a(G31_4),.b(n151_1),.q(_w_2459));
  or_bb g478(.a(n361_8),.b(n477),.q(_w_2453));
  spl3L g392_s_1(.a(n392_2),.q0(n392_4),.q1(n392_5),.q2(n392_6));
  and_bb g473(.a(n315_0),.b(n338_1),.q(n473));
  spl2 g123_s_0(.a(n123),.q0(n123_0),.q1(_w_2452));
  and_bi g190(.a(n187),.b(n189_0),.q(n190));
  or_bb g431(.a(n428_0),.b(n430),.q(n431));
  bfr _b_2283(.a(_w_3099),.q(_w_3100));
  bfr _b_1339(.a(_w_2155),.q(_w_2156));
  or_bi g841(.a(n839),.b(n840),.q(G3539));
  bfr _b_1557(.a(_w_2373),.q(n406));
  bfr _b_1801(.a(_w_2617),.q(n56_2));
  and_bi g158(.a(n157),.b(n147_2),.q(_w_2451));
  or_bb g685(.a(n500_4),.b(n511_1),.q(n685));
  spl4L g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1),.q2(n149_2),.q3(_w_2450));
  spl2 g379_s_3(.a(n379_10),.q0(n379_11),.q1(_w_2442));
  and_bi g568(.a(n566_1),.b(n553_3),.q(n568));
  and_bb g219(.a(G10_3),.b(n137_5),.q(n219));
  bfr _b_1395(.a(_w_2211),.q(_w_2212));
  spl4L g392_s_2(.a(n392_3),.q0(n392_7),.q1(n392_8),.q2(n392_9),.q3(n392_10));
  and_bb g307(.a(G36_6),.b(n283_1),.q(n307));
  or_bb g161(.a(n142_0),.b(n160),.q(n161));
  and_bb g321(.a(n299_0),.b(n320_3),.q(n321));
  or_bb g162(.a(G23_0),.b(G24_4),.q(n162));
  and_bi g630(.a(n392_6),.b(G11_11),.q(n630));
  bfr _b_1584(.a(_w_2400),.q(_w_2401));
  and_bi g548(.a(n535_1),.b(n547),.q(n548));
  and_bi g563(.a(n561),.b(n562),.q(_w_2441));
  and_bb g417(.a(n413),.b(n416),.q(n417));
  bfr _b_2523(.a(_w_3339),.q(_w_3340));
  and_bb g435(.a(n215_2),.b(n433_1),.q(n435));
  bfr _b_2077(.a(_w_2893),.q(_w_2894));
  and_bi g170(.a(n137_1),.b(G9_6),.q(n170));
  spl2 g145_s_1(.a(n145_2),.q0(n145_3),.q1(n145_4));
  bfr _b_1507(.a(_w_2323),.q(n481));
  bfr _b_1782(.a(_w_2598),.q(n129_4));
  bfr _b_2032(.a(_w_2848),.q(_w_2849));
  or_bb g98(.a(n94_0),.b(n97_0),.q(n98));
  bfr _b_1828(.a(_w_2644),.q(_w_2645));
  spl3L G21_s_2(.a(G21_4),.q0(G21_5),.q1(G21_6),.q2(G21_7));
  bfr _b_1953(.a(_w_2769),.q(_w_2770));
  bfr _b_1683(.a(_w_2499),.q(_w_2500));
  spl2 g135_s_1(.a(n135_2),.q0(n135_3),.q1(n135_4));
  and_bi g524(.a(G7_20),.b(G9_18),.q(n524));
  spl2 g317_s_0(.a(n317),.q0(n317_0),.q1(_w_2439));
  and_bb g452(.a(G40_8),.b(n395_14),.q(n452));
  bfr _b_2255(.a(_w_3071),.q(_w_3072));
  spl3L G10_s_4(.a(G10_12),.q0(G10_13),.q1(G10_14),.q2(G10_15));
  bfr _b_2153(.a(_w_2969),.q(_w_2970));
  spl4L g382_s_0(.a(n382),.q0(n382_0),.q1(n382_1),.q2(n382_2),.q3(n382_3));
  spl4L g377_s_0(.a(n377),.q0(_w_2437),.q1(n377_1),.q2(n377_2),.q3(n377_3));
  and_bi g171(.a(G22_0),.b(G3_10),.q(n171));
  or_bb g110(.a(n108),.b(n109),.q(n110));
  and_bi g309(.a(G40_0),.b(G4_17),.q(n309));
  or_bb g196(.a(G8_8),.b(n135_3),.q(n196));
  bfr _b_2734(.a(_w_3550),.q(_w_3551));
  bfr _b_2655(.a(G33),.q(_w_3471));
  or_bb g310(.a(n308),.b(n309),.q(n310));
  spl2 g517_s_0(.a(n517),.q0(n517_0),.q1(n517_1));
  bfr _b_2608(.a(_w_3424),.q(_w_3425));
  or_bb g485(.a(n481_1),.b(n484_1),.q(_w_2436));
  and_bi g147(.a(n126_0),.b(n146_0),.q(n147));
  spl2 g500_s_0(.a(n500),.q0(n500_0),.q1(_w_2433));
  and_bb g539(.a(n428_3),.b(n537_1),.q(n539));
  bfr _b_1733(.a(_w_2549),.q(_w_2550));
  spl4L G14_s_6(.a(G14_15),.q0(G14_16),.q1(G14_17),.q2(G14_18),.q3(_w_3231));
  bfr _b_2289(.a(_w_3105),.q(n764));
  or_bb g51(.a(G8_2),.b(G9_2),.q(n51));
  and_bb g104(.a(G8_4),.b(G9_4),.q(n104));
  and_bi g380(.a(G3_27),.b(G23_1),.q(n380));
  bfr _b_1310(.a(_w_2126),.q(n494_4));
  bfr _b_2333(.a(_w_3149),.q(n329_3));
  and_bb g362(.a(n306_3),.b(n361_4),.q(n362));
  and_bb g278(.a(G13_8),.b(G4_34),.q(n278));
  and_bb g127(.a(G1_4),.b(G3_2),.q(n127));
  and_bi g311(.a(G34_7),.b(n151_5),.q(n311));
  or_bb g312(.a(n310),.b(n311),.q(n312));
  and_bi g675(.a(n674),.b(n381_7),.q(_w_2431));
  and_bb g512(.a(n500_2),.b(n511_0),.q(n512));
  and_bi g504(.a(n503),.b(n502),.q(n504));
  and_bb g96(.a(G32_2),.b(G33_2),.q(n96));
  or_bb g395(.a(n382_1),.b(n394_0),.q(n395));
  and_bi g320(.a(n319),.b(n317_0),.q(n320));
  and_bi g361(.a(n360_0),.b(n77_1),.q(n361));
  bfr _b_1815(.a(_w_2631),.q(_w_2632));
  spl3L g381_s_1(.a(n381_1),.q0(n381_3),.q1(n381_4),.q2(n381_5));
  and_bi g567(.a(n553_2),.b(n566_0),.q(n567));
  bfr _b_1532(.a(_w_2348),.q(_w_2349));
  or_bb g498(.a(n190_1),.b(n497_0),.q(n498));
  bfr _b_2256(.a(_w_3072),.q(_w_3073));
  or_bb g391(.a(G24_2),.b(n143_0),.q(n391));
  and_bi g637(.a(n636),.b(n381_6),.q(_w_2984));
  spl4L G14_s_5(.a(G14_11),.q0(G14_12),.q1(G14_13),.q2(_w_2430),.q3(G14_15));
  or_bb g731(.a(n700),.b(n730),.q(G3534_0));
  bfr _b_1418(.a(_w_2234),.q(_w_2235));
  and_bi g323(.a(G14_12),.b(n322),.q(n323));
  bfr _b_2514(.a(_w_3330),.q(_w_3331));
  bfr _b_1392(.a(_w_2208),.q(G22_9));
  bfr _b_1860(.a(_w_2676),.q(_w_2677));
  or_bb g402(.a(G42_0),.b(_w_3494),.q(_w_2425));
  spl2 g535_s_0(.a(n535),.q0(n535_0),.q1(n535_1));
  spl4L g401_s_2(.a(n401_3),.q0(n401_8),.q1(n401_9),.q2(_w_2424),.q3(n401_11));
  bfr _b_1963(.a(_w_2779),.q(_w_2780));
  bfr _b_2564(.a(_w_3380),.q(_w_3381));
  or_bb g349(.a(n267_1),.b(n348),.q(_w_3212));
  bfr _b_1921(.a(_w_2737),.q(n153_1));
  bfr _b_2219(.a(_w_3035),.q(_w_3036));
  spl3L g361_s_3(.a(n361_9),.q0(n361_10),.q1(n361_11),.q2(n361_12));
  bfr _b_1544(.a(_w_2360),.q(n477));
  and_bi g218(.a(G7_5),.b(n135_4),.q(n218));
  bfr _b_1633(.a(_w_2449),.q(n379_12));
  and_bi g709(.a(G39_11),.b(n398_20),.q(n709));
  spl3L G7_s_1(.a(G7_1),.q0(G7_2),.q1(G7_3),.q2(G7_4));
  bfr _b_1328(.a(_w_2144),.q(n237_3));
  bfr _b_2644(.a(_w_3460),.q(_w_3461));
  bfr _b_2117(.a(_w_2933),.q(_w_2934));
  or_bb g328(.a(n324),.b(n327),.q(n328));
  or_bb g293(.a(n284_0),.b(n292),.q(n293));
  spl4L G4_s_5(.a(G4_11),.q0(G4_19),.q1(G4_20),.q2(G4_21),.q3(G4_22));
  spl2 g164_s_0(.a(n164),.q0(n164_0),.q1(_w_3160));
  spl2 G11_s_2(.a(G11_3),.q0(G11_4),.q1(G11_5));
  spl2 G40_s_0(.a(_w_3480),.q0(G40_0),.q1(_w_2746));
  bfr _b_1750(.a(_w_2566),.q(_w_2567));
  and_bb g330(.a(G37_3),.b(n283_2),.q(n330));
  or_bb g54(.a(G12_2),.b(G13_4),.q(n54));
  spl4L g381_s_2(.a(n381_2),.q0(n381_6),.q1(n381_7),.q2(n381_8),.q3(n381_9));
  and_bi g334(.a(G35_6),.b(n151_6),.q(n334));
  bfr _b_1935(.a(_w_2751),.q(_w_2752));
  and_bb g413(.a(n411_0),.b(n412),.q(n413));
  or_bb g336(.a(n330),.b(n335),.q(n336));
  and_bi g583(.a(n582),.b(n581_1),.q(n583));
  and_bb g353(.a(n214_1),.b(n235_1),.q(n353));
  or_bb g338(.a(n284_2),.b(n337_0),.q(n338));
  and_bi g590(.a(G42_5),.b(n398_16),.q(n590));
  or_bb g576(.a(n574),.b(n575),.q(n576));
  or_bb g342(.a(n329_2),.b(n341),.q(n342));
  and_bi g343(.a(n342),.b(n340_0),.q(n343));
  and_bi g246(.a(n245),.b(n242),.q(n246));
  and_bi g507(.a(n506),.b(n358_1),.q(n507));
  spl2 g237_s_0(.a(n237),.q0(n237_0),.q1(n237_1));
  spl2 G5_s_2(.a(G5_4),.q0(G5_5),.q1(G5_6));
  and_bi g244(.a(n137_2),.b(G12_7),.q(n244));
  bfr _b_2046(.a(_w_2862),.q(_w_2863));
  or_bb g459(.a(G13_21),.b(n407_13),.q(n459));
  or_bb g582(.a(G8_17),.b(n407_5),.q(n582));
  or_bb g350(.a(n347),.b(n349),.q(_w_2422));
  bfr _b_2641(.a(_w_3457),.q(_w_3458));
  or_bb g809(.a(n807),.b(n808),.q(_w_2419));
  spl3L G8_s_7(.a(G8_15),.q0(G8_16),.q1(G8_17),.q2(G8_18));
  bfr _b_1548(.a(_w_2364),.q(n152));
  and_bb g502(.a(n240_4),.b(n501_0),.q(n502));
  spl3L G10_s_0(.a(_w_3407),.q0(G10_0),.q1(G10_1),.q2(_w_3344));
  and_bi g650(.a(n649),.b(n645),.q(n650));
  spl2 g551_s_0(.a(n551),.q0(n551_0),.q1(_w_2418));
  or_bb g283(.a(G5_3),.b(n260_2),.q(n283));
  or_bb g354(.a(n237_2),.b(n353),.q(_w_2417));
  or_bb g121(.a(n110_1),.b(n119_1),.q(n121));
  or_bb g357(.a(n164_1),.b(n356),.q(_w_2414));
  or_bb g682(.a(n643),.b(n681),.q(_w_3051));
  or_bb g359(.a(n352),.b(n358_0),.q(_w_2385));
  bfr _b_2668(.a(_w_3484),.q(_w_3485));
  and_bb g272(.a(G12_10),.b(n250_1),.q(n272));
  and_bb g364(.a(n320_1),.b(n362_1),.q(n364));
  bfr _b_1880(.a(_w_2696),.q(_w_2697));
  and_bb g462(.a(G4_49),.b(n461),.q(n462));
  spl2 g549_s_0(.a(n549),.q0(n549_0),.q1(n549_1));
  and_bi g322(.a(n250_3),.b(n192_2),.q(n322));
  or_bb g784(.a(n385_15),.b(n783),.q(n784));
  bfr _b_2023(.a(_w_2839),.q(n460_1));
  or_bb g367(.a(n343_0),.b(n366_0),.q(n367));
  and_bb g368(.a(n343_1),.b(n366_1),.q(n368));
  and_bb g370(.a(G47_3),.b(n369_3),.q(n370));
  bfr _b_1754(.a(_w_2570),.q(n762));
  and_bi g727(.a(n726),.b(n381_8),.q(_w_2382));
  and_bb g242(.a(G3_20),.b(n241),.q(n242));
  bfr _b_2556(.a(_w_3372),.q(_w_3373));
  and_bi g61(.a(G37_0),.b(G14_0),.q(n61));
  and_bb g598(.a(n589),.b(n597),.q(n598));
  bfr _b_1613(.a(_w_2429),.q(n402));
  and_bi g372(.a(G5_6),.b(n77_3),.q(_w_2380));
  and_bi g374(.a(n351_1),.b(n361_19),.q(n374));
  bfr _b_2354(.a(_w_3170),.q(G12_8));
  and_bi g679(.a(n678),.b(n533_2),.q(n679));
  bfr _b_2232(.a(_w_3048),.q(_w_3049));
  bfr _b_1855(.a(_w_2671),.q(_w_2672));
  bfr _b_2675(.a(_w_3491),.q(_w_3492));
  and_bi g492(.a(n238_1),.b(n491_0),.q(n492));
  and_bi g377(.a(n137_6),.b(G2_7),.q(_w_2374));
  bfr _b_1596(.a(_w_2412),.q(_w_2413));
  and_bi g406(.a(n390),.b(n405),.q(_w_2371));
  bfr _b_2294(.a(_w_3110),.q(_w_3111));
  bfr _b_2435(.a(_w_3251),.q(_w_3252));
  bfr _b_2363(.a(_w_3179),.q(_w_3180));
  and_bi g387(.a(n386_0),.b(n385_0),.q(n387));
  spl2 g371_s_0(.a(G3526_0),.q0(G3526_1),.q1(G3526_2));
  and_bb g366(.a(n329_3),.b(n361_0),.q(n366));
  bfr _b_1856(.a(_w_2672),.q(_w_2673));
  bfr _b_1490(.a(_w_2306),.q(_w_2307));
  bfr _b_2617(.a(_w_3433),.q(_w_3434));
  spl2 g315_s_1(.a(n315_1),.q0(n315_2),.q1(_w_2370));
  or_bb g397(.a(n393),.b(n396),.q(n397));
  and_bi g398(.a(n384_1),.b(n382_2),.q(n398));
  and_bi g403(.a(n402),.b(n401_0),.q(n403));
  or_bb g411(.a(G9_9),.b(n385_4),.q(n411));
  spl2 g669_s_0(.a(n669),.q0(n669_0),.q1(n669_1));
  bfr _b_1382(.a(_w_2198),.q(n340_1));
  bfr _b_2321(.a(_w_3137),.q(_w_3138));
  or_bb g261(.a(G38_0),.b(n260_0),.q(n261));
  bfr _b_1928(.a(_w_2744),.q(n292));
  bfr _b_2430(.a(_w_3246),.q(_w_3247));
  spl4L g395_s_3(.a(n395_7),.q0(n395_12),.q1(n395_13),.q2(_w_2749),.q3(n395_15));
  and_bi g85(.a(n83),.b(n84),.q(n85));
  bfr _b_1724(.a(_w_2540),.q(_w_2541));
  and_bi g415(.a(n395_9),.b(G8_14),.q(n415));
  spl3L g298_s_0(.a(n298),.q0(n298_0),.q1(n298_1),.q2(n298_2));
  and_bi g420(.a(n392_11),.b(G12_13),.q(n420));
  or_bb g424(.a(n406),.b(n423),.q(n424));
  spl2 G16_s_0(.a(_w_3413),.q0(G16_0),.q1(_w_3221));
  bfr _b_1706(.a(_w_2522),.q(n399));
  or_bb g561(.a(n270_1),.b(n560_0),.q(n561));
  and_bi g425(.a(n424),.b(n381_3),.q(_w_2365));
  bfr _b_1517(.a(_w_2333),.q(_w_2334));
  bfr _b_1331(.a(_w_2147),.q(_w_2148));
  and_bi g152(.a(_w_3464),.b(n151_0),.q(_w_2364));
  spl3L g490_s_0(.a(n490),.q0(n490_0),.q1(n490_1),.q2(n490_2));
  or_bb g511(.a(n508),.b(n510),.q(n511));
  bfr _b_2244(.a(_w_3060),.q(_w_3061));
  and_bi g427(.a(n426),.b(n378),.q(_w_2363));
  or_bb g83(.a(G36_1),.b(G37_1),.q(n83));
  and_bb g490(.a(G47_4),.b(n480_0),.q(n490));
  bfr _b_2241(.a(_w_3057),.q(n686));
  or_bb g430(.a(n379_11),.b(n429),.q(n430));
  spl2 G32_s_1(.a(G32_3),.q0(G32_4),.q1(G32_5));
  and_bb g302(.a(G14_4),.b(G4_30),.q(n302));
  and_bb g644(.a(n377_2),.b(n546_0),.q(n644));
  spl2 g372_s_1(.a(n372_1),.q0(n372_2),.q1(_w_2362));
  bfr _b_1583(.a(_w_2399),.q(_w_2400));
  bfr _b_1867(.a(_w_2683),.q(_w_2684));
  and_bi g482(.a(n436_4),.b(n374_0),.q(n482));
  bfr _b_2667(.a(_w_3483),.q(_w_3484));
  and_bb g649(.a(n646),.b(n648),.q(n649));
  bfr _b_1934(.a(_w_2750),.q(_w_2751));
  spl2 g159_s_0(.a(n159),.q0(n159_0),.q1(n159_1));
  and_bi g448(.a(n447),.b(n445),.q(n448));
  and_bb g450(.a(n444),.b(n449),.q(n450));
  spl2 g100_s_0(.a(n100),.q0(n100_0),.q1(n100_1));
  and_bi g451(.a(n450),.b(n443),.q(n451));
  and_bi g180(.a(G4_26),.b(G30_5),.q(n180));
  spl3L G40_s_1(.a(G40_1),.q0(G40_2),.q1(G40_3),.q2(_w_2361));
  or_bb g824(.a(n814_0),.b(n823),.q(n824));
  or_bb g453(.a(n420_1),.b(n452),.q(n453));
  spl3L g277_s_0(.a(n277),.q0(n277_0),.q1(n277_1),.q2(n277_2));
  and_bi g184(.a(n183),.b(n147_10),.q(n184));
  spl2 g509_s_0(.a(n509),.q0(n509_0),.q1(_w_3400));
  bfr _b_2194(.a(_w_3010),.q(_w_3011));
  and_bi g458(.a(n457),.b(n453),.q(n458));
  and_bi g58(.a(G31_0),.b(G8_0),.q(n58));
  and_bi g460(.a(G14_6),.b(G42_2),.q(n460));
  bfr _b_1380(.a(_w_2196),.q(_w_2197));
  spl3L g533_s_2(.a(n533_3),.q0(n533_4),.q1(n533_5),.q2(_w_2412));
  or_bb g230(.a(n226),.b(n229),.q(n230));
  or_bb g469(.a(n314_1),.b(n337_1),.q(n469));
  bfr _b_2337(.a(_w_3153),.q(n533_1));
  spl2 g147_s_0(.a(n147),.q0(n147_0),.q1(n147_1));
  and_bi g477(.a(n472),.b(n476),.q(_w_2359));
  spl3L g811_s_0(.a(n811),.q0(n811_0),.q1(n811_1),.q2(n811_2));
  bfr _b_2349(.a(_w_3165),.q(_w_3166));
  spl2 G27_s_1(.a(G27_1),.q0(G27_2),.q1(_w_2325));
  or_bb g721(.a(n385_7),.b(n572_1),.q(_w_2324));
  and_bb g476(.a(n473),.b(n475),.q(n476));
  bfr _b_1550(.a(_w_2366),.q(_w_2367));
  and_bi g251(.a(G11_7),.b(n250_0),.q(n251));
  bfr _b_1784(.a(_w_2600),.q(_w_2601));
  and_bi g181(.a(n179_0),.b(n180),.q(n181));
  and_bi g481(.a(G47_5),.b(n480_1),.q(_w_2322));
  spl2 g105_s_1(.a(n105_1),.q0(n105_2),.q1(_w_2983));
  and_bb g378(.a(n369_0),.b(n377_0),.q(n378));
  and_bi g483(.a(n374_3),.b(n215_3),.q(n483));
  bfr _b_1906(.a(_w_2722),.q(_w_2723));
  bfr _b_2130(.a(_w_2946),.q(_w_2947));
  bfr _b_2562(.a(_w_3378),.q(_w_3379));
  spl2 g74_s_0(.a(n74),.q0(_w_2321),.q1(n74_1));
  bfr _b_1915(.a(_w_2731),.q(G33_6));
  and_bi g546(.a(n544),.b(n545),.q(_w_2320));
  and_bb g495(.a(n436_2),.b(n494_3),.q(n495));
  spl2 G9_s_5(.a(G9_12),.q0(G9_13),.q1(G9_14));
  and_bb g499(.a(n190_2),.b(n497_1),.q(n499));
  bfr _b_2585(.a(_w_3401),.q(_w_3402));
  or_bb g813(.a(G3531_1),.b(G3533_1),.q(n813));
  bfr _b_2410(.a(_w_3226),.q(G20_6));
  bfr _b_1641(.a(_w_2457),.q(_w_2458));
  or_bb g503(.a(n240_5),.b(n501_1),.q(n503));
  spl4L G12_s_4(.a(G12_8),.q0(G12_9),.q1(G12_10),.q2(G12_11),.q3(G12_12));
  bfr _b_2300(.a(_w_3116),.q(_w_3117));
  or_bb g319(.a(n306_2),.b(n318),.q(n319));
  and_bb g760(.a(n751),.b(n759),.q(n760));
  or_bb g95(.a(G32_1),.b(G33_1),.q(n95));
  and_bi g258(.a(n256),.b(n257),.q(n258));
  bfr _b_1811(.a(_w_2627),.q(_w_2628));
  spl3L G4_s_3(.a(G4_9),.q0(G4_12),.q1(G4_13),.q2(G4_14));
  bfr _b_1873(.a(_w_2689),.q(_w_2690));
  bfr _b_2731(.a(_w_3547),.q(_w_3548));
  and_bi g508(.a(n237_3),.b(n361_13),.q(_w_2319));
  spl2 G33_s_2(.a(G33_5),.q0(_w_2731),.q1(G33_7));
  and_bi g510(.a(n494_0),.b(n509_0),.q(n510));
  bfr _b_2469(.a(_w_3285),.q(_w_3286));
  bfr _b_2013(.a(_w_2829),.q(_w_2830));
  bfr _b_2263(.a(_w_3079),.q(_w_3080));
  and_bb g515(.a(n507_0),.b(n514_3),.q(n515));
  bfr _b_2215(.a(_w_3031),.q(_w_3032));
  and_bb g736(.a(n437_1),.b(n735_0),.q(n736));
  bfr _b_2129(.a(_w_2945),.q(n601));
  bfr _b_2594(.a(G13),.q(_w_3410));
  or_bb g516(.a(n507_1),.b(n514_4),.q(n516));
  and_bb g518(.a(n505_0),.b(n517_0),.q(n518));
  or_bb g519(.a(n505_1),.b(n517_1),.q(n519));
  and_bi g619(.a(n618),.b(n614),.q(_w_2978));
  or_bb g800(.a(n798),.b(n799),.q(n800));
  spl2 g85_s_0(.a(n85),.q0(n85_0),.q1(n85_1));
  and_bb g522(.a(n521_1),.b(n56_2),.q(_w_2300));
  bfr _b_2604(.a(_w_3420),.q(_w_3413));
  spl3L G12_s_6(.a(G12_15),.q0(G12_16),.q1(G12_17),.q2(G12_18));
  or_bb g78(.a(G35_9),.b(G36_7),.q(n78));
  and_bi g523(.a(n522),.b(n520),.q(n523));
  spl3L g54_s_0(.a(n54),.q0(n54_0),.q1(n54_1),.q2(_w_2296));
  and_bb g756(.a(n753),.b(n755),.q(n756));
  and_bi g528(.a(n74_1),.b(G14_19),.q(n528));
  spl2 G21_s_0(.a(_w_3438),.q0(G21_0),.q1(G21_1));
  spl2 G29_s_0(.a(_w_3467),.q0(G29_0),.q1(_w_2293));
  and_bi g429(.a(n369_2),.b(G47_1),.q(n429));
  and_bi g529(.a(n528),.b(n275_1),.q(_w_2292));
  bfr _b_1922(.a(_w_2738),.q(n186));
  spl4L G31_s_0(.a(_w_3469),.q0(G31_0),.q1(G31_1),.q2(G31_2),.q3(G31_3));
  or_bi g531(.a(n523),.b(n530),.q(_w_2275));
  and_bi g532(.a(n260_3),.b(n125_1),.q(_w_2272));
  and_bi g533(.a(n532),.b(n73_5),.q(_w_2257));
  and_bi g558(.a(n295_2),.b(n361_20),.q(_w_2255));
  spl2 g543_s_0(.a(n543),.q0(n543_0),.q1(n543_1));
  and_bi g534(.a(n340_2),.b(n361_11),.q(n534));
  or_bb g535(.a(n365_0),.b(n534_0),.q(n535));
  bfr _b_2278(.a(_w_3094),.q(_w_3095));
  bfr _b_1663(.a(_w_2479),.q(_w_2480));
  bfr _b_1809(.a(_w_2625),.q(_w_2626));
  bfr _b_1575(.a(_w_2391),.q(_w_2392));
  spl2 G3_s_8(.a(G3_23),.q0(G3_24),.q1(G3_25));
  spl2 g826_s_0(.a(n826),.q0(n826_0),.q1(n826_1));
  spl3L g295_s_0(.a(n295),.q0(n295_0),.q1(n295_1),.q2(_w_2246));
  and_bb g550(.a(n546_3),.b(n548_1),.q(_w_2245));
  spl4L G30_s_0(.a(_w_3468),.q0(G30_0),.q1(G30_1),.q2(G30_2),.q3(_w_2244));
  and_bi g103(.a(n101),.b(n102),.q(_w_2662));
  spl2 G13_s_5(.a(G13_9),.q0(G13_10),.q1(G13_11));
  spl2 G9_s_7(.a(G9_17),.q0(G9_18),.q1(G9_19));
  bfr _b_1455(.a(_w_2271),.q(n533));
  spl4L G7_s_5(.a(G7_14),.q0(G7_15),.q1(G7_16),.q2(G7_17),.q3(G7_18));
  spl4L g151_s_1(.a(n151_3),.q0(n151_4),.q1(n151_5),.q2(n151_6),.q3(n151_7));
  bfr _b_2587(.a(_w_3403),.q(_w_3404));
  or_bb g404(.a(n400),.b(n403),.q(n404));
  or_bb g176(.a(n168),.b(n175),.q(n176));
  bfr _b_2414(.a(_w_3230),.q(n696));
  and_bi g552(.a(n551_1),.b(G3526_3),.q(n552));
  or_bb g775(.a(n773),.b(n774),.q(_w_3108));
  bfr _b_1892(.a(_w_2708),.q(_w_2709));
  bfr _b_2654(.a(G32),.q(_w_3470));
  and_bi g611(.a(n399_1),.b(n401_7),.q(n611));
  and_bi g255(.a(G32_6),.b(n151_2),.q(n255));
  and_bi g341(.a(n143_8),.b(n338_2),.q(n341));
  and_bi g553(.a(G3526_1),.b(n551_0),.q(n553));
  bfr _b_1838(.a(_w_2654),.q(_w_2655));
  or_bb g573(.a(n401_5),.b(n572_0),.q(n573));
  bfr _b_1655(.a(_w_2471),.q(_w_2472));
  spl2 g73_s_1(.a(n73_1),.q0(n73_2),.q1(n73_3));
  bfr _b_1334(.a(_w_2150),.q(n365_2));
  spl2 g73_s_2(.a(n73_3),.q0(n73_4),.q1(n73_5));
  bfr _b_1875(.a(_w_2691),.q(_w_2692));
  bfr _b_2073(.a(_w_2889),.q(_w_2890));
  spl2 g162_s_1(.a(n162_0),.q0(n162_2),.q1(n162_3));
  or_bb g718(.a(n714),.b(n717),.q(_w_2243));
  and_bi g365(.a(n363),.b(n364),.q(n365));
  and_bb g710(.a(G4_46),.b(n409_0),.q(n710));
  bfr _b_1342(.a(_w_2158),.q(_w_2159));
  and_bb g560(.a(n254_2),.b(n361_2),.q(n560));
  or_bb g569(.a(n567),.b(n568),.q(_w_2241));
  and_bi g570(.a(n569),.b(n557),.q(n570));
  and_bb g571(.a(n377_1),.b(n563_0),.q(n571));
  bfr _b_1401(.a(_w_2217),.q(_w_2218));
  bfr _b_1530(.a(_w_2346),.q(_w_2347));
  bfr _b_1674(.a(_w_2490),.q(_w_2491));
  and_bi g714(.a(G16_1),.b(n401_18),.q(n714));
  spl2 G2_s_2(.a(G2_4),.q0(G2_5),.q1(G2_6));
  and_bi g572(.a(G7_3),.b(G19_2),.q(n572));
  bfr _b_2524(.a(_w_3340),.q(_w_3341));
  spl3L g123_s_2(.a(n123_2),.q0(n123_4),.q1(n123_5),.q2(n123_6));
  bfr _b_1924(.a(_w_2740),.q(_w_2741));
  bfr _b_1780(.a(_w_2596),.q(n468));
  and_bb g385(.a(n382_0),.b(n384_0),.q(n385));
  bfr _b_2691(.a(_w_3507),.q(_w_3508));
  bfr _b_1436(.a(_w_2252),.q(_w_2253));
  bfr _b_1478(.a(_w_2294),.q(_w_2295));
  bfr _b_2651(.a(G29),.q(_w_3467));
  spl2 G41_s_0(.a(G41),.q0(G41_0),.q1(_w_2240));
  or_bb g657(.a(n653_0),.b(n656),.q(n657));
  and_bb g382(.a(G25_1),.b(G3_5),.q(n382));
  and_bi g586(.a(n386_1),.b(n401_23),.q(n586));
  or_bb g484(.a(n482_0),.b(n483),.q(n484));
  spl3L g385_s_5(.a(n385_16),.q0(n385_17),.q1(n385_18),.q2(n385_19));
  and_bi g587(.a(G12_14),.b(G40_5),.q(n587));
  bfr _b_1745(.a(_w_2561),.q(G3523));
  spl4L G4_s_4(.a(G4_10),.q0(G4_15),.q1(G4_16),.q2(G4_17),.q3(G4_18));
  and_bi g823(.a(G3532_3),.b(G3528_3),.q(n823));
  spl2 G40_s_3(.a(G40_7),.q0(G40_8),.q1(G40_9));
  or_bb g421(.a(n419_0),.b(n420_0),.q(n421));
  bfr _b_1737(.a(_w_2553),.q(_w_2554));
  or_bb g588(.a(n385_20),.b(n587_0),.q(n588));
  spl4L G7_s_4(.a(G7_10),.q0(G7_11),.q1(G7_12),.q2(G7_13),.q3(G7_14));
  spl4L g293_s_0(.a(n293),.q0(n293_0),.q1(n293_1),.q2(n293_2),.q3(_w_2239));
  spl3L g52_s_0(.a(n52),.q0(n52_0),.q1(n52_1),.q2(n52_2));
  or_bb g487(.a(n379_12),.b(n486),.q(n487));
  spl2 g105_s_2(.a(n105_3),.q0(n105_4),.q1(n105_5));
  spl3L g238_s_0(.a(n238),.q0(n238_0),.q1(n238_1),.q2(n238_2));
  bfr _b_1947(.a(_w_2763),.q(G3528_0));
  bfr _b_2228(.a(_w_3044),.q(_w_3045));
  spl2 g731_s_0(.a(G3534_0),.q0(G3534_1),.q1(G3534_2));
  spl2 g731_s_1(.a(G3534_2),.q0(G3534_3),.q1(_w_2230));
  bfr _b_2698(.a(_w_3514),.q(_w_3495));
  or_bb g525(.a(n105_2),.b(n52_1),.q(n525));
  bfr _b_2142(.a(_w_2958),.q(_w_2959));
  spl4L g250_s_0(.a(n250),.q0(n250_0),.q1(n250_1),.q2(n250_2),.q3(n250_3));
  spl2 g834_s_0(.a(n834),.q0(n834_0),.q1(n834_1));
  bfr _b_2161(.a(_w_2977),.q(n305));
  bfr _b_1621(.a(_w_2437),.q(n377_0));
  and_bi g112(.a(G11_16),.b(G13_19),.q(n112));
  spl2 g834_s_1(.a(n834_1),.q0(n834_2),.q1(_w_2228));
  spl2 g563_s_1(.a(n563_1),.q0(n563_2),.q1(n563_3));
  spl2 g265_s_2(.a(n265_3),.q0(n265_4),.q1(n265_5));
  bfr _b_1943(.a(_w_2759),.q(_w_2760));
  bfr _b_2070(.a(_w_2886),.q(_w_2887));
  spl4L g407_s_1(.a(n407_2),.q0(n407_4),.q1(n407_5),.q2(n407_6),.q3(n407_7));
  bfr _b_1348(.a(_w_2164),.q(_w_2165));
  spl4L g407_s_2(.a(n407_3),.q0(n407_8),.q1(n407_9),.q2(n407_10),.q3(n407_11));
  spl2 g282_s_1(.a(n282_1),.q0(n282_2),.q1(_w_2227));
  bfr _b_2575(.a(_w_3391),.q(n536));
  and_bb g464(.a(n458),.b(n463),.q(n464));
  spl2 g384_s_0(.a(n384),.q0(n384_0),.q1(n384_1));
  bfr _b_1973(.a(_w_2789),.q(_w_2790));
  spl4L g283_s_0(.a(n283),.q0(n283_0),.q1(n283_1),.q2(n283_2),.q3(_w_2225));
  spl2 g822_s_0(.a(n822),.q0(n822_0),.q1(n822_1));
  spl2 g491_s_0(.a(n491),.q0(n491_0),.q1(n491_1));
  spl2 G7_s_0(.a(_w_3570),.q0(G7_0),.q1(_w_2222));
  bfr _b_1713(.a(_w_2529),.q(_w_2530));
  spl4L G7_s_3(.a(G7_6),.q0(G7_7),.q1(G7_8),.q2(G7_9),.q3(G7_10));
  spl2 G7_s_6(.a(G7_18),.q0(G7_19),.q1(G7_20));
  bfr _b_1388(.a(_w_2204),.q(n260_3));
  and_bb g123(.a(G3_4),.b(n73_0),.q(n123));
  or_bb g335(.a(n333),.b(n334),.q(n335));
  bfr _b_1700(.a(_w_2516),.q(_w_2517));
  spl2 g372_s_0(.a(n372),.q0(n372_0),.q1(_w_2211));
  spl2 g372_s_2(.a(n372_3),.q0(n372_4),.q1(n372_5));
  bfr _b_2597(.a(G16),.q(_w_3414));
  spl2 g351_s_0(.a(n351),.q0(n351_0),.q1(n351_1));
  spl2 g372_s_4(.a(n372_7),.q0(n372_8),.q1(n372_9));
  spl3L g372_s_5(.a(n372_9),.q0(n372_10),.q1(n372_11),.q2(n372_12));
  bfr _b_2368(.a(_w_3184),.q(_w_3185));
  spl2 g408_s_0(.a(n408),.q0(n408_0),.q1(n408_1));
  spl2 G22_s_0(.a(_w_3443),.q0(G22_0),.q1(_w_2210));
  bfr _b_2095(.a(_w_2911),.q(_w_2912));
  bfr _b_2515(.a(_w_3331),.q(_w_3332));
  spl2 G22_s_1(.a(G22_1),.q0(G22_2),.q1(_w_2209));
  bfr _b_2736(.a(_w_3552),.q(_w_3553));
  bfr _b_2252(.a(_w_3068),.q(n399_1));
  spl3L G22_s_2(.a(G22_3),.q0(G22_4),.q1(G22_5),.q2(G22_6));
  spl3L G22_s_3(.a(G22_6),.q0(G22_7),.q1(G22_8),.q2(_w_2208));
  spl4L g398_s_1(.a(n398_3),.q0(n398_4),.q1(n398_5),.q2(n398_6),.q3(n398_7));
  or_bb g579(.a(n385_12),.b(n578),.q(n579));
  bfr _b_1964(.a(_w_2780),.q(_w_2781));
  spl2 g732_s_0(.a(n732),.q0(n732_0),.q1(n732_1));
  spl4L g398_s_5(.a(n398_15),.q0(n398_18),.q1(n398_19),.q2(n398_20),.q3(n398_21));
  bfr _b_2519(.a(_w_3335),.q(_w_3336));
  bfr _b_2152(.a(_w_2968),.q(_w_2969));
  spl4L g407_s_0(.a(n407),.q0(n407_0),.q1(n407_1),.q2(n407_2),.q3(n407_3));
  spl2 g306_s_0(.a(n306),.q0(n306_0),.q1(n306_1));
  bfr _b_1356(.a(_w_2172),.q(_w_2173));
  and_bi g493(.a(n491_1),.b(n238_2),.q(n493));
  spl2 g306_s_1(.a(n306_1),.q0(n306_2),.q1(_w_2207));
  spl3L g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1),.q2(_w_2205));
  bfr _b_1937(.a(_w_2753),.q(_w_2754));
  bfr _b_1353(.a(_w_2169),.q(_w_2170));
  bfr _b_2614(.a(_w_3430),.q(_w_3431));
  spl4L g260_s_0(.a(n260),.q0(n260_0),.q1(n260_1),.q2(n260_2),.q3(_w_2202));
  bfr _b_1338(.a(_w_2154),.q(_w_2155));
  spl3L g320_s_0(.a(n320),.q0(n320_0),.q1(n320_1),.q2(n320_2));
  bfr _b_2607(.a(_w_3423),.q(_w_3424));
  spl2 g320_s_1(.a(n320_2),.q0(n320_3),.q1(_w_2200));
  spl2 g329_s_0(.a(n329),.q0(n329_0),.q1(n329_1));
  or_bb g840(.a(n832_1),.b(n838_1),.q(n840));
  spl2 G8_s_1(.a(G8_1),.q0(G8_2),.q1(G8_3));
  and_bi g769(.a(n768),.b(n533_8),.q(n769));
  spl2 g383_s_0(.a(n383),.q0(n383_0),.q1(n383_1));
  spl2 G8_s_4(.a(G8_7),.q0(G8_8),.q1(G8_9));
  bfr _b_1336(.a(_w_2152),.q(_w_2153));
  spl2 g481_s_0(.a(n481),.q0(n481_0),.q1(n481_1));
  spl2 G8_s_6(.a(G8_13),.q0(G8_14),.q1(G8_15));
  bfr _b_1628(.a(_w_2444),.q(_w_2445));
  bfr _b_2179(.a(_w_2995),.q(n511_1));
  or_bb g730(.a(n702),.b(n729),.q(n730));
  spl3L g338_s_0(.a(n338),.q0(n338_0),.q1(n338_1),.q2(_w_2199));
  spl2 g420_s_0(.a(n420),.q0(n420_0),.q1(n420_1));
  bfr _b_2566(.a(_w_3382),.q(_w_3383));
  spl2 g682_s_0(.a(G3533_0),.q0(G3533_1),.q1(G3533_2));
  spl2 g340_s_0(.a(n340),.q0(n340_0),.q1(_w_2196));
  and_bi g440(.a(n392_14),.b(G8_16),.q(n440));
  spl2 g340_s_1(.a(n340_1),.q0(n340_2),.q1(_w_2194));
  spl2 G19_s_0(.a(G19),.q0(G19_0),.q1(_w_2190));
  spl2 G19_s_1(.a(G19_1),.q0(G19_2),.q1(_w_2188));
  spl2 G19_s_2(.a(G19_3),.q0(G19_4),.q1(_w_2187));
  bfr _b_1768(.a(_w_2584),.q(_w_2585));
  spl3L g385_s_0(.a(n385),.q0(_w_2186),.q1(n385_1),.q2(n385_2));
  bfr _b_1433(.a(_w_2249),.q(_w_2250));
  bfr _b_2160(.a(_w_2976),.q(n608));
  and_bi g715(.a(G17_2),.b(n398_9),.q(n715));
  spl3L g365_s_0(.a(n365),.q0(n365_0),.q1(n365_1),.q2(_w_2145));
  spl2 g366_s_0(.a(n366),.q0(n366_0),.q1(n366_1));
  and_bi g194(.a(G10_14),.b(n193),.q(n194));
  spl2 g374_s_1(.a(n374_2),.q0(n374_3),.q1(n374_4));
  bfr _b_1354(.a(_w_2170),.q(_w_2171));
  spl2 g374_s_3(.a(n374_6),.q0(n374_7),.q1(n374_8));
  bfr _b_1905(.a(_w_2721),.q(_w_2722));
  bfr _b_2009(.a(_w_2825),.q(_w_2826));
  spl4L g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1),.q2(n379_2),.q3(n379_3));
  spl3L g379_s_1(.a(n379_2),.q0(n379_4),.q1(n379_5),.q2(n379_6));
  and_bi g577(.a(n573),.b(n576),.q(n577));
  spl2 g237_s_1(.a(n237_1),.q0(n237_2),.q1(_w_2142));
  bfr _b_2060(.a(_w_2876),.q(_w_2877));
  spl2 G24_s_1(.a(G24_1),.q0(G24_2),.q1(_w_2137));
  or_bb g281(.a(n276),.b(n280),.q(n281));
  spl2 G24_s_2(.a(G24_3),.q0(G24_4),.q1(G24_5));
  bfr _b_1978(.a(_w_2794),.q(_w_2795));
  spl2 G24_s_3(.a(G24_5),.q0(G24_6),.q1(_w_2136));
  bfr _b_2112(.a(_w_2928),.q(_w_2929));
  bfr _b_1383(.a(_w_2199),.q(n338_2));
  spl4L g385_s_1(.a(n385_1),.q0(n385_3),.q1(n385_4),.q2(n385_5),.q3(n385_6));
  spl4L g385_s_2(.a(n385_2),.q0(n385_7),.q1(n385_8),.q2(n385_9),.q3(n385_10));
  spl4L G4_s_0(.a(G4),.q0(G4_0),.q1(G4_1),.q2(G4_2),.q3(G4_3));
  spl2 g385_s_3(.a(n385_9),.q0(n385_11),.q1(n385_12));
  spl4L g385_s_4(.a(n385_10),.q0(n385_13),.q1(n385_14),.q2(n385_15),.q3(n385_16));
  spl2 g385_s_6(.a(n385_19),.q0(n385_20),.q1(n385_21));
  bfr _b_2716(.a(_w_3532),.q(_w_3533));
  bfr _b_2565(.a(_w_3381),.q(_w_3382));
  bfr _b_1954(.a(_w_2770),.q(_w_2771));
  bfr _b_2022(.a(_w_2838),.q(G1_13));
  spl4L g401_s_0(.a(n401),.q0(n401_0),.q1(n401_1),.q2(n401_2),.q3(n401_3));
  and_bi g808(.a(n533_5),.b(n695_2),.q(n808));
  spl4L g401_s_1(.a(n401_2),.q0(n401_4),.q1(n401_5),.q2(n401_6),.q3(n401_7));
  bfr _b_2358(.a(_w_3174),.q(_w_3175));
  spl4L g401_s_3(.a(n401_11),.q0(n401_12),.q1(n401_13),.q2(n401_14),.q3(n401_15));
  and_bi g314(.a(n313),.b(n147_7),.q(n314));
  spl3L g401_s_4(.a(n401_14),.q0(n401_16),.q1(n401_17),.q2(n401_18));
  bfr _b_2737(.a(_w_3553),.q(_w_3554));
  spl2 g401_s_6(.a(n401_22),.q0(n401_23),.q1(n401_24));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(n119_1));
  or_bb g801(.a(n797),.b(n800),.q(n801));
  or_bb g443(.a(n439),.b(n442),.q(n443));
  spl3L g437_s_0(.a(n437),.q0(n437_0),.q1(n437_1),.q2(n437_2));
  spl2 g437_s_1(.a(n437_2),.q0(n437_3),.q1(n437_4));
  spl2 g411_s_0(.a(n411),.q0(n411_0),.q1(n411_1));
  spl2 g433_s_0(.a(n433),.q0(n433_0),.q1(n433_1));
  spl2 g436_s_0(.a(n436),.q0(n436_0),.q1(_w_2134));
  and_bi g326(.a(n227_1),.b(n325),.q(n326));
  bfr _b_2168(.a(_w_2984),.q(_w_2985));
  spl3L G4_s_10(.a(G4_35),.q0(G4_36),.q1(_w_2840),.q2(G4_38));
  and_bi g205(.a(G4_12),.b(G32_4),.q(n205));
  bfr _b_1686(.a(_w_2502),.q(n145));
  spl2 g436_s_2(.a(n436_3),.q0(n436_4),.q1(_w_2131));
  bfr _b_1524(.a(_w_2340),.q(_w_2341));
  spl2 g51_s_2(.a(n51_3),.q0(n51_4),.q1(_w_2130));
  bfr _b_1825(.a(_w_2641),.q(_w_2642));
  and_bi g422(.a(n417),.b(n421),.q(n422));
  spl3L g496_s_0(.a(n496),.q0(n496_0),.q1(n496_1),.q2(n496_2));
  bfr _b_1914(.a(_w_2730),.q(G18_1));
  spl3L g189_s_0(.a(n189),.q0(n189_0),.q1(n189_1),.q2(n189_2));
  spl2 g267_s_0(.a(n267),.q0(n267_0),.q1(_w_2129));
  bfr _b_1512(.a(_w_2328),.q(_w_2329));
  and_bb g347(.a(n299_1),.b(n317_2),.q(n347));
  spl2 g482_s_0(.a(n482),.q0(n482_0),.q1(n482_1));
  bfr _b_1863(.a(_w_2679),.q(_w_2680));
  spl2 G42_s_1(.a(G42_1),.q0(G42_2),.q1(G42_3));
  bfr _b_1520(.a(_w_2336),.q(_w_2337));
  spl3L g695_s_0(.a(n695),.q0(n695_0),.q1(n695_1),.q2(n695_2));
  spl3L g494_s_0(.a(n494),.q0(n494_0),.q1(n494_1),.q2(_w_2127));
  bfr _b_1440(.a(_w_2256),.q(n558));
  spl2 g494_s_1(.a(n494_2),.q0(n494_3),.q1(_w_2122));
  spl2 G13_s_2(.a(G13_3),.q0(G13_4),.q1(G13_5));
  spl2 G13_s_3(.a(G13_5),.q0(G13_6),.q1(G13_7));
  spl3L G13_s_7(.a(G13_14),.q0(G13_15),.q1(G13_16),.q2(G13_17));
  spl4L g143_s_1(.a(n143_1),.q0(n143_2),.q1(n143_3),.q2(n143_4),.q3(n143_5));
  bfr _b_2538(.a(_w_3354),.q(_w_3355));
  spl3L g270_s_0(.a(n270),.q0(n270_0),.q1(n270_1),.q2(n270_2));
  spl4L g143_s_2(.a(n143_5),.q0(n143_6),.q1(n143_7),.q2(n143_8),.q3(n143_9));
  bfr _b_2454(.a(_w_3270),.q(_w_3271));
  bfr _b_2390(.a(_w_3206),.q(_w_3207));
  spl2 g500_s_1(.a(n500_1),.q0(n500_2),.q1(n500_3));
  spl2 g500_s_2(.a(n500_3),.q0(n500_4),.q1(_w_2121));
  and_bi g67(.a(G33_0),.b(G10_0),.q(n67));
  bfr _b_1371(.a(_w_2187),.q(G19_5));
  and_bi g799(.a(G20_3),.b(n385_8),.q(n799));
  spl3L g507_s_0(.a(n507),.q0(n507_0),.q1(n507_1),.q2(_w_2120));
  spl2 g512_s_0(.a(n512),.q0(n512_0),.q1(n512_1));
  bfr _b_1691(.a(_w_2507),.q(n750));
  bfr _b_2119(.a(_w_2935),.q(_w_2936));
  spl2 G13_s_4(.a(G13_7),.q0(G13_8),.q1(G13_9));
  spl2 g514_s_1(.a(n514_2),.q0(n514_3),.q1(n514_4));
  bfr _b_1748(.a(_w_2564),.q(n372_7));
  spl4L g215_s_0(.a(n215),.q0(n215_0),.q1(n215_1),.q2(n215_2),.q3(_w_2111));
  or_bb g282(.a(n273),.b(n281),.q(n282));
  bfr _b_1409(.a(_w_2225),.q(_w_2226));
  and_bb g742(.a(G17_0),.b(n395_2),.q(n742));
  spl2 g521_s_0(.a(n521),.q0(n521_0),.q1(n521_1));
  bfr _b_1296(.a(_w_2112),.q(_w_2113));
  bfr _b_1297(.a(_w_2113),.q(_w_2114));
  bfr _b_1299(.a(_w_2115),.q(_w_2116));
  bfr _b_2116(.a(_w_2932),.q(_w_2933));
  spl2 g233_s_0(.a(n233),.q0(n233_0),.q1(n233_1));
  bfr _b_1303(.a(_w_2119),.q(n215_3));
  spl2 G23_s_0(.a(_w_3446),.q0(G23_0),.q1(_w_3227));
  bfr _b_1851(.a(_w_2667),.q(_w_2668));
  bfr _b_1304(.a(_w_2120),.q(n507_2));
  and_bi g488(.a(n485),.b(n487),.q(n488));
  bfr _b_2123(.a(_w_2939),.q(G3529));
  bfr _b_2631(.a(_w_3447),.q(_w_3448));
  bfr _b_1306(.a(_w_2122),.q(_w_2123));
  bfr _b_1307(.a(_w_2123),.q(_w_2124));
  bfr _b_1890(.a(_w_2706),.q(n72));
  bfr _b_1308(.a(_w_2124),.q(_w_2125));
  bfr _b_1311(.a(_w_2127),.q(_w_2128));
  bfr _b_1397(.a(_w_2213),.q(_w_2214));
  bfr _b_1312(.a(_w_2128),.q(n494_2));
  and_bi g669(.a(G13_10),.b(G41_5),.q(n669));
  bfr _b_2207(.a(_w_3023),.q(_w_3024));
  bfr _b_2006(.a(_w_2822),.q(_w_2823));
  bfr _b_1314(.a(_w_2130),.q(n51_5));
  bfr _b_1897(.a(_w_2713),.q(_w_2714));
  bfr _b_1317(.a(_w_2133),.q(n436_3));
  spl2 g360_s_0(.a(n360),.q0(n360_0),.q1(_w_2151));
  bfr _b_1525(.a(_w_2341),.q(_w_2342));
  bfr _b_1320(.a(_w_2136),.q(G24_7));
  bfr _b_1899(.a(_w_2715),.q(_w_2716));
  bfr _b_1321(.a(_w_2137),.q(_w_2138));
  bfr _b_1322(.a(_w_2138),.q(_w_2139));
  bfr _b_1669(.a(_w_2485),.q(_w_2486));
  bfr _b_2502(.a(_w_3318),.q(_w_3319));
  bfr _b_1810(.a(_w_2626),.q(_w_2627));
  bfr _b_1323(.a(_w_2139),.q(G24_3));
  bfr _b_1370(.a(_w_2186),.q(n385_0));
  bfr _b_1324(.a(_w_2140),.q(_w_2141));
  bfr _b_1325(.a(_w_2141),.q(G24_1));
  bfr _b_1326(.a(_w_2142),.q(_w_2143));
  bfr _b_1772(.a(_w_2588),.q(_w_2589));
  bfr _b_1329(.a(_w_2145),.q(_w_2146));
  or_bb g678(.a(n372_4),.b(n604_1),.q(n678));
  bfr _b_1330(.a(_w_2146),.q(_w_2147));
  bfr _b_1333(.a(_w_2149),.q(_w_2150));
  bfr _b_1488(.a(_w_2304),.q(_w_2305));
  bfr _b_2708(.a(G49),.q(_w_3524));
  bfr _b_1335(.a(_w_2151),.q(_w_2152));
  bfr _b_1337(.a(_w_2153),.q(_w_2154));
  bfr _b_1341(.a(_w_2157),.q(_w_2158));
  bfr _b_1626(.a(_w_2442),.q(_w_2443));
  bfr _b_2505(.a(_w_3321),.q(_w_3322));
  bfr _b_2143(.a(_w_2959),.q(n602));
  bfr _b_1343(.a(_w_2159),.q(_w_2160));
  bfr _b_2385(.a(_w_3201),.q(n224_2));
  bfr _b_1393(.a(_w_2209),.q(G22_3));
  bfr _b_1451(.a(_w_2267),.q(_w_2268));
  spl4L G33_s_0(.a(_w_3471),.q0(G33_0),.q1(G33_1),.q2(G33_2),.q3(G33_3));
  bfr _b_2251(.a(_w_3067),.q(n700));
  bfr _b_1345(.a(_w_2161),.q(_w_2162));
  bfr _b_1460(.a(_w_2276),.q(_w_2277));
  bfr _b_2021(.a(_w_2837),.q(_w_2838));
  bfr _b_1715(.a(_w_2531),.q(_w_2532));
  bfr _b_1346(.a(_w_2162),.q(_w_2163));
  bfr _b_2206(.a(_w_3022),.q(_w_3023));
  bfr _b_1347(.a(_w_2163),.q(_w_2164));
  bfr _b_2423(.a(_w_3239),.q(_w_3240));
  bfr _b_1349(.a(_w_2165),.q(_w_2166));
  bfr _b_1350(.a(_w_2166),.q(_w_2167));
  bfr _b_1355(.a(_w_2171),.q(_w_2172));
  and_bi g537(.a(n535_0),.b(n536),.q(n537));
  bfr _b_1660(.a(_w_2476),.q(_w_2477));
  spl2 g374_s_2(.a(n374_4),.q0(n374_5),.q1(n374_6));
  bfr _b_1357(.a(_w_2173),.q(_w_2174));
  bfr _b_1358(.a(_w_2174),.q(_w_2175));
  and_bi g480(.a(n478),.b(n479),.q(n480));
  bfr _b_1359(.a(_w_2175),.q(_w_2176));
  or_bb g412(.a(G7_12),.b(n398_13),.q(n412));
  bfr _b_1834(.a(_w_2650),.q(n146_1));
  and_bi g418(.a(G22_4),.b(n401_4),.q(n418));
  bfr _b_1361(.a(_w_2177),.q(_w_2178));
  bfr _b_1518(.a(_w_2334),.q(_w_2335));
  bfr _b_2203(.a(_w_3019),.q(_w_3020));
  bfr _b_1365(.a(_w_2181),.q(_w_2182));
  bfr _b_2327(.a(_w_3143),.q(_w_3144));
  or_bb g291(.a(n285),.b(n290),.q(n291));
  bfr _b_1639(.a(_w_2455),.q(_w_2456));
  bfr _b_2646(.a(_w_3462),.q(_w_3463));
  bfr _b_1368(.a(_w_2184),.q(_w_2185));
  bfr _b_1369(.a(_w_2185),.q(n360_1));
  bfr _b_1707(.a(_w_2523),.q(_w_2524));
  and_bb g835(.a(G50_1),.b(n834_2),.q(n835));
  bfr _b_1492(.a(_w_2308),.q(_w_2309));
  bfr _b_1372(.a(_w_2188),.q(_w_2189));
  bfr _b_1771(.a(_w_2587),.q(_w_2588));
  bfr _b_1374(.a(_w_2190),.q(_w_2191));
  bfr _b_1375(.a(_w_2191),.q(_w_2192));
  bfr _b_1413(.a(_w_2229),.q(n834_3));
  spl2 g489_s_1(.a(G3529_2),.q0(G3529_3),.q1(_w_2932));
  bfr _b_1376(.a(_w_2192),.q(_w_2193));
  bfr _b_1428(.a(_w_2244),.q(G30_3));
  bfr _b_1377(.a(_w_2193),.q(G19_1));
  bfr _b_1378(.a(_w_2194),.q(_w_2195));
  bfr _b_1385(.a(_w_2201),.q(n320_4));
  bfr _b_1477(.a(_w_2293),.q(_w_2294));
  bfr _b_1386(.a(_w_2202),.q(_w_2203));
  bfr _b_1389(.a(_w_2205),.q(_w_2206));
  bfr _b_1396(.a(_w_2212),.q(_w_2213));
  bfr _b_1399(.a(_w_2215),.q(_w_2216));
  bfr _b_1864(.a(_w_2680),.q(_w_2681));
  bfr _b_1402(.a(_w_2218),.q(_w_2219));
  bfr _b_1403(.a(_w_2219),.q(_w_2220));
  bfr _b_2271(.a(_w_3087),.q(n688));
  bfr _b_1404(.a(_w_2220),.q(_w_2221));
  bfr _b_1635(.a(_w_2451),.q(n158));
  and_bi g369(.a(n367),.b(n368),.q(_w_2613));
  bfr _b_1405(.a(_w_2221),.q(n372_1));
  bfr _b_1795(.a(_w_2611),.q(_w_2612));
  bfr _b_1407(.a(_w_2223),.q(_w_2224));
  and_bi g68(.a(G30_0),.b(G7_0),.q(n68));
  bfr _b_2284(.a(_w_3100),.q(_w_3101));
  bfr _b_1410(.a(_w_2226),.q(n283_3));
  bfr _b_1411(.a(_w_2227),.q(n282_3));
  bfr _b_1571(.a(_w_2387),.q(_w_2388));
  and_bi g248(.a(G4_24),.b(G1_8),.q(n248));
  bfr _b_1417(.a(_w_2233),.q(_w_2234));
  bfr _b_1419(.a(_w_2235),.q(_w_2236));
  bfr _b_1420(.a(_w_2236),.q(_w_2237));
  or_bb g640(.a(n606),.b(n639),.q(_w_2993));
  spl2 g73_s_0(.a(n73),.q0(n73_0),.q1(_w_2903));
  bfr _b_1673(.a(_w_2489),.q(_w_2490));
  bfr _b_1426(.a(_w_2242),.q(n569));
  bfr _b_1427(.a(_w_2243),.q(n718));
  spl4L g77_s_0(.a(n77),.q0(n77_0),.q1(n77_1),.q2(n77_2),.q3(n77_3));
  bfr _b_1429(.a(_w_2245),.q(n550));
  bfr _b_2656(.a(G34),.q(_w_3472));
  bfr _b_1430(.a(_w_2246),.q(_w_2247));
  bfr _b_1437(.a(_w_2253),.q(_w_2254));
  bfr _b_2706(.a(_w_3522),.q(_w_3523));
  bfr _b_2366(.a(_w_3182),.q(G3535));
  bfr _b_1438(.a(_w_2254),.q(n295_2));
  bfr _b_1443(.a(_w_2259),.q(_w_2260));
  bfr _b_1444(.a(_w_2260),.q(_w_2261));
  bfr _b_2287(.a(_w_3103),.q(_w_3104));
  bfr _b_1446(.a(_w_2262),.q(_w_2263));
  bfr _b_1447(.a(_w_2263),.q(_w_2264));
  bfr _b_2445(.a(_w_3261),.q(G3529_2));
  bfr _b_1448(.a(_w_2264),.q(_w_2265));
  and_bb g608(.a(G39_6),.b(n392_5),.q(_w_2976));
  bfr _b_1676(.a(_w_2492),.q(_w_2493));
  and_bi g165(.a(n161_0),.b(n164_0),.q(n165));
  bfr _b_1449(.a(_w_2265),.q(_w_2266));
  bfr _b_2315(.a(_w_3131),.q(G3538));
  bfr _b_1450(.a(_w_2266),.q(_w_2267));
  bfr _b_1452(.a(_w_2268),.q(_w_2269));
  bfr _b_1453(.a(_w_2269),.q(_w_2270));
  bfr _b_2586(.a(_w_3402),.q(_w_3403));
  bfr _b_1756(.a(_w_2572),.q(_w_2573));
  bfr _b_1454(.a(_w_2270),.q(_w_2271));
  bfr _b_1886(.a(_w_2702),.q(_w_2703));
  bfr _b_2316(.a(_w_3132),.q(G8_5));
  bfr _b_1456(.a(_w_2272),.q(_w_2273));
  bfr _b_2267(.a(_w_3083),.q(n743));
  spl3L g381_s_0(.a(n381),.q0(n381_0),.q1(n381_1),.q2(n381_2));
  bfr _b_1458(.a(_w_2274),.q(n532));
  bfr _b_2664(.a(G40),.q(_w_3481));
  bfr _b_1755(.a(_w_2571),.q(_w_2572));
  spl2 G24_s_0(.a(G24),.q0(G24_0),.q1(_w_2140));
  bfr _b_1459(.a(_w_2275),.q(_w_2276));
  bfr _b_1462(.a(_w_2278),.q(_w_2279));
  spl2 g176_s_1(.a(n176_1),.q0(n176_2),.q1(_w_3256));
  and_bi g437(.a(G4_52),.b(G2_8),.q(_w_2571));
  or_bb g811(.a(G3534_1),.b(G3535_1),.q(n811));
  bfr _b_2212(.a(_w_3028),.q(_w_3029));
  bfr _b_1463(.a(_w_2279),.q(_w_2280));
  bfr _b_1826(.a(_w_2642),.q(_w_2643));
  bfr _b_1465(.a(_w_2281),.q(_w_2282));
  bfr _b_1466(.a(_w_2282),.q(_w_2283));
  bfr _b_2069(.a(_w_2885),.q(_w_2886));
  bfr _b_1734(.a(_w_2550),.q(_w_2551));
  or_bb g556(.a(n542_1),.b(n555),.q(n556));
  bfr _b_1468(.a(_w_2284),.q(_w_2285));
  spl3L G39_s_2(.a(G39_4),.q0(G39_5),.q1(G39_6),.q2(G39_7));
  bfr _b_1469(.a(_w_2285),.q(_w_2286));
  and_bi g73(.a(G2_0),.b(G1_0),.q(n73));
  bfr _b_1470(.a(_w_2286),.q(_w_2287));
  bfr _b_2242(.a(_w_3058),.q(_w_3059));
  bfr _b_1472(.a(_w_2288),.q(_w_2289));
  bfr _b_2181(.a(_w_2997),.q(n645));
  bfr _b_2498(.a(_w_3314),.q(_w_3315));
  spl2 g105_s_0(.a(n105),.q0(n105_0),.q1(_w_2565));
  bfr _b_1473(.a(_w_2289),.q(_w_2290));
  bfr _b_1785(.a(_w_2601),.q(_w_2602));
  bfr _b_1475(.a(_w_2291),.q(G3530));
  bfr _b_2572(.a(_w_3388),.q(_w_3389));
  bfr _b_1476(.a(_w_2292),.q(n529));
  bfr _b_1479(.a(_w_2295),.q(G29_1));
  bfr _b_1480(.a(_w_2296),.q(_w_2297));
  bfr _b_2238(.a(_w_3054),.q(G3533_0));
  bfr _b_2276(.a(_w_3092),.q(_w_3093));
  bfr _b_2632(.a(_w_3448),.q(_w_3449));
  bfr _b_2356(.a(_w_3172),.q(G31_7));
  and_bb g433(.a(n201_3),.b(n361_5),.q(n433));
  bfr _b_1483(.a(_w_2299),.q(n54_2));
  bfr _b_1911(.a(_w_2727),.q(_w_2728));
  and_bb g713(.a(n705),.b(n712),.q(n713));
  bfr _b_1485(.a(_w_2301),.q(_w_2302));
  bfr _b_1487(.a(_w_2303),.q(_w_2304));
  bfr _b_1489(.a(_w_2305),.q(_w_2306));
  bfr _b_1491(.a(_w_2307),.q(_w_2308));
  bfr _b_1881(.a(_w_2697),.q(_w_2698));
  bfr _b_1494(.a(_w_2310),.q(_w_2311));
  bfr _b_1495(.a(_w_2311),.q(_w_2312));
  bfr _b_1497(.a(_w_2313),.q(_w_2314));
  bfr _b_1499(.a(_w_2315),.q(_w_2316));
  bfr _b_1883(.a(_w_2699),.q(_w_2700));
  bfr _b_2376(.a(_w_3192),.q(_w_3193));
  bfr _b_2254(.a(_w_3070),.q(_w_3071));
  bfr _b_1502(.a(_w_2318),.q(n522));
  bfr _b_1503(.a(_w_2319),.q(n508));
  bfr _b_2051(.a(_w_2867),.q(_w_2868));
  bfr _b_1505(.a(_w_2321),.q(n74_0));
  bfr _b_2702(.a(_w_3518),.q(_w_3519));
  bfr _b_1506(.a(_w_2322),.q(_w_2323));
  bfr _b_1508(.a(_w_2324),.q(n721));
  bfr _b_2747(.a(_w_3563),.q(_w_3564));
  and_bi g763(.a(n379_1),.b(n762),.q(_w_2423));
  bfr _b_1956(.a(_w_2772),.q(_w_2773));
  bfr _b_1511(.a(_w_2327),.q(_w_2328));
  bfr _b_1513(.a(_w_2329),.q(_w_2330));
  bfr _b_2086(.a(_w_2902),.q(G42_1));
  spl2 g265_s_0(.a(n265),.q0(n265_0),.q1(n265_1));
  bfr _b_1514(.a(_w_2330),.q(_w_2331));
  bfr _b_1516(.a(_w_2332),.q(_w_2333));
  or_bb g456(.a(n385_17),.b(n455_0),.q(n456));
  bfr _b_1519(.a(_w_2335),.q(_w_2336));
  bfr _b_1521(.a(_w_2337),.q(_w_2338));
  bfr _b_2234(.a(_w_3050),.q(n677));
  bfr _b_1523(.a(_w_2339),.q(_w_2340));
  bfr _b_1526(.a(_w_2342),.q(_w_2343));
  bfr _b_1528(.a(_w_2344),.q(_w_2345));
  bfr _b_1541(.a(_w_2357),.q(_w_2358));
  bfr _b_2528(.a(_w_3344),.q(_w_3345));
  and_bi g390(.a(n389),.b(n387),.q(n390));
  bfr _b_1533(.a(_w_2349),.q(_w_2350));
  or_bb g613(.a(n611),.b(n612),.q(_w_2503));
  bfr _b_1534(.a(_w_2350),.q(_w_2351));
  or_bb g376(.a(n373),.b(n375),.q(_w_2960));
  bfr _b_1538(.a(_w_2354),.q(_w_2355));
  bfr _b_2038(.a(_w_2854),.q(_w_2855));
  bfr _b_1802(.a(_w_2618),.q(n467));
  and_bi g496(.a(G27_2),.b(n77_2),.q(n496));
  bfr _b_1539(.a(_w_2355),.q(_w_2356));
  bfr _b_1604(.a(_w_2420),.q(_w_2421));
  bfr _b_1540(.a(_w_2356),.q(_w_2357));
  bfr _b_1542(.a(_w_2358),.q(G27_3));
  bfr _b_1576(.a(_w_2392),.q(_w_2393));
  bfr _b_2428(.a(_w_3244),.q(_w_3245));
  and_bb g352(.a(n240_0),.b(n351_0),.q(n352));
  bfr _b_1545(.a(_w_2361),.q(G40_4));
  bfr _b_1546(.a(_w_2362),.q(n372_3));
  and_bi g188(.a(n162_3),.b(n185_0),.q(n188));
  bfr _b_1547(.a(_w_2363),.q(n427));
  bfr _b_1549(.a(_w_2365),.q(_w_2366));
  bfr _b_1551(.a(_w_2367),.q(n425));
  spl2 G3_s_4(.a(G3_11),.q0(G3_12),.q1(G3_13));
  bfr _b_1871(.a(_w_2687),.q(_w_2688));
  bfr _b_2028(.a(_w_2844),.q(_w_2845));
  bfr _b_1552(.a(_w_2368),.q(_w_2369));
  bfr _b_1366(.a(_w_2182),.q(_w_2183));
  bfr _b_1554(.a(_w_2370),.q(n315_3));
  bfr _b_1605(.a(_w_2421),.q(n809));
  bfr _b_1962(.a(_w_2778),.q(_w_2779));
  bfr _b_1555(.a(_w_2371),.q(_w_2372));
  spl4L g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1),.q2(n192_2),.q3(_w_2438));
  bfr _b_1556(.a(_w_2372),.q(_w_2373));
  bfr _b_1558(.a(_w_2374),.q(_w_2375));
  bfr _b_1559(.a(_w_2375),.q(_w_2376));
  bfr _b_1561(.a(_w_2377),.q(_w_2378));
  bfr _b_2066(.a(_w_2882),.q(n466));
  bfr _b_1562(.a(_w_2378),.q(_w_2379));
  bfr _b_1565(.a(_w_2381),.q(n372));
  or_bb g472(.a(n293_1),.b(n471),.q(_w_3393));
  bfr _b_1566(.a(_w_2382),.q(_w_2383));
  spl4L g147_s_1(.a(n147_1),.q0(_w_2816),.q1(_w_2817),.q2(_w_2818),.q3(n147_5));
  bfr _b_2335(.a(_w_3151),.q(_w_3152));
  bfr _b_1569(.a(_w_2385),.q(_w_2386));
  bfr _b_1570(.a(_w_2386),.q(_w_2387));
  bfr _b_2397(.a(_w_3213),.q(_w_3214));
  spl2 g97_s_0(.a(n97),.q0(n97_0),.q1(n97_1));
  bfr _b_1719(.a(_w_2535),.q(_w_2536));
  bfr _b_2373(.a(_w_3189),.q(_w_3190));
  bfr _b_1572(.a(_w_2388),.q(_w_2389));
  bfr _b_1945(.a(_w_2761),.q(_w_2762));
  bfr _b_1573(.a(_w_2389),.q(_w_2390));
  spl3L g254_s_0(.a(n254),.q0(n254_0),.q1(n254_1),.q2(_w_2727));
  bfr _b_2182(.a(_w_2998),.q(n667));
  bfr _b_1574(.a(_w_2390),.q(_w_2391));
  bfr _b_2230(.a(_w_3046),.q(_w_3047));
  bfr _b_1577(.a(_w_2393),.q(_w_2394));
  bfr _b_1578(.a(_w_2394),.q(_w_2395));
  bfr _b_1580(.a(_w_2396),.q(_w_2397));
  bfr _b_1586(.a(_w_2402),.q(_w_2403));
  bfr _b_1588(.a(_w_2404),.q(_w_2405));
  bfr _b_1590(.a(_w_2406),.q(_w_2407));
  bfr _b_1591(.a(_w_2407),.q(_w_2408));
  bfr _b_1594(.a(_w_2410),.q(_w_2411));
  bfr _b_2190(.a(_w_3006),.q(_w_3007));
  and_bi g217(.a(n216_0),.b(G9_15),.q(n217));
  bfr _b_1597(.a(_w_2413),.q(n533_6));
  bfr _b_1598(.a(_w_2414),.q(_w_2415));
  bfr _b_1806(.a(_w_2622),.q(G30_4));
  bfr _b_2221(.a(_w_3037),.q(_w_3038));
  bfr _b_1599(.a(_w_2415),.q(_w_2416));
  bfr _b_1608(.a(_w_2424),.q(n401_10));
  bfr _b_1609(.a(_w_2425),.q(_w_2426));
  or_bb g599(.a(n585),.b(n598),.q(n599));
  bfr _b_1610(.a(_w_2426),.q(_w_2427));
  bfr _b_1611(.a(_w_2427),.q(_w_2428));
  spl2 g398_s_4(.a(n398_14),.q0(n398_16),.q1(n398_17));
  bfr _b_1612(.a(_w_2428),.q(_w_2429));
  bfr _b_1614(.a(_w_2430),.q(G14_14));
  bfr _b_2155(.a(_w_2971),.q(_w_2972));
  bfr _b_1615(.a(_w_2431),.q(_w_2432));
  bfr _b_1616(.a(_w_2432),.q(n675));
  bfr _b_1618(.a(_w_2434),.q(_w_2435));
  bfr _b_1619(.a(_w_2435),.q(n500_1));
  bfr _b_1620(.a(_w_2436),.q(n485));
  and_bi g209(.a(n208),.b(n147_3),.q(_w_2506));
  bfr _b_2208(.a(_w_3024),.q(_w_3025));
  bfr _b_2479(.a(_w_3295),.q(_w_3296));
  bfr _b_1624(.a(_w_2440),.q(n317_1));
  bfr _b_1625(.a(_w_2441),.q(n563));
  bfr _b_1627(.a(_w_2443),.q(_w_2444));
  bfr _b_1637(.a(_w_2453),.q(_w_2454));
  bfr _b_1629(.a(_w_2445),.q(_w_2446));
  bfr _b_1630(.a(_w_2446),.q(_w_2447));
  spl2 G17_s_0(.a(_w_3421),.q0(G17_0),.q1(_w_3222));
  bfr _b_1631(.a(_w_2447),.q(_w_2448));
  bfr _b_1632(.a(_w_2448),.q(_w_2449));
  bfr _b_1634(.a(_w_2450),.q(n149_3));
  bfr _b_1439(.a(_w_2255),.q(_w_2256));
  bfr _b_1900(.a(_w_2716),.q(_w_2717));
  bfr _b_1729(.a(_w_2545),.q(_w_2546));
  bfr _b_1638(.a(_w_2454),.q(_w_2455));
  or_bb g743(.a(_w_3412),.b(G19_0),.q(_w_3079));
  bfr _b_1645(.a(_w_2461),.q(_w_2462));
  bfr _b_1646(.a(_w_2462),.q(_w_2463));
  bfr _b_1379(.a(_w_2195),.q(n340_3));
  bfr _b_1648(.a(_w_2464),.q(_w_2465));
  bfr _b_1649(.a(_w_2465),.q(_w_2466));
  bfr _b_1651(.a(_w_2467),.q(_w_2468));
  bfr _b_2302(.a(_w_3118),.q(_w_3119));
  bfr _b_1654(.a(_w_2470),.q(_w_2471));
  bfr _b_1656(.a(_w_2472),.q(_w_2473));
  bfr _b_1938(.a(_w_2754),.q(_w_2755));
  or_bb g159(.a(n149_0),.b(n158),.q(n159));
  bfr _b_1657(.a(_w_2473),.q(_w_2474));
  bfr _b_1658(.a(_w_2474),.q(_w_2475));
  bfr _b_1661(.a(_w_2477),.q(_w_2478));
  and_bi g436(.a(n434),.b(n435),.q(n436));
  bfr _b_1664(.a(_w_2480),.q(_w_2481));
  bfr _b_1665(.a(_w_2481),.q(_w_2482));
  bfr _b_1667(.a(_w_2483),.q(_w_2484));
  and_bi g687(.a(n686),.b(n684_0),.q(n687));
  bfr _b_2062(.a(_w_2878),.q(_w_2879));
  bfr _b_1668(.a(_w_2484),.q(_w_2485));
  bfr _b_1672(.a(_w_2488),.q(_w_2489));
  bfr _b_1840(.a(_w_2656),.q(_w_2657));
  bfr _b_1675(.a(_w_2491),.q(_w_2492));
  bfr _b_2262(.a(_w_3078),.q(n201_3));
  bfr _b_1764(.a(_w_2580),.q(_w_2581));
  and_bi g555(.a(n374_9),.b(n554_0),.q(n555));
  bfr _b_1677(.a(_w_2493),.q(_w_2494));
  bfr _b_1680(.a(_w_2496),.q(_w_2497));
  bfr _b_1681(.a(_w_2497),.q(_w_2498));
  or_bb g414(.a(G10_11),.b(n401_10),.q(n414));
  bfr _b_1685(.a(_w_2501),.q(G3520));
  bfr _b_1918(.a(_w_2734),.q(n358));
  bfr _b_2010(.a(_w_2826),.q(_w_2827));
  bfr _b_1687(.a(_w_2503),.q(n613));
  bfr _b_2336(.a(_w_3152),.q(_w_3153));
  bfr _b_1689(.a(_w_2505),.q(n154));
  bfr _b_1694(.a(_w_2510),.q(_w_2511));
  bfr _b_2637(.a(G25),.q(_w_3453));
  bfr _b_1501(.a(_w_2317),.q(_w_2318));
  bfr _b_1695(.a(_w_2511),.q(n374_9));
  bfr _b_2427(.a(_w_3243),.q(_w_3244));
  bfr _b_1696(.a(_w_2512),.q(_w_2513));
  and_bb g712(.a(n708),.b(n711),.q(n712));
  bfr _b_2053(.a(_w_2869),.q(_w_2870));
  bfr _b_2186(.a(_w_3002),.q(_w_3003));
  bfr _b_1697(.a(_w_2513),.q(_w_2514));
  bfr _b_1761(.a(_w_2577),.q(_w_2578));
  bfr _b_2595(.a(G14),.q(_w_3411));
  bfr _b_1699(.a(_w_2515),.q(_w_2516));
  bfr _b_2673(.a(_w_3489),.q(_w_3490));
  and_bi g724(.a(n723),.b(n653_1),.q(n724));
  bfr _b_1701(.a(_w_2517),.q(_w_2518));
  bfr _b_1702(.a(_w_2518),.q(n375));
  or_bb g173(.a(n170),.b(n172),.q(n173));
  bfr _b_1703(.a(_w_2519),.q(_w_2520));
  bfr _b_2732(.a(_w_3548),.q(_w_3549));
  spl2 G4_s_15(.a(G4_50),.q0(G4_51),.q1(G4_52));
  bfr _b_1704(.a(_w_2520),.q(_w_2521));
  bfr _b_1705(.a(_w_2521),.q(_w_2522));
  bfr _b_1711(.a(_w_2527),.q(n392_14));
  bfr _b_1712(.a(_w_2528),.q(_w_2529));
  bfr _b_1714(.a(_w_2530),.q(_w_2531));
  bfr _b_1406(.a(_w_2222),.q(_w_2223));
  bfr _b_2205(.a(_w_3021),.q(_w_3022));
  and_bi g642(.a(n604_2),.b(n372_6),.q(n642));
  bfr _b_2246(.a(_w_3062),.q(_w_3063));
  bfr _b_1716(.a(_w_2532),.q(_w_2533));
  bfr _b_1717(.a(_w_2533),.q(_w_2534));
  bfr _b_1698(.a(_w_2514),.q(_w_2515));
  bfr _b_1718(.a(_w_2534),.q(_w_2535));
  bfr _b_1720(.a(_w_2536),.q(_w_2537));
  bfr _b_1722(.a(_w_2538),.q(_w_2539));
  bfr _b_1510(.a(_w_2326),.q(_w_2327));
  bfr _b_1723(.a(_w_2539),.q(_w_2540));
  bfr _b_2467(.a(_w_3283),.q(n623_1));
  bfr _b_1725(.a(_w_2541),.q(_w_2542));
  spl2 g834_s_2(.a(n834_3),.q0(n834_4),.q1(n834_5));
  bfr _b_1726(.a(_w_2542),.q(_w_2543));
  bfr _b_1732(.a(_w_2548),.q(_w_2549));
  bfr _b_1735(.a(_w_2551),.q(_w_2552));
  spl2 G43_s_1(.a(G43_1),.q0(G43_2),.q1(G43_3));
  bfr _b_1740(.a(_w_2556),.q(_w_2557));
  bfr _b_1741(.a(_w_2557),.q(_w_2558));
  bfr _b_1839(.a(_w_2655),.q(_w_2656));
  bfr _b_1742(.a(_w_2558),.q(_w_2559));
  bfr _b_1747(.a(_w_2563),.q(_w_2564));
  bfr _b_1749(.a(_w_2565),.q(_w_2566));
  bfr _b_1751(.a(_w_2567),.q(n105_1));
  spl2 g147_s_3(.a(n147_9),.q0(n147_10),.q1(_w_3367));
  bfr _b_1752(.a(_w_2568),.q(n439));
  bfr _b_1757(.a(_w_2573),.q(_w_2574));
  bfr _b_1758(.a(_w_2574),.q(_w_2575));
  bfr _b_1988(.a(_w_2804),.q(n71));
  bfr _b_1763(.a(_w_2579),.q(_w_2580));
  bfr _b_1765(.a(_w_2581),.q(_w_2582));
  bfr _b_1606(.a(_w_2422),.q(n350));
  bfr _b_1766(.a(_w_2582),.q(_w_2583));
  bfr _b_1767(.a(_w_2583),.q(_w_2584));
  bfr _b_1774(.a(_w_2590),.q(_w_2591));
  bfr _b_1775(.a(_w_2591),.q(_w_2592));
  and_bi g57(.a(G32_0),.b(G9_0),.q(n57));
  bfr _b_1916(.a(_w_2732),.q(_w_2733));
  spl2 G26_s_1(.a(G26_1),.q0(G26_2),.q1(G26_3));
  bfr _b_2326(.a(_w_3142),.q(_w_3143));
  bfr _b_2375(.a(_w_3191),.q(n240_3));
  bfr _b_1776(.a(_w_2592),.q(_w_2593));
  bfr _b_1778(.a(_w_2594),.q(_w_2595));
  bfr _b_1728(.a(_w_2544),.q(_w_2545));
  bfr _b_1781(.a(_w_2597),.q(n210_1));
  spl2 g587_s_0(.a(n587),.q0(n587_0),.q1(n587_1));
  bfr _b_1783(.a(_w_2599),.q(_w_2600));
  bfr _b_1786(.a(_w_2602),.q(_w_2603));
  bfr _b_1788(.a(_w_2604),.q(_w_2605));
  bfr _b_1989(.a(_w_2805),.q(_w_2806));
  bfr _b_1367(.a(_w_2183),.q(_w_2184));
  spl4L g398_s_2(.a(n398_6),.q0(n398_8),.q1(n398_9),.q2(n398_10),.q3(n398_11));
  bfr _b_2174(.a(_w_2990),.q(_w_2991));
  or_bb g394(.a(G26_3),.b(n383_1),.q(n394));
  bfr _b_1789(.a(_w_2605),.q(_w_2606));
  and_bi g620(.a(n395_17),.b(G7_17),.q(n620));
  spl2 g436_s_1(.a(n436_1),.q0(n436_2),.q1(_w_2133));
  bfr _b_1790(.a(_w_2606),.q(G3536));
  bfr _b_1794(.a(_w_2610),.q(G13_21));
  bfr _b_2125(.a(_w_2941),.q(_w_2942));
  bfr _b_2570(.a(_w_3386),.q(_w_3387));
  bfr _b_1796(.a(_w_2612),.q(n426));
  bfr _b_1791(.a(_w_2607),.q(_w_2608));
  bfr _b_1798(.a(_w_2614),.q(n369));
  bfr _b_1803(.a(_w_2619),.q(_w_2620));
  spl2 g130_s_1(.a(n130_2),.q0(n130_3),.q1(n130_4));
  bfr _b_2197(.a(_w_3013),.q(_w_3014));
  bfr _b_1746(.a(_w_2562),.q(_w_2563));
  bfr _b_1804(.a(_w_2620),.q(n317_3));
  bfr _b_1805(.a(_w_2621),.q(G50_1));
  bfr _b_1884(.a(_w_2700),.q(_w_2701));
  bfr _b_2323(.a(_w_3139),.q(n688_1));
  bfr _b_2578(.a(_w_3394),.q(G9_8));
  bfr _b_1807(.a(_w_2623),.q(G30_6));
  spl2 g227_s_0(.a(n227),.q0(n227_0),.q1(_w_3392));
  and_bi g75(.a(n51_4),.b(G7_15),.q(n75));
  bfr _b_1976(.a(_w_2792),.q(_w_2793));
  bfr _b_1808(.a(_w_2624),.q(_w_2625));
  bfr _b_2621(.a(_w_3437),.q(_w_3432));
  or_bb g444(.a(G7_19),.b(n407_12),.q(n444));
  bfr _b_1813(.a(_w_2629),.q(n143_1));
  and_bi g60(.a(G36_0),.b(G13_0),.q(n60));
  bfr _b_1814(.a(_w_2630),.q(_w_2631));
  and_bi g633(.a(n629_0),.b(n632),.q(n633));
  or_bb g399(.a(G41_0),.b(_w_3493),.q(_w_2519));
  bfr _b_1819(.a(_w_2635),.q(n303));
  bfr _b_1820(.a(_w_2636),.q(_w_2637));
  bfr _b_1821(.a(_w_2637),.q(_w_2638));
  bfr _b_1822(.a(_w_2638),.q(_w_2639));
  bfr _b_1332(.a(_w_2148),.q(_w_2149));
  bfr _b_1824(.a(_w_2640),.q(n79));
  or_bb g538(.a(n428_2),.b(n537_0),.q(n538));
  bfr _b_1391(.a(_w_2207),.q(n306_3));
  bfr _b_1827(.a(_w_2643),.q(_w_2644));
  bfr _b_1829(.a(_w_2645),.q(n344_1));
  bfr _b_1832(.a(_w_2648),.q(_w_2649));
  bfr _b_1853(.a(_w_2669),.q(_w_2670));
  bfr _b_1833(.a(_w_2649),.q(_w_2650));
  bfr _b_2676(.a(_w_3492),.q(_w_3487));
  bfr _b_1319(.a(_w_2135),.q(n436_1));
  bfr _b_1835(.a(_w_2651),.q(_w_2652));
  bfr _b_2432(.a(_w_3248),.q(_w_3249));
  bfr _b_1836(.a(_w_2652),.q(_w_2653));
  spl4L g392_s_0(.a(n392),.q0(n392_0),.q1(n392_1),.q2(n392_2),.q3(n392_3));
  bfr _b_2227(.a(_w_3043),.q(_w_3044));
  bfr _b_1842(.a(_w_2658),.q(G5_4));
  bfr _b_1844(.a(_w_2660),.q(_w_2661));
  bfr _b_2332(.a(_w_3148),.q(n495_1));
  spl3L g540_s_0(.a(n540),.q0(n540_0),.q1(n540_1),.q2(_w_3150));
  bfr _b_1846(.a(_w_2662),.q(_w_2663));
  bfr _b_1847(.a(_w_2663),.q(_w_2664));
  bfr _b_1850(.a(_w_2666),.q(_w_2667));
  bfr _b_2048(.a(_w_2864),.q(G3524));
  bfr _b_2338(.a(_w_3154),.q(_w_3155));
  and_bi g578(.a(G10_5),.b(G22_5),.q(n578));
  bfr _b_1852(.a(_w_2668),.q(_w_2669));
  bfr _b_2404(.a(_w_3220),.q(G44_2));
  bfr _b_1854(.a(_w_2670),.q(_w_2671));
  bfr _b_1858(.a(_w_2674),.q(_w_2675));
  bfr _b_2056(.a(_w_2872),.q(_w_2873));
  bfr _b_1861(.a(_w_2677),.q(_w_2678));
  bfr _b_1862(.a(_w_2678),.q(_w_2679));
  bfr _b_2677(.a(G45),.q(_w_3493));
  bfr _b_1866(.a(_w_2682),.q(_w_2683));
  bfr _b_1868(.a(_w_2684),.q(_w_2685));
  bfr _b_1869(.a(_w_2685),.q(_w_2686));
  bfr _b_1872(.a(_w_2688),.q(_w_2689));
  bfr _b_2195(.a(_w_3011),.q(_w_3012));
  bfr _b_1876(.a(_w_2692),.q(_w_2693));
  bfr _b_1878(.a(_w_2694),.q(_w_2695));
  bfr _b_1885(.a(_w_2701),.q(_w_2702));
  bfr _b_1887(.a(_w_2703),.q(G3522));
  bfr _b_1891(.a(_w_2707),.q(_w_2708));
  bfr _b_1893(.a(_w_2709),.q(_w_2710));
  or_bb g624(.a(G9_16),.b(n401_17),.q(n624));
  bfr _b_1895(.a(_w_2711),.q(_w_2712));
  bfr _b_1898(.a(_w_2714),.q(_w_2715));
  spl2 g697_s_0(.a(n697),.q0(n697_0),.q1(n697_1));
  bfr _b_1901(.a(_w_2717),.q(_w_2718));
  bfr _b_1412(.a(_w_2228),.q(_w_2229));
  bfr _b_1902(.a(_w_2718),.q(_w_2719));
  and_bi g621(.a(G22_9),.b(n398_18),.q(n621));
  bfr _b_1903(.a(_w_2719),.q(_w_2720));
  bfr _b_1302(.a(_w_2118),.q(_w_2119));
  bfr _b_1904(.a(_w_2720),.q(_w_2721));
  bfr _b_1969(.a(_w_2785),.q(_w_2786));
  bfr _b_1831(.a(_w_2647),.q(_w_2648));
  bfr _b_1907(.a(_w_2723),.q(_w_2724));
  bfr _b_2279(.a(_w_3095),.q(_w_3096));
  bfr _b_1910(.a(_w_2726),.q(G11_3));
  and_bi g118(.a(n116_1),.b(n113_1),.q(n118));
  bfr _b_1912(.a(_w_2728),.q(n254_2));
  spl2 G14_s_3(.a(G14_5),.q0(G14_6),.q1(G14_7));
  bfr _b_2225(.a(_w_3041),.q(_w_3042));
  bfr _b_1913(.a(_w_2729),.q(_w_2730));
  bfr _b_1925(.a(_w_2741),.q(_w_2742));
  bfr _b_1926(.a(_w_2742),.q(n386_1));
  bfr _b_1515(.a(_w_2331),.q(_w_2332));
  bfr _b_1923(.a(_w_2739),.q(n638));
  bfr _b_1927(.a(_w_2743),.q(G14_5));
  bfr _b_1929(.a(_w_2745),.q(n226));
  bfr _b_2431(.a(_w_3247),.q(_w_3248));
  bfr _b_1930(.a(_w_2746),.q(_w_2747));
  and_bi g400(.a(n399_0),.b(n398_1),.q(n400));
  bfr _b_1931(.a(_w_2747),.q(_w_2748));
  bfr _b_1933(.a(_w_2749),.q(n395_14));
  bfr _b_1936(.a(_w_2752),.q(_w_2753));
  bfr _b_1939(.a(_w_2755),.q(_w_2756));
  bfr _b_1940(.a(_w_2756),.q(_w_2757));
  and_bb g479(.a(n344_0),.b(n361_17),.q(n479));
  bfr _b_1941(.a(_w_2757),.q(_w_2758));
  bfr _b_1942(.a(_w_2758),.q(_w_2759));
  bfr _b_1946(.a(_w_2762),.q(_w_2763));
  bfr _b_1948(.a(_w_2764),.q(_w_2765));
  bfr _b_1949(.a(_w_2765),.q(_w_2766));
  bfr _b_1950(.a(_w_2766),.q(_w_2767));
  spl2 g314_s_0(.a(n314),.q0(n314_0),.q1(n314_1));
  bfr _b_1684(.a(_w_2500),.q(_w_2501));
  bfr _b_1951(.a(_w_2767),.q(_w_2768));
  bfr _b_1957(.a(_w_2773),.q(_w_2774));
  bfr _b_1958(.a(_w_2774),.q(_w_2775));
  or_bb g69(.a(n67),.b(n68),.q(n69));
  bfr _b_1896(.a(_w_2712),.q(_w_2713));
  bfr _b_2102(.a(_w_2918),.q(_w_2919));
  spl2 g553_s_0(.a(n553),.q0(n553_0),.q1(n553_1));
  bfr _b_1482(.a(_w_2298),.q(_w_2299));
  bfr _b_1959(.a(_w_2775),.q(_w_2776));
  bfr _b_1961(.a(_w_2777),.q(_w_2778));
  bfr _b_1500(.a(_w_2316),.q(_w_2317));
  bfr _b_1965(.a(_w_2781),.q(_w_2782));
  bfr _b_1966(.a(_w_2782),.q(_w_2783));
  bfr _b_1967(.a(_w_2783),.q(_w_2784));
  bfr _b_2707(.a(_w_3523),.q(_w_3515));
  bfr _b_1968(.a(_w_2784),.q(_w_2785));
  bfr _b_1300(.a(_w_2116),.q(_w_2117));
  bfr _b_1970(.a(_w_2786),.q(_w_2787));
  bfr _b_1971(.a(_w_2787),.q(_w_2788));
  bfr _b_1972(.a(_w_2788),.q(_w_2789));
  bfr _b_1727(.a(_w_2543),.q(_w_2544));
  bfr _b_1974(.a(_w_2790),.q(_w_2791));
  bfr _b_1975(.a(_w_2791),.q(_w_2792));
  bfr _b_2035(.a(_w_2851),.q(_w_2852));
  bfr _b_2224(.a(_w_3040),.q(_w_3041));
  bfr _b_1977(.a(_w_2793),.q(_w_2794));
  bfr _b_1979(.a(_w_2795),.q(_w_2796));
  bfr _b_1981(.a(_w_2797),.q(_w_2798));
  bfr _b_1982(.a(_w_2798),.q(_w_2799));
  bfr _b_1983(.a(_w_2799),.q(_w_2800));
  bfr _b_1984(.a(_w_2800),.q(G3521));
  bfr _b_1640(.a(_w_2456),.q(_w_2457));
  bfr _b_1985(.a(_w_2801),.q(_w_2802));
  bfr _b_1986(.a(_w_2802),.q(_w_2803));
  or_bb g405(.a(n397),.b(n404),.q(n405));
  bfr _b_1799(.a(_w_2615),.q(_w_2616));
  bfr _b_1991(.a(_w_2807),.q(_w_2808));
  bfr _b_1993(.a(_w_2809),.q(_w_2810));
  bfr _b_1994(.a(_w_2810),.q(_w_2811));
  bfr _b_2058(.a(_w_2874),.q(_w_2875));
  bfr _b_1992(.a(_w_2808),.q(_w_2809));
  bfr _b_1995(.a(_w_2811),.q(_w_2812));
  bfr _b_1996(.a(_w_2812),.q(_w_2813));
  bfr _b_2199(.a(_w_3015),.q(_w_3016));
  bfr _b_1997(.a(_w_2813),.q(_w_2814));
  spl2 g812_s_0(.a(n812),.q0(n812_0),.q1(_w_2893));
  bfr _b_1509(.a(_w_2325),.q(_w_2326));
  bfr _b_1998(.a(_w_2814),.q(_w_2815));
  bfr _b_2455(.a(_w_3271),.q(_w_3272));
  bfr _b_2000(.a(_w_2816),.q(n147_2));
  spl2 g240_s_0(.a(n240),.q0(n240_0),.q1(_w_3187));
  or_bb g461(.a(n401_19),.b(n460_1),.q(n461));
  bfr _b_2001(.a(_w_2817),.q(n147_3));
  bfr _b_2002(.a(_w_2818),.q(n147_4));
  bfr _b_2003(.a(_w_2819),.q(n210));
  bfr _b_2004(.a(_w_2820),.q(n653_1));
  bfr _b_2005(.a(_w_2821),.q(_w_2822));
  bfr _b_2622(.a(G21),.q(_w_3439));
  bfr _b_2007(.a(_w_2823),.q(_w_2824));
  bfr _b_2601(.a(_w_3417),.q(_w_3418));
  bfr _b_2011(.a(_w_2827),.q(_w_2828));
  bfr _b_2012(.a(_w_2828),.q(_w_2829));
  bfr _b_2014(.a(_w_2830),.q(_w_2831));
  bfr _b_2016(.a(_w_2832),.q(_w_2833));
  bfr _b_2027(.a(_w_2843),.q(_w_2844));
  spl3L g696_s_0(.a(n696),.q0(n696_0),.q1(n696_1),.q2(n696_2));
  bfr _b_2017(.a(_w_2833),.q(_w_2834));
  bfr _b_1363(.a(_w_2179),.q(_w_2180));
  bfr _b_2018(.a(_w_2834),.q(_w_2835));
  bfr _b_1908(.a(_w_2724),.q(n729));
  bfr _b_2019(.a(_w_2835),.q(_w_2836));
  bfr _b_2709(.a(G50),.q(_w_3526));
  bfr _b_2024(.a(_w_2840),.q(G4_37));
  bfr _b_2025(.a(_w_2841),.q(_w_2842));
  bfr _b_2026(.a(_w_2842),.q(_w_2843));
  bfr _b_2029(.a(_w_2845),.q(_w_2846));
  bfr _b_2072(.a(_w_2888),.q(_w_2889));
  bfr _b_2030(.a(_w_2846),.q(_w_2847));
  bfr _b_2034(.a(_w_2850),.q(_w_2851));
  spl3L g224_s_0(.a(n224),.q0(n224_0),.q1(n224_1),.q2(_w_3200));
  bfr _b_2036(.a(_w_2852),.q(_w_2853));
  bfr _b_2037(.a(_w_2853),.q(_w_2854));
  or_bb g656(.a(n654_0),.b(n655),.q(n656));
  bfr _b_1531(.a(_w_2347),.q(_w_2348));
  bfr _b_1593(.a(_w_2409),.q(_w_2410));
  bfr _b_2039(.a(_w_2855),.q(_w_2856));
  bfr _b_2040(.a(_w_2856),.q(_w_2857));
  bfr _b_1434(.a(_w_2250),.q(_w_2251));
  bfr _b_2041(.a(_w_2857),.q(_w_2858));
  bfr _b_2042(.a(_w_2858),.q(_w_2859));
  bfr _b_1688(.a(_w_2504),.q(n151_2));
  bfr _b_2043(.a(_w_2859),.q(_w_2860));
  bfr _b_2044(.a(_w_2860),.q(_w_2861));
  bfr _b_2047(.a(_w_2863),.q(_w_2864));
  bfr _b_1603(.a(_w_2419),.q(_w_2420));
  bfr _b_2049(.a(_w_2865),.q(_w_2866));
  bfr _b_2050(.a(_w_2866),.q(_w_2867));
  bfr _b_2055(.a(_w_2871),.q(_w_2872));
  or_bb g527(.a(n521_0),.b(n526),.q(n527));
  bfr _b_2057(.a(_w_2873),.q(_w_2874));
  bfr _b_2059(.a(_w_2875),.q(_w_2876));
  bfr _b_2723(.a(_w_3539),.q(_w_3540));
  bfr _b_2061(.a(_w_2877),.q(_w_2878));
  bfr _b_2472(.a(_w_3288),.q(n126_3));
  spl3L G44_s_0(.a(_w_3487),.q0(G44_0),.q1(G44_1),.q2(_w_3219));
  bfr _b_2141(.a(_w_2957),.q(_w_2958));
  bfr _b_2064(.a(_w_2880),.q(_w_2881));
  bfr _b_2065(.a(_w_2881),.q(_w_2882));
  spl4L g379_s_2(.a(n379_3),.q0(n379_7),.q1(n379_8),.q2(n379_9),.q3(_w_2368));
  bfr _b_2067(.a(_w_2883),.q(_w_2884));
  bfr _b_2071(.a(_w_2887),.q(_w_2888));
  bfr _b_2074(.a(_w_2890),.q(_w_2891));
  bfr _b_2075(.a(_w_2891),.q(_w_2892));
  bfr _b_2243(.a(_w_3059),.q(_w_3060));
  spl2 G12_s_0(.a(_w_3409),.q0(G12_0),.q1(_w_3168));
  bfr _b_2079(.a(_w_2895),.q(n748));
  bfr _b_2259(.a(_w_3075),.q(_w_3076));
  bfr _b_2080(.a(_w_2896),.q(_w_2897));
  or_bb g94(.a(n92),.b(n93),.q(n94));
  bfr _b_2082(.a(_w_2898),.q(_w_2899));
  bfr _b_1408(.a(_w_2224),.q(G7_1));
  bfr _b_2083(.a(_w_2899),.q(_w_2900));
  bfr _b_2085(.a(_w_2901),.q(_w_2902));
  bfr _b_2474(.a(_w_3290),.q(_w_3291));
  bfr _b_2088(.a(_w_2904),.q(_w_2905));
  bfr _b_2089(.a(_w_2905),.q(_w_2906));
  bfr _b_2091(.a(_w_2907),.q(n73_1));
  bfr _b_1461(.a(_w_2277),.q(_w_2278));
  bfr _b_2093(.a(_w_2909),.q(_w_2910));
  and_bb g192(.a(G3_14),.b(n129_1),.q(n192));
  bfr _b_1920(.a(_w_2736),.q(_w_2737));
  bfr _b_2097(.a(_w_2913),.q(_w_2914));
  spl2 g148_s_0(.a(n148),.q0(n148_0),.q1(n148_1));
  bfr _b_2103(.a(_w_2919),.q(_w_2920));
  bfr _b_2099(.a(_w_2915),.q(_w_2916));
  bfr _b_2100(.a(_w_2916),.q(_w_2917));
  bfr _b_2101(.a(_w_2917),.q(_w_2918));
  or_bb g182(.a(n178),.b(n181),.q(n182));
  bfr _b_2105(.a(_w_2921),.q(_w_2922));
  bfr _b_2106(.a(_w_2922),.q(_w_2923));
  bfr _b_2107(.a(_w_2923),.q(_w_2924));
  bfr _b_2108(.a(_w_2924),.q(_w_2925));
  spl3L g284_s_0(.a(n284),.q0(n284_0),.q1(n284_1),.q2(n284_2));
  bfr _b_2136(.a(_w_2952),.q(_w_2953));
  bfr _b_2109(.a(_w_2925),.q(_w_2926));
  and_bi g111(.a(G13_18),.b(G11_15),.q(n111));
  bfr _b_2110(.a(_w_2926),.q(n530));
  bfr _b_2111(.a(_w_2927),.q(n179_1));
  bfr _b_2286(.a(_w_3102),.q(_w_3103));
  spl2 G7_s_2(.a(G7_4),.q0(G7_5),.q1(G7_6));
  bfr _b_2113(.a(_w_2929),.q(n765_1));
  bfr _b_2120(.a(_w_2936),.q(_w_2937));
  bfr _b_2545(.a(_w_3361),.q(_w_3362));
  bfr _b_2351(.a(_w_3167),.q(n343_2));
  and_bi g692(.a(n691),.b(n684_1),.q(n692));
  bfr _b_2121(.a(_w_2937),.q(_w_2938));
  bfr _b_2122(.a(_w_2938),.q(_w_2939));
  bfr _b_2417(.a(_w_3233),.q(_w_3234));
  bfr _b_2126(.a(_w_2942),.q(G42_5));
  bfr _b_2343(.a(_w_3159),.q(n171_1));
  bfr _b_2128(.a(_w_2944),.q(G38_1));
  bfr _b_2131(.a(_w_2947),.q(_w_2948));
  bfr _b_2133(.a(_w_2949),.q(_w_2950));
  bfr _b_2134(.a(_w_2950),.q(_w_2951));
  bfr _b_2138(.a(_w_2954),.q(_w_2955));
  bfr _b_2139(.a(_w_2955),.q(_w_2956));
  bfr _b_2140(.a(_w_2956),.q(_w_2957));
  bfr _b_1770(.a(_w_2586),.q(G3532));
  bfr _b_2144(.a(_w_2960),.q(_w_2961));
  bfr _b_2145(.a(_w_2961),.q(_w_2962));
  and_bb g221(.a(n129_8),.b(n220),.q(n221));
  bfr _b_2285(.a(_w_3101),.q(_w_3102));
  bfr _b_2147(.a(_w_2963),.q(_w_2964));
  bfr _b_2214(.a(_w_3030),.q(_w_3031));
  bfr _b_2148(.a(_w_2964),.q(_w_2965));
  bfr _b_2149(.a(_w_2965),.q(_w_2966));
  bfr _b_2150(.a(_w_2966),.q(_w_2967));
  spl2 g432_s_1(.a(G3528_2),.q0(G3528_3),.q1(_w_3348));
  and_bi g327(.a(n277_2),.b(n326),.q(n327));
  bfr _b_2151(.a(_w_2967),.q(_w_2968));
  bfr _b_2481(.a(_w_3297),.q(_w_3298));
  bfr _b_2156(.a(_w_2972),.q(_w_2973));
  bfr _b_2158(.a(_w_2974),.q(_w_2975));
  bfr _b_2162(.a(_w_2978),.q(n619));
  bfr _b_2163(.a(_w_2979),.q(_w_2980));
  spl3L g130_s_0(.a(n130),.q0(n130_0),.q1(n130_1),.q2(n130_2));
  bfr _b_2164(.a(_w_2980),.q(_w_2981));
  bfr _b_2400(.a(_w_3216),.q(_w_3217));
  bfr _b_2166(.a(_w_2982),.q(n805));
  bfr _b_2261(.a(_w_3077),.q(n719));
  bfr _b_2295(.a(_w_3111),.q(_w_3112));
  bfr _b_2169(.a(_w_2985),.q(_w_2986));
  bfr _b_2171(.a(_w_2987),.q(_w_2988));
  bfr _b_1692(.a(_w_2508),.q(n547));
  bfr _b_2313(.a(_w_3129),.q(_w_3130));
  bfr _b_2172(.a(_w_2988),.q(_w_2989));
  bfr _b_2319(.a(_w_3135),.q(_w_3136));
  bfr _b_2173(.a(_w_2989),.q(_w_2990));
  bfr _b_2176(.a(_w_2992),.q(n639));
  bfr _b_1812(.a(_w_2628),.q(_w_2629));
  bfr _b_2180(.a(_w_2996),.q(n643));
  bfr _b_2189(.a(_w_3005),.q(_w_3006));
  bfr _b_2191(.a(_w_3007),.q(_w_3008));
  bfr _b_2192(.a(_w_3008),.q(_w_3009));
  bfr _b_2612(.a(_w_3428),.q(_w_3429));
  and_bb g491(.a(n224_2),.b(n361_6),.q(n491));
  bfr _b_2196(.a(_w_3012),.q(_w_3013));
  bfr _b_2303(.a(_w_3119),.q(_w_3120));
  bfr _b_2200(.a(_w_3016),.q(_w_3017));
  and_bi g446(.a(G9_10),.b(G21_5),.q(n446));
  bfr _b_2201(.a(_w_3017),.q(_w_3018));
  bfr _b_2202(.a(_w_3018),.q(_w_3019));
  and_bi g802(.a(n629_2),.b(n801),.q(n802));
  bfr _b_2211(.a(_w_3027),.q(_w_3028));
  bfr _b_2216(.a(_w_3032),.q(_w_3033));
  bfr _b_2217(.a(_w_3033),.q(_w_3034));
  bfr _b_2220(.a(_w_3036),.q(_w_3037));
  and_bi g236(.a(n162_9),.b(n233_1),.q(n236));
  bfr _b_2258(.a(_w_3074),.q(_w_3075));
  bfr _b_2222(.a(_w_3038),.q(_w_3039));
  bfr _b_2226(.a(_w_3042),.q(_w_3043));
  bfr _b_2229(.a(_w_3045),.q(_w_3046));
  bfr _b_2231(.a(_w_3047),.q(_w_3048));
  bfr _b_2235(.a(_w_3051),.q(_w_3052));
  bfr _b_2236(.a(_w_3052),.q(_w_3053));
  bfr _b_2237(.a(_w_3053),.q(_w_3054));
  bfr _b_2245(.a(_w_3061),.q(_w_3062));
  bfr _b_2248(.a(_w_3064),.q(n563_1));
  bfr _b_2249(.a(_w_3065),.q(_w_3066));
  bfr _b_2250(.a(_w_3066),.q(n689));
  bfr _b_2260(.a(_w_3076),.q(G3532_0));
  bfr _b_2264(.a(_w_3080),.q(_w_3081));
  bfr _b_2265(.a(_w_3081),.q(_w_3082));
  bfr _b_2266(.a(_w_3082),.q(_w_3083));
  bfr _b_2268(.a(_w_3084),.q(_w_3085));
  bfr _b_2269(.a(_w_3085),.q(n818));
  bfr _b_2270(.a(_w_3086),.q(_w_3087));
  bfr _b_1568(.a(_w_2384),.q(n727));
  bfr _b_2273(.a(_w_3089),.q(_w_3090));
  bfr _b_2275(.a(_w_3091),.q(_w_3092));
  spl2 G27_s_0(.a(_w_3455),.q0(G27_0),.q1(_w_3257));
  bfr _b_2277(.a(_w_3093),.q(_w_3094));
  bfr _b_2280(.a(_w_3096),.q(_w_3097));
  bfr _b_2052(.a(_w_2868),.q(_w_2869));
  and_bi g229(.a(n227_0),.b(n228),.q(n229));
  bfr _b_2281(.a(_w_3097),.q(_w_3098));
  bfr _b_2272(.a(_w_3088),.q(_w_3089));
  bfr _b_2282(.a(_w_3098),.q(_w_3099));
  bfr _b_1563(.a(_w_2379),.q(n377));
  bfr _b_2288(.a(_w_3104),.q(_w_3105));
  bfr _b_2290(.a(_w_3106),.q(G11_7));
  bfr _b_2292(.a(_w_3108),.q(_w_3109));
  bfr _b_2298(.a(_w_3114),.q(G14_3));
  bfr _b_2299(.a(_w_3115),.q(_w_3116));
  bfr _b_1600(.a(_w_2416),.q(n357));
  bfr _b_2304(.a(_w_3120),.q(_w_3121));
  bfr _b_2308(.a(_w_3124),.q(_w_3125));
  bfr _b_2310(.a(_w_3126),.q(_w_3127));
  and_bi g301(.a(G13_12),.b(n250_2),.q(n301));
  bfr _b_2311(.a(_w_3127),.q(n807));
  bfr _b_2312(.a(_w_3128),.q(_w_3129));
  bfr _b_2341(.a(_w_3157),.q(_w_3158));
  bfr _b_2314(.a(_w_3130),.q(_w_3131));
  bfr _b_2317(.a(_w_3133),.q(G39_4));
  bfr _b_2318(.a(_w_3134),.q(_w_3135));
  bfr _b_2638(.a(G26),.q(_w_3454));
  and_bi g332(.a(G41_2),.b(G4_19),.q(n332));
  bfr _b_2322(.a(_w_3138),.q(_w_3139));
  bfr _b_2213(.a(_w_3029),.q(_w_3030));
  bfr _b_2324(.a(_w_3140),.q(_w_3141));
  bfr _b_2325(.a(_w_3141),.q(_w_3142));
  bfr _b_2330(.a(_w_3146),.q(n735_1));
  and_bb g659(.a(n650),.b(n658),.q(n659));
  bfr _b_2331(.a(_w_3147),.q(_w_3148));
  bfr _b_2334(.a(_w_3150),.q(n540_2));
  or_bb g142(.a(n132),.b(n141),.q(n142));
  bfr _b_2339(.a(_w_3155),.q(_w_3156));
  spl2 G41_s_1(.a(G41_1),.q0(G41_2),.q1(_w_3284));
  bfr _b_2340(.a(_w_3156),.q(G47_2));
  bfr _b_2348(.a(_w_3164),.q(_w_3165));
  spl2 g537_s_0(.a(n537),.q0(n537_0),.q1(n537_1));
  bfr _b_1471(.a(_w_2287),.q(_w_2288));
  bfr _b_2352(.a(_w_3168),.q(G12_1));
  bfr _b_2146(.a(_w_2962),.q(_w_2963));
  bfr _b_2353(.a(_w_3169),.q(G4_8));
  bfr _b_2581(.a(_w_3397),.q(_w_3398));
  bfr _b_2355(.a(_w_3171),.q(n806));
endmodule
