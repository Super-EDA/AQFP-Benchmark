module counter_64 (in_15_,in_0_,in_4_,in_29_,in_38_,in_53_,in_42_,in_11_,in_59_,in_48_,in_54_,in_16_,in_43_,in_37_,in_61_,in_14_,in_62_,in_60_,in_40_,in_5_,in_28_,in_7_,in_6_,in_34_,in_57_,in_3_,in_56_,in_45_,in_10_,in_27_,in_21_,in_25_,in_22_,in_12_,in_58_,in_36_,in_51_,in_18_,in_9_,in_39_,in_24_,in_26_,in_8_,in_41_,in_55_,in_2_,in_49_,in_19_,in_35_,in_50_,in_32_,in_30_,in_33_,in_17_,in_31_,in_44_,in_1_,in_23_,in_52_,in_20_,in_46_,in_13_,in_63_,in_47_,out_1_,out_3_,out_6_,out_2_,out_0_,out_4_,out_5_);
  input in_15_,in_0_,in_4_,in_29_,in_38_,in_53_,in_42_,in_11_,in_59_,in_48_,in_54_,in_16_,in_43_,in_37_,in_61_,in_14_,in_62_,in_60_,in_40_,in_5_,in_28_,in_7_,in_6_,in_34_,in_57_,in_3_,in_56_,in_45_,in_10_,in_27_,in_21_,in_25_,in_22_,in_12_,in_58_,in_36_,in_51_,in_18_,in_9_,in_39_,in_24_,in_26_,in_8_,in_41_,in_55_,in_2_,in_49_,in_19_,in_35_,in_50_,in_32_,in_30_,in_33_,in_17_,in_31_,in_44_,in_1_,in_23_,in_52_,in_20_,in_46_,in_13_,in_63_,in_47_;
  output out_1_,out_3_,out_6_,out_2_,out_0_,out_4_,out_5_;
  wire _w_804,_w_800,_w_796,_w_794,_w_788,_w_786,_w_783,_w_781,_w_780,_w_778,_w_777,_w_776,_w_775,_w_774,_w_771,_w_770,_w_769,_w_768,_w_766,_w_765,_w_762,_w_758,_w_757,_w_756,_w_755,_w_767,_w_753,_w_748,_w_747,_w_745,_w_744,_w_739,_w_735,_w_734,_w_772,_w_733,_w_732,_w_731,_w_729,_w_728,_w_727,_w_723,_w_721,_w_716,_w_714,_w_713,_w_712,_w_710,_w_708,_w_707,_w_706,_w_705,_w_704,_w_702,_w_699,_w_698,_w_694,_w_693,_w_692,_w_691,_w_696,_w_689,_w_688,_w_685,_w_750,_w_684,_w_680,_w_784,_w_677,_w_672,_w_673,_w_671,_w_670,_w_669,_w_668,_w_666,_w_799,_w_665,_w_754,_w_664,_w_663,_w_662,_w_661,_w_667,_w_660,_w_686,_w_656,_w_655,_w_654,_w_650,_w_648,_w_647,_w_803,_w_646,_w_645,_w_751,_w_644,_w_643,_w_640,_w_637,_w_636,_w_635,_w_632,_w_631,_w_629,_w_634,_w_628,_w_627,_w_623,_w_618,_w_615,_w_614,_w_613,_w_612,_w_611,_w_608,_w_607,_w_606,_w_605,_w_601,_w_740,n238_2,n238_1,n238_0,n235_0,n232_1,n107_1,n107_0,_w_641,n239_1,n226_2,n225_1,n225_0,n219_1,n219_0,n244_1,n212_1,n212_0,n209_1,n209_0,n115_1,n66_2,n66_0,n203_2,n203_1,n99_4,n99_0,n229_1,n190_4,n229_0,n190_3,_w_797,n190_2,n189_1,n200_3,n200_1,n200_0,n188_0,n251,n99_1,n80,n68_1,_w_617,n98_0,n232,n89_0,n230,n154_1,n227,n197_1,n174_1,n239,n134,n225,n165_0,n164_0,n220,n179_0,n219,n217,n212,n209,n208,_w_610,n115,n66_1,n203,n75_1,n191,n229,n228,n190,_w_801,_w_791,n125_0,n189,n188,_w_759,n245,n238,n181_0,_w_749,n180,n177,n218,n94_1,n173,n171,n98,n167,n166,n165,n164,n74,n160,n214,n185,n137_0,n143,n158_3,n193,n136_1,n157,n86_2,n175_3,n155,n84_1,_w_743,n236,n151,n202,n147,_w_622,n145,n105_1,n87_1,n144,n207,_w_679,n140,_w_760,n138,n111_0,n204,n66,n78_1,n168,n235_1,n118,n218_1,n86_0,n182_1,n135,_w_711,n167_0,n133,n165_3,n86_1,n81_1,n175,n130,n129,n132,n196,n190_1,n146,_w_675,n256,n127,n239_0,n125,n125_1,_w_715,n122,n107,n147_0,n121,n99,n150,_w_676,n165_4,n69,n252,n188_1,n156,n116_2,n242,n221,n206,_w_792,n189_0,n126,n84_0,n130_1,n246,n237,n102_1,_w_764,_w_652,_w_630,n101,n137,n98_1,n123,n149,n174_2,n243,n195_1,n118_1,_w_657,n92,n248,n128,n129_1,n74_0,n181,_w_625,n115_0,n113_2,n133_3,n213,n88,n158,n90_2,n160_1,_w_709,n109,_w_678,n239_2,n136,n216,n102_0,_w_722,_w_638,n256_1,_w_600,n219_3,n233,n111,n130_0,n68,n120,n89,n211,n88_0,n192,n158_1,n172,n131,n75,n67_1,n89_1,n138_1,n112,n165_2,n102,n100,n71,n164_1,n255,n254,n108,_w_658,n240,_w_789,n84,n67_0,n192_0,_w_790,n172_1,n146_0,n232_0,n67,_w_609,n110_2,n154,n178,n163_0,n93,_w_626,n99_2,n167_1,_w_683,n113_3,_w_695,n111_1,n92_1,_w_763,n174,n70,_w_624,n104,n82,n179,n187,_w_779,n108_0,n186,n110,n76,n91,n179_3,n65,n72,n176,_w_674,n244_0,n197_0,n77,_w_730,n183,n142_3,n116,_w_687,_w_752,n78,_w_726,n195,n79_2,n156_0,_w_798,n83,_w_736,n161,n85,n87,n86,n119_1,n87_2,n146_2,n154_3,n132_0,n119,n226_1,n157_1,n94,n224_2,_w_737,n95,n85_0,n79,n96,n142_2,n122_0,n219_2,n97,n234,n103,n199,n90,n109_1,n122_4,n162,n127_1,_w_639,n106,n113,n137_1,n184,n223_2,n257,n258,n158_2,n70_0,n113_0,n235,n113_1,n90_0,_w_795,n90_1,n163_1,n90_3,n200_2,n223_0,n105_0,n226,n72_1,n73_2,n105_2,n105_3,n183_4,n210,n199_0,n65_1,n199_1,n223_1,n199_2,_w_616,n82_1,_w_787,n88_1,n96_2,n96_0,n96_1,n96_3,n79_0,n129_2,n79_1,n79_4,n160_2,n95_1,n119_0,n124_1,n157_0,_w_724,n185_0,n119_2,_w_719,n119_3,n197_2,n87_0,_w_741,_w_651,n161_0,n141,n161_1,n73,n161_2,_w_782,n182,n161_3,_w_620,n81_0,n116_0,n72_0,n76_0,n76_1,n76_2,n226_0,n76_3,_w_725,n110_0,n110_1,n82_2,n154_0,n175_0,n186_0,n186_1,n186_2,n144_1,_w_603,n159,n105_4,n179_1,n190_0,n148,n179_2,n224,n82_0,n70_1,_w_785,n70_3,n215_0,n175_1,_w_619,n138_0,n93_1,_w_718,n101_0,n186_3,n93_2,n178_0,n146_1,n178_1,n178_2,_w_761,_w_746,n152,n65_0,n67_2,_w_653,n117_0,n117_1,_w_649,n136_0,n240_0,_w_701,n231,n240_1,n185_2,n142,n108_1,n240_2,_w_633,n139_0,_w_700,n158_0,n158_4,_w_802,_w_773,n157_2,n183_2,n194,n132_1,n139_2,n139_3,n225_2,n151_1,n201,n102_2,_w_659,n112_0,n112_1,n215,n151_5,n95_0,n75_0,n172_0,_w_604,n172_2,n192_1,n192_2,_w_805,_w_720,n195_0,n68_0,n135_0,n142_0,n203_0,n85_1,n73_1,n142_1,n109_0,n148_1,n109_2,n81,n181_1,n92_0,n101_1,n170,n206_0,n99_3,n206_1,_w_682,n69_1,n156_1,_w_703,_w_697,n69_0,n198,n79_3,n121_0,n130_2,n78_0,n150_1,n124_0,n93_0,n150_0,n175_2,n121_1,n116_1,n122_1,n122_2,n122_3,n174_0,n125_2,n127_0,n169,n128_0,n244,n128_1,n70_2,n129_0,n232_2,n205,n131_1,n215_1,n250_1,n131_0,n249,n114,n224_0,n200,n151_4,n224_1,n189_2,n250_0,n139_1,n133_0,n133_1,n133_2,n73_0,n135_1,_w_742,n223,n118_0,n136_2,n104_0,n250,n141_0,n141_1,_w_717,n94_0,n144_0,_w_642,_w_621,n147_1,n148_0,_w_793,n148_2,n148_3,n148_4,n151_0,_w_602,n151_2,n151_3,n142_4,n170_0,n212_2,n154_2,n185_1,_w_681,n160_0,n104_1,n74_1,n124,n117,n197,n164_2,n165_1,n167_2,n163,n105,n218_0,n218_2,n182_0,n139,n182_2,n183_1,_w_690,n183_0,n183_3,_w_738,n170_1,n256_0;

  bfr _b_544(.a(_w_803),.q(n139_1));
  bfr _b_541(.a(_w_800),.q(out_2_));
  spl3L g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1),.q2(_w_804));
  spl2 g68_s_0(.a(n68),.q0(n68_0),.q1(n68_1));
  spl3L g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1),.q2(n192_2));
  spl2 g139_s_0(.a(n139),.q0(n139_0),.q1(_w_801));
  bfr _b_471(.a(_w_730),.q(_w_731));
  bfr _b_348(.a(_w_607),.q(n66_2));
  spl2 g84_s_0(.a(n84),.q0(n84_0),.q1(n84_1));
  and_bi g247(.a(n246),.b(n245),.q(_w_798));
  spl2 g70_s_0(.a(n70),.q0(n70_0),.q1(_w_795));
  spl3L g102_s_0(.a(n102),.q0(n102_0),.q1(n102_1),.q2(n102_2));
  bfr _b_417(.a(_w_676),.q(n110_2));
  spl2 g72_s_0(.a(n72),.q0(n72_0),.q1(n72_1));
  and_bb g89(.a(in_18_),.b(in_19_),.q(n89));
  bfr _b_458(.a(_w_717),.q(_w_718));
  bfr _b_533(.a(_w_792),.q(_w_793));
  bfr _b_507(.a(_w_766),.q(_w_767));
  spl2 g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1));
  spl2 g108_s_0(.a(n108),.q0(n108_0),.q1(n108_1));
  and_bb g85(.a(in_30_),.b(in_31_),.q(_w_782));
  bfr _b_462(.a(_w_721),.q(_w_722));
  bfr _b_442(.a(_w_701),.q(_w_702));
  spl3L g87_s_0(.a(n87),.q0(n87_0),.q1(n87_1),.q2(_w_780));
  or_bb g221(.a(n206_1),.b(n219_3),.q(n221));
  and_bb g116(.a(in_42_),.b(in_43_),.q(n116));
  spl2 g186_s_0(.a(n186),.q0(n186_0),.q1(_w_777));
  bfr _b_545(.a(_w_804),.q(_w_805));
  spl3L g178_s_0(.a(n178),.q0(n178_0),.q1(n178_1),.q2(n178_2));
  spl2 g113_s_1(.a(n113_1),.q0(n113_2),.q1(_w_774));
  and_bb g213(.a(n197_1),.b(n199_1),.q(n213));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(_w_768));
  and_bi g244(.a(n243),.b(n242),.q(n244));
  or_bb g177(.a(n170_1),.b(n175_3),.q(n177));
  or_bb g243(.a(n212_2),.b(n218_2),.q(n243));
  maj_bbb g142(.a(n129_0),.b(n135_0),.c(n141_0),.q(n142));
  and_bb g242(.a(n212_1),.b(n218_1),.q(n242));
  and_bi g235(.a(n234),.b(n233),.q(n235));
  and_bb g233(.a(n183_2),.b(n190_2),.q(n233));
  and_bi g232(.a(n231),.b(n230),.q(n232));
  spl2 g175_s_1(.a(n175_1),.q0(n175_2),.q1(n175_3));
  spl2 g89_s_0(.a(n89),.q0(n89_0),.q1(n89_1));
  or_bb g231(.a(n223_2),.b(n229_1),.q(n231));
  bfr _b_439(.a(_w_698),.q(_w_699));
  maj_bbb g219(.a(n151_2),.b(n212_0),.c(n218_0),.q(n219));
  and_bi g238(.a(n237),.b(n236),.q(n238));
  maj_bbi g121(.a(n116_2),.b(n120),.c(n119_0),.q(n121));
  and_bb g69(.a(in_2_),.b(in_3_),.q(n69));
  bfr _b_531(.a(_w_790),.q(_w_791));
  and_bb g227(.a(n158_2),.b(n165_2),.q(n227));
  maj_bbb g224(.a(n158_4),.b(n165_4),.c(n223_0),.q(_w_760));
  or_bb g205(.a(n178_1),.b(n203_1),.q(n205));
  or_bb g68(.a(in_0_),.b(in_1_),.q(n68));
  maj_bbb g223(.a(n160_2),.b(n167_2),.c(n175_0),.q(n223));
  spl2 g79_s_1(.a(n79_2),.q0(n79_3),.q1(_w_759));
  and_bb g117(.a(in_38_),.b(in_39_),.q(n117));
  and_bb g148(.a(n127_0),.b(n147_0),.q(n148));
  bfr _b_343(.a(_w_602),.q(n238_2));
  and_bi g229(.a(n228),.b(n227),.q(n229));
  or_bb g237(.a(n225_2),.b(n235_1),.q(n237));
  maj_bbi g81(.a(n66_2),.b(n80),.c(n79_0),.q(n81));
  and_bi g218(.a(n217),.b(n216),.q(n218));
  or_bb g217(.a(n148_4),.b(n215_1),.q(n217));
  maj_bbb g225(.a(n185_2),.b(n192_2),.c(n200_0),.q(n225));
  spl3L g240_s_0(.a(n240),.q0(n240_0),.q1(n240_1),.q2(n240_2));
  spl2 g215_s_0(.a(n215),.q0(n215_0),.q1(n215_1));
  and_bi g215(.a(n214),.b(n213),.q(n215));
  bfr _b_460(.a(_w_719),.q(n99_4));
  or_bb g214(.a(n197_2),.b(n199_2),.q(n214));
  or_bb g67(.a(in_4_),.b(in_5_),.q(n67));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(_w_756));
  or_bb g211(.a(n105_4),.b(n209_1),.q(n211));
  spl3L g223_s_0(.a(n223),.q0(n223_0),.q1(n223_1),.q2(n223_2));
  or_bb g159(.a(n154_3),.b(n157_2),.q(_w_755));
  spl2 g119_s_1(.a(n119_1),.q0(n119_2),.q1(_w_754));
  bfr _b_503(.a(_w_762),.q(n224));
  and_bb g210(.a(n105_3),.b(n209_0),.q(n210));
  bfr _b_437(.a(_w_696),.q(n67_2));
  and_bb g207(.a(n172_1),.b(n174_1),.q(n207));
  and_bi g206(.a(n205),.b(n204),.q(n206));
  maj_bbi g71(.a(n68_1),.b(n69_1),.c(n67_1),.q(_w_751));
  or_bb g258(.a(n240_1),.b(n256_1),.q(n258));
  and_bb g82(.a(n65_0),.b(n81_0),.q(n82));
  maj_bbb g226(.a(n183_4),.b(n190_4),.c(n225_0),.q(_w_748));
  bfr _b_466(.a(_w_725),.q(n183_4));
  spl2 g161_s_0(.a(n161),.q0(n161_0),.q1(_w_742));
  and_bi g199(.a(n198),.b(n189_1),.q(n199));
  spl2 g163_s_0(.a(n163),.q0(n163_0),.q1(n163_1));
  bfr _b_382(.a(_w_641),.q(_w_642));
  spl2 g139_s_1(.a(n139_1),.q0(n139_2),.q1(_w_741));
  maj_bbi g187(.a(n133_3),.b(n139_3),.c(n142_3),.q(n187));
  or_bb g196(.a(n125_2),.b(n181_1),.q(_w_740));
  spl2 g70_s_1(.a(n70_1),.q0(n70_2),.q1(_w_739));
  maj_bbi g120(.a(n117_1),.b(n118_1),.c(n116_1),.q(_w_737));
  spl2 g179_s_1(.a(n179_1),.q0(n179_2),.q1(n179_3));
  or_bb g118(.a(in_40_),.b(in_41_),.q(n118));
  spl2 g95_s_0(.a(n95),.q0(n95_0),.q1(n95_1));
  or_bb g166(.a(n161_3),.b(n164_2),.q(_w_736));
  and_bi g104(.a(n103),.b(n102_0),.q(n104));
  or_bb g234(.a(n183_3),.b(n190_3),.q(n234));
  spl2 g181_s_0(.a(n181),.q0(n181_0),.q1(n181_1));
  and_bb g112(.a(in_34_),.b(in_35_),.q(n112));
  bfr _b_368(.a(_w_627),.q(n130_2));
  or_bb g228(.a(n158_3),.b(n165_3),.q(n228));
  and_bb g216(.a(n148_3),.b(n215_0),.q(n216));
  and_bb g108(.a(in_46_),.b(in_47_),.q(_w_728));
  or_bb g111(.a(in_32_),.b(in_33_),.q(n111));
  spl3L g86_s_0(.a(n86),.q0(n86_0),.q1(n86_1),.q2(_w_726));
  or_bb g75(.a(in_8_),.b(in_9_),.q(n75));
  spl2 g206_s_0(.a(n206),.q0(n206_0),.q1(n206_1));
  spl2 g94_s_0(.a(n94),.q0(n94_0),.q1(n94_1));
  or_bb g249(.a(n232_1),.b(n238_1),.q(n249));
  and_bb g157(.a(n156_0),.b(n82_1),.q(n157));
  spl2 g124_s_0(.a(n124),.q0(n124_0),.q1(n124_1));
  bfr _b_356(.a(_w_615),.q(_w_616));
  and_bb g201(.a(n195_0),.b(n200_2),.q(n201));
  maj_bbb g113(.a(n110_0),.b(n111_0),.c(n112_0),.q(n113));
  maj_bbb g79(.a(n66_0),.b(n72_0),.c(n78_0),.q(n79));
  and_bb g164(.a(n102_1),.b(n163_0),.q(n164));
  spl3L g73_s_0(.a(n73),.q0(n73_0),.q1(n73_1),.q2(_w_792));
  and_bb g102(.a(n101_0),.b(n85_0),.q(n102));
  and_bb g168(.a(n160_0),.b(n167_0),.q(n168));
  or_bb g208(.a(n172_2),.b(n174_2),.q(n208));
  spl3L g183_s_1(.a(n183_1),.q0(n183_2),.q1(n183_3),.q2(_w_723));
  and_bb g236(.a(n225_1),.b(n235_0),.q(n236));
  bfr _b_386(.a(_w_645),.q(_w_646));
  and_bi g256(.a(n255),.b(n254),.q(n256));
  spl2 g76_s_0(.a(n76),.q0(n76_0),.q1(_w_765));
  bfr _b_423(.a(_w_682),.q(out_6_));
  maj_bbb g119(.a(n116_0),.b(n117_0),.c(n118_0),.q(n119));
  spl2 g99_s_1(.a(n99_2),.q0(n99_3),.q1(_w_719));
  maj_bbb g99(.a(n86_0),.b(n92_0),.c(n98_0),.q(n99));
  bfr _b_496(.a(_w_755),.q(n159));
  bfr _b_431(.a(_w_690),.q(_w_691));
  spl2 g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1));
  and_bb g146(.a(n128_1),.b(n144_1),.q(n146));
  bfr _b_376(.a(_w_635),.q(n171));
  spl3L g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1),.q2(n199_2));
  spl2 g105_s_1(.a(n105_2),.q0(n105_3),.q1(n105_4));
  and_bi g212(.a(n211),.b(n210),.q(n212));
  maj_bbb g70(.a(n67_0),.b(n68_0),.c(n69_0),.q(n70));
  or_bb g202(.a(n195_1),.b(n200_3),.q(n202));
  bfr _b_350(.a(_w_609),.q(n219_1));
  bfr _b_492(.a(_w_751),.q(n71));
  maj_bbi g77(.a(n74_1),.b(n75_1),.c(n73_1),.q(_w_714));
  maj_bbb g175(.a(n105_1),.b(n172_0),.c(n174_0),.q(n175));
  or_bb g198(.a(n146_2),.b(n188_1),.q(_w_713));
  bfr _b_525(.a(_w_784),.q(_w_785));
  or_bb g169(.a(n160_1),.b(n167_1),.q(n169));
  maj_bbb g239(.a(n178_2),.b(n203_2),.c(n219_0),.q(n239));
  bfr _b_453(.a(_w_712),.q(n114));
  and_bb g220(.a(n206_0),.b(n219_2),.q(n220));
  and_bi g222(.a(n221),.b(n220),.q(_w_711));
  or_bb g106(.a(n104_1),.b(n84_1),.q(_w_710));
  and_bb g74(.a(in_6_),.b(in_7_),.q(n74));
  or_bb g66(.a(in_12_),.b(in_13_),.q(_w_704));
  or_bb g246(.a(n151_5),.b(n244_1),.q(n246));
  spl2 g81_s_0(.a(n81),.q0(n81_0),.q1(n81_1));
  and_bb g136(.a(in_58_),.b(in_59_),.q(n136));
  maj_bbi g92(.a(n87_2),.b(n91),.c(n90_0),.q(n92));
  spl3L g232_s_0(.a(n232),.q0(n232_0),.q1(n232_1),.q2(_w_701));
  spl2 g76_s_1(.a(n76_1),.q0(n76_2),.q1(_w_794));
  and_bb g183(.a(n179_2),.b(n182_0),.q(n183));
  spl2 g90_s_0(.a(n90),.q0(n90_0),.q1(_w_698));
  maj_bbb g96(.a(n93_0),.b(n94_0),.c(n95_0),.q(n96));
  bfr _b_425(.a(_w_684),.q(_w_685));
  and_bb g73(.a(in_10_),.b(in_11_),.q(n73));
  and_bb g245(.a(n151_4),.b(n244_0),.q(n245));
  spl2 g85_s_0(.a(n85),.q0(n85_0),.q1(n85_1));
  spl3L g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1),.q2(n182_2));
  bfr _b_387(.a(_w_646),.q(out_1_));
  and_bi g107(.a(n106),.b(n105_0),.q(n107));
  maj_bbb g76(.a(n73_0),.b(n74_0),.c(n75_0),.q(n76));
  bfr _b_512(.a(_w_771),.q(_w_772));
  maj_bbi g100(.a(n92_1),.b(n98_1),.c(n86_1),.q(_w_697));
  spl3L g67_s_0(.a(n67),.q0(n67_0),.q1(n67_1),.q2(_w_695));
  maj_bbi g80(.a(n72_1),.b(n78_1),.c(n66_1),.q(_w_694));
  or_bb g87(.a(in_20_),.b(in_21_),.q(n87));
  and_bi g84(.a(n83),.b(n82_0),.q(n84));
  and_bb g94(.a(in_22_),.b(in_23_),.q(n94));
  maj_bbi g143(.a(n135_1),.b(n141_1),.c(n129_1),.q(_w_692));
  bfr _b_344(.a(_w_603),.q(_w_604));
  maj_bbb g122(.a(n109_0),.b(n115_0),.c(n121_0),.q(n122));
  and_bb g165(.a(n161_2),.b(n164_0),.q(n165));
  bfr _b_506(.a(_w_765),.q(_w_766));
  or_bb g109(.a(in_44_),.b(in_45_),.q(_w_688));
  or_bb g86(.a(in_28_),.b(in_29_),.q(_w_684));
  and_bi g197(.a(n196),.b(n182_1),.q(n197));
  bfr _b_406(.a(_w_665),.q(n129));
  spl2 g132_s_0(.a(n132),.q0(n132_0),.q1(n132_1));
  maj_bbi g91(.a(n88_1),.b(n89_1),.c(n87_1),.q(_w_683));
  spl2 g148_s_1(.a(n148_2),.q0(n148_3),.q1(n148_4));
  spl2 g131_s_0(.a(n131),.q0(n131_0),.q1(n131_1));
  maj_bbb g241(.a(n224_2),.b(n226_2),.c(n240_2),.q(_w_682));
  bfr _b_363(.a(_w_622),.q(_w_623));
  maj_bbi g134(.a(n131_1),.b(n132_1),.c(n130_1),.q(_w_681));
  and_bi g259(.a(n258),.b(n257),.q(out_5_));
  maj_bbi g123(.a(n115_1),.b(n121_1),.c(n109_1),.q(_w_680));
  spl2 g118_s_0(.a(n118),.q0(n118_0),.q1(n118_1));
  and_bb g204(.a(n178_0),.b(n203_0),.q(n204));
  spl2 g96_s_1(.a(n96_1),.q0(n96_2),.q1(_w_679));
  maj_bbi g124(.a(n109_2),.b(n123),.c(n122_0),.q(n124));
  or_bb g194(.a(n185_1),.b(n192_1),.q(n194));
  and_bb g125(.a(n108_0),.b(n124_0),.q(n125));
  bfr _b_427(.a(_w_686),.q(_w_687));
  bfr _b_475(.a(_w_734),.q(_w_735));
  bfr _b_443(.a(_w_702),.q(_w_703));
  or_bb g255(.a(n224_1),.b(n226_1),.q(n255));
  bfr _b_459(.a(_w_718),.q(n96_1));
  and_bi g195(.a(n194),.b(n193),.q(n195));
  spl3L g129_s_0(.a(n129),.q0(n129_0),.q1(n129_1),.q2(_w_677));
  spl3L g110_s_0(.a(n110),.q0(n110_0),.q1(n110_1),.q2(_w_675));
  or_bb g126(.a(n108_1),.b(n124_1),.q(_w_674));
  and_bi g127(.a(n126),.b(n125_0),.q(n127));
  and_bb g193(.a(n185_0),.b(n192_0),.q(n193));
  and_bb g128(.a(in_62_),.b(in_63_),.q(_w_666));
  or_bb g129(.a(in_60_),.b(in_61_),.q(_w_662));
  and_bb g248(.a(n232_0),.b(n238_0),.q(n248));
  or_bb g130(.a(in_52_),.b(in_53_),.q(n130));
  or_bb g152(.a(n107_1),.b(n150_1),.q(_w_661));
  spl2 g161_s_1(.a(n161_1),.q0(n161_2),.q1(n161_3));
  and_bb g254(.a(n224_0),.b(n226_0),.q(n254));
  bfr _b_444(.a(_w_703),.q(n232_2));
  or_bb g103(.a(n101_1),.b(n85_1),.q(_w_660));
  and_bb g230(.a(n223_1),.b(n229_0),.q(n230));
  bfr _b_491(.a(_w_750),.q(n226));
  and_bi g160(.a(n159),.b(n158_0),.q(n160));
  bfr _b_416(.a(_w_675),.q(_w_676));
  and_bi g250(.a(n249),.b(n248),.q(n250));
  and_bi g174(.a(n173),.b(n164_1),.q(n174));
  spl3L g116_s_0(.a(n116),.q0(n116_0),.q1(n116_1),.q2(_w_790));
  bfr _b_487(.a(_w_746),.q(_w_747));
  and_bi g209(.a(n208),.b(n207),.q(n209));
  or_bb g95(.a(in_24_),.b(in_25_),.q(n95));
  bfr _b_384(.a(_w_643),.q(_w_644));
  bfr _b_370(.a(_w_629),.q(_w_630));
  spl3L g203_s_0(.a(n203),.q0(n203_0),.q1(n203_1),.q2(n203_2));
  maj_bbb g200(.a(n148_1),.b(n197_0),.c(n199_0),.q(n200));
  maj_bbb g154(.a(n70_2),.b(n76_2),.c(n79_1),.q(n154));
  spl2 g133_s_0(.a(n133),.q0(n133_0),.q1(_w_657));
  and_bb g137(.a(in_54_),.b(in_55_),.q(n137));
  spl2 g115_s_0(.a(n115),.q0(n115_0),.q1(n115_1));
  bfr _b_375(.a(_w_634),.q(n173));
  bfr _b_529(.a(_w_788),.q(_w_789));
  spl3L g79_s_0(.a(n79),.q0(n79_0),.q1(n79_1),.q2(n79_2));
  bfr _b_451(.a(_w_710),.q(n106));
  spl2 g104_s_0(.a(n104),.q0(n104_0),.q1(n104_1));
  maj_bbi g140(.a(n137_1),.b(n138_1),.c(n136_1),.q(_w_656));
  bfr _b_474(.a(_w_733),.q(_w_734));
  bfr _b_361(.a(_w_620),.q(n133_3));
  maj_bbi g144(.a(n129_2),.b(n143),.c(n142_0),.q(n144));
  bfr _b_412(.a(_w_671),.q(_w_672));
  and_bb g151(.a(n107_0),.b(n150_0),.q(n151));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(n250_1));
  spl2 g113_s_0(.a(n113),.q0(n113_0),.q1(_w_771));
  bfr _b_498(.a(_w_757),.q(_w_758));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(n112_1));
  maj_bbb g139(.a(n136_0),.b(n137_0),.c(n138_0),.q(n139));
  bfr _b_369(.a(_w_628),.q(n122_4));
  and_bb g65(.a(in_14_),.b(in_15_),.q(_w_647));
  maj_bbb g240(.a(n232_2),.b(n238_2),.c(n239_0),.q(n240));
  and_bi g147(.a(n145),.b(n146_0),.q(n147));
  bfr _b_420(.a(_w_679),.q(n96_3));
  bfr _b_411(.a(_w_670),.q(_w_671));
  maj_bbi g115(.a(n110_2),.b(n114),.c(n113_0),.q(n115));
  and_bi g153(.a(n152),.b(n151_0),.q(_w_638));
  maj_bbi g155(.a(n70_3),.b(n76_3),.c(n79_3),.q(n155));
  spl2 g186_s_1(.a(n186_1),.q0(n186_2),.q1(n186_3));
  spl3L g136_s_0(.a(n136),.q0(n136_0),.q1(n136_1),.q2(_w_636));
  spl3L g99_s_0(.a(n99),.q0(n99_0),.q1(n99_1),.q2(n99_2));
  bfr _b_440(.a(_w_699),.q(_w_700));
  and_bb g190(.a(n186_2),.b(n189_0),.q(n190));
  spl2 g121_s_0(.a(n121),.q0(n121_0),.q1(n121_1));
  and_bb g158(.a(n154_2),.b(n157_0),.q(n158));
  bfr _b_438(.a(_w_697),.q(n100));
  maj_bbb g161(.a(n90_2),.b(n96_2),.c(n99_1),.q(n161));
  maj_bbi g162(.a(n90_3),.b(n96_3),.c(n99_3),.q(n162));
  bfr _b_449(.a(_w_708),.q(_w_709));
  and_bi g185(.a(n184),.b(n183_0),.q(n185));
  bfr _b_452(.a(_w_711),.q(out_3_));
  maj_bbi g163(.a(n162),.b(n99_4),.c(n161_0),.q(n163));
  spl2 g92_s_0(.a(n92),.q0(n92_0),.q1(n92_1));
  spl3L g82_s_0(.a(n82),.q0(n82_0),.q1(n82_1),.q2(n82_2));
  maj_bbb g179(.a(n113_2),.b(n119_2),.c(n122_1),.q(n179));
  bfr _b_521(.a(_w_780),.q(_w_781));
  and_bi g167(.a(n166),.b(n165_0),.q(n167));
  and_bi g170(.a(n169),.b(n168),.q(n170));
  bfr _b_441(.a(_w_700),.q(n90_1));
  bfr _b_405(.a(_w_664),.q(_w_665));
  maj_bbi g98(.a(n93_2),.b(n97),.c(n96_0),.q(n98));
  maj_bbi g78(.a(n73_2),.b(n77),.c(n76_0),.q(n78));
  bfr _b_502(.a(_w_761),.q(_w_762));
  or_bb g171(.a(n156_1),.b(n82_2),.q(_w_635));
  bfr _b_527(.a(_w_786),.q(_w_787));
  or_bb g252(.a(n239_2),.b(n250_1),.q(n252));
  bfr _b_349(.a(_w_608),.q(_w_609));
  spl2 g195_s_0(.a(n195),.q0(n195_0),.q1(n195_1));
  or_bb g173(.a(n102_2),.b(n163_1),.q(_w_634));
  spl2 g142_s_1(.a(n142_2),.q0(n142_3),.q1(_w_633));
  bfr _b_429(.a(_w_688),.q(_w_689));
  or_bb g110(.a(in_36_),.b(in_37_),.q(n110));
  and_bb g257(.a(n240_0),.b(n256_0),.q(n257));
  maj_bbi g101(.a(n100),.b(n86_2),.c(n99_0),.q(n101));
  maj_bbi g180(.a(n113_3),.b(n119_3),.c(n122_3),.q(n180));
  spl3L g93_s_0(.a(n93),.q0(n93_0),.q1(n93_1),.q2(_w_708));
  and_bi g178(.a(n177),.b(n176),.q(n178));
  maj_bbb g186(.a(n133_2),.b(n139_2),.c(n142_1),.q(n186));
  maj_bbb g133(.a(n130_0),.b(n131_0),.c(n132_0),.q(n133));
  maj_bbb g90(.a(n87_0),.b(n88_0),.c(n89_0),.q(n90));
  or_bb g184(.a(n179_3),.b(n182_2),.q(_w_632));
  spl3L g190_s_1(.a(n190_1),.q0(n190_2),.q1(n190_3),.q2(_w_629));
  bfr _b_413(.a(_w_672),.q(_w_673));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(n88_1));
  spl2 g101_s_0(.a(n101),.q0(n101_0),.q1(n101_1));
  spl3L g125_s_0(.a(n125),.q0(n125_0),.q1(n125_1),.q2(n125_2));
  bfr _b_515(.a(_w_774),.q(n113_3));
  spl3L g174_s_0(.a(n174),.q0(n174_0),.q1(n174_1),.q2(n174_2));
  spl2 g156_s_0(.a(n156),.q0(n156_0),.q1(n156_1));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  maj_bbi g141(.a(n136_2),.b(n140),.c(n139_0),.q(n141));
  spl3L g122_s_0(.a(n122),.q0(n122_0),.q1(n122_1),.q2(n122_2));
  bfr _b_403(.a(_w_662),.q(_w_663));
  spl2 g122_s_1(.a(n122_2),.q0(n122_3),.q1(_w_628));
  spl2 g127_s_0(.a(n127),.q0(n127_0),.q1(n127_1));
  spl3L g146_s_0(.a(n146),.q0(n146_0),.q1(n146_1),.q2(n146_2));
  and_bi g192(.a(n191),.b(n190_0),.q(n192));
  bfr _b_407(.a(_w_666),.q(_w_667));
  bfr _b_341(.a(_w_600),.q(_w_601));
  or_bb g83(.a(n65_1),.b(n81_1),.q(_w_693));
  spl2 g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1));
  spl3L g130_s_0(.a(n130),.q0(n130_0),.q1(n130_1),.q2(_w_626));
  bfr _b_430(.a(_w_689),.q(_w_690));
  spl2 g111_s_0(.a(n111),.q0(n111_0),.q1(n111_1));
  spl2 g175_s_0(.a(n175),.q0(n175_0),.q1(_w_624));
  spl2 g117_s_0(.a(n117),.q0(n117_0),.q1(n117_1));
  spl3L g157_s_0(.a(n157),.q0(n157_0),.q1(n157_1),.q2(n157_2));
  maj_bbi g72(.a(n67_2),.b(n71),.c(n70_0),.q(n72));
  bfr _b_472(.a(_w_731),.q(_w_732));
  spl3L g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1),.q2(n142_2));
  spl3L g224_s_0(.a(n224),.q0(n224_0),.q1(n224_1),.q2(_w_621));
  spl2 g133_s_1(.a(n133_1),.q0(n133_2),.q1(_w_620));
  spl2 g135_s_0(.a(n135),.q0(n135_0),.q1(n135_1));
  bfr _b_389(.a(_w_648),.q(_w_649));
  and_bb g105(.a(n104_0),.b(n84_0),.q(n105));
  and_bi g203(.a(n202),.b(n201),.q(n203));
  spl2 g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1));
  and_bi g172(.a(n171),.b(n157_1),.q(n172));
  spl2 g138_s_0(.a(n138),.q0(n138_0),.q1(n138_1));
  spl2 g141_s_0(.a(n141),.q0(n141_0),.q1(n141_1));
  spl2 g147_s_0(.a(n147),.q0(n147_0),.q1(n147_1));
  spl3L g148_s_0(.a(n148),.q0(n148_0),.q1(n148_1),.q2(_w_618));
  spl3L g239_s_0(.a(n239),.q0(n239_0),.q1(n239_1),.q2(n239_2));
  or_bb g88(.a(in_16_),.b(in_17_),.q(n88));
  spl2 g151_s_0(.a(n151),.q0(n151_0),.q1(_w_617));
  spl2 g229_s_0(.a(n229),.q0(n229_0),.q1(n229_1));
  bfr _b_352(.a(_w_611),.q(n200_1));
  and_bb g176(.a(n170_0),.b(n175_2),.q(n176));
  spl2 g151_s_1(.a(n151_1),.q0(n151_2),.q1(_w_615));
  bfr _b_393(.a(_w_652),.q(_w_653));
  spl2 g170_s_0(.a(n170),.q0(n170_0),.q1(n170_1));
  spl2 g154_s_1(.a(n154_1),.q0(n154_2),.q1(n154_3));
  spl3L g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1),.q2(n185_2));
  spl3L g160_s_0(.a(n160),.q0(n160_0),.q1(n160_1),.q2(n160_2));
  spl3L g164_s_0(.a(n164),.q0(n164_0),.q1(n164_1),.q2(n164_2));
  spl3L g165_s_1(.a(n165_1),.q0(n165_2),.q1(n165_3),.q2(_w_612));
  spl3L g167_s_0(.a(n167),.q0(n167_0),.q1(n167_1),.q2(n167_2));
  spl2 g98_s_0(.a(n98),.q0(n98_0),.q1(n98_1));
  spl3L g218_s_0(.a(n218),.q0(n218_0),.q1(n218_1),.q2(n218_2));
  spl2 g183_s_0(.a(n183),.q0(n183_0),.q1(n183_1));
  bfr _b_408(.a(_w_667),.q(_w_668));
  spl2 g200_s_0(.a(n200),.q0(n200_0),.q1(_w_610));
  bfr _b_543(.a(_w_802),.q(_w_803));
  spl2 g219_s_0(.a(n219),.q0(n219_0),.q1(_w_608));
  bfr _b_546(.a(_w_805),.q(n109_2));
  bfr _b_456(.a(_w_715),.q(n149));
  spl2 g200_s_1(.a(n200_1),.q0(n200_2),.q1(n200_3));
  and_bb g189(.a(n146_1),.b(n188_0),.q(n189));
  spl3L g66_s_0(.a(n66),.q0(n66_0),.q1(n66_1),.q2(_w_606));
  spl2 g209_s_0(.a(n209),.q0(n209_0),.q1(n209_1));
  spl2 g96_s_0(.a(n96),.q0(n96_0),.q1(_w_716));
  spl3L g212_s_0(.a(n212),.q0(n212_0),.q1(n212_1),.q2(n212_2));
  bfr _b_345(.a(_w_604),.q(_w_605));
  spl2 g256_s_0(.a(n256),.q0(n256_0),.q1(n256_1));
  spl2 g244_s_0(.a(n244),.q0(n244_0),.q1(n244_1));
  bfr _b_373(.a(_w_632),.q(n184));
  spl2 g219_s_1(.a(n219_1),.q0(n219_2),.q1(n219_3));
  spl2 g74_s_0(.a(n74),.q0(n74_0),.q1(n74_1));
  spl3L g225_s_0(.a(n225),.q0(n225_0),.q1(n225_1),.q2(n225_2));
  bfr _b_461(.a(_w_720),.q(_w_721));
  spl3L g226_s_0(.a(n226),.q0(n226_0),.q1(n226_1),.q2(_w_603));
  spl2 g107_s_0(.a(n107),.q0(n107_0),.q1(n107_1));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(n235_1));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(n75_1));
  spl3L g238_s_0(.a(n238),.q0(n238_0),.q1(n238_1),.q2(_w_600));
  bfr _b_342(.a(_w_601),.q(_w_602));
  bfr _b_346(.a(_w_605),.q(n226_2));
  bfr _b_347(.a(_w_606),.q(_w_607));
  and_bi g253(.a(n252),.b(n251),.q(_w_752));
  bfr _b_501(.a(_w_760),.q(_w_761));
  bfr _b_351(.a(_w_610),.q(_w_611));
  bfr _b_354(.a(_w_613),.q(_w_614));
  spl3L g105_s_0(.a(n105),.q0(n105_0),.q1(n105_1),.q2(_w_775));
  bfr _b_374(.a(_w_633),.q(n142_4));
  bfr _b_419(.a(_w_678),.q(n129_2));
  bfr _b_355(.a(_w_614),.q(n165_4));
  bfr _b_540(.a(_w_799),.q(_w_800));
  bfr _b_357(.a(_w_616),.q(n151_3));
  spl2 g90_s_1(.a(n90_1),.q0(n90_2),.q1(_w_763));
  bfr _b_509(.a(_w_768),.q(_w_769));
  bfr _b_479(.a(_w_738),.q(n191));
  or_bb g131(.a(in_48_),.b(in_49_),.q(n131));
  bfr _b_358(.a(_w_617),.q(n151_1));
  spl2 g158_s_0(.a(n158),.q0(n158_0),.q1(n158_1));
  and_bi g150(.a(n149),.b(n148_0),.q(n150));
  bfr _b_359(.a(_w_618),.q(_w_619));
  bfr _b_360(.a(_w_619),.q(n148_2));
  spl2 g65_s_0(.a(n65),.q0(n65_0),.q1(n65_1));
  bfr _b_362(.a(_w_621),.q(_w_622));
  bfr _b_364(.a(_w_623),.q(n224_2));
  spl2 g154_s_0(.a(n154),.q0(n154_0),.q1(_w_720));
  bfr _b_500(.a(_w_759),.q(n79_4));
  bfr _b_365(.a(_w_624),.q(_w_625));
  bfr _b_371(.a(_w_630),.q(_w_631));
  bfr _b_398(.a(_w_657),.q(_w_658));
  bfr _b_372(.a(_w_631),.q(n190_4));
  bfr _b_377(.a(_w_636),.q(_w_637));
  and_bb g251(.a(n239_1),.b(n250_0),.q(n251));
  spl2 g151_s_2(.a(n151_3),.q0(n151_4),.q1(n151_5));
  bfr _b_379(.a(_w_638),.q(_w_639));
  bfr _b_380(.a(_w_639),.q(_w_640));
  bfr _b_381(.a(_w_640),.q(_w_641));
  bfr _b_383(.a(_w_642),.q(_w_643));
  or_bb g138(.a(in_56_),.b(in_57_),.q(n138));
  bfr _b_518(.a(_w_777),.q(_w_778));
  bfr _b_385(.a(_w_644),.q(_w_645));
  bfr _b_388(.a(_w_647),.q(_w_648));
  bfr _b_390(.a(_w_649),.q(_w_650));
  bfr _b_391(.a(_w_650),.q(_w_651));
  spl2 g150_s_0(.a(n150),.q0(n150_0),.q1(n150_1));
  bfr _b_395(.a(_w_654),.q(n65));
  bfr _b_493(.a(_w_752),.q(_w_753));
  bfr _b_396(.a(_w_655),.q(n145));
  maj_bbi g188(.a(n142_4),.b(n187),.c(n186_0),.q(n188));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  bfr _b_397(.a(_w_656),.q(n140));
  bfr _b_399(.a(_w_658),.q(_w_659));
  spl3L g197_s_0(.a(n197),.q0(n197_0),.q1(n197_1),.q2(n197_2));
  bfr _b_516(.a(_w_775),.q(_w_776));
  bfr _b_400(.a(_w_659),.q(n133_1));
  bfr _b_409(.a(_w_668),.q(_w_669));
  bfr _b_542(.a(_w_801),.q(_w_802));
  bfr _b_410(.a(_w_669),.q(_w_670));
  bfr _b_505(.a(_w_764),.q(n97));
  bfr _b_378(.a(_w_637),.q(n136_2));
  bfr _b_415(.a(_w_674),.q(n126));
  bfr _b_418(.a(_w_677),.q(_w_678));
  bfr _b_367(.a(_w_626),.q(_w_627));
  bfr _b_421(.a(_w_680),.q(n123));
  or_bb g145(.a(n128_0),.b(n144_0),.q(_w_655));
  spl2 g144_s_0(.a(n144),.q0(n144_0),.q1(n144_1));
  bfr _b_497(.a(_w_756),.q(_w_757));
  bfr _b_422(.a(_w_681),.q(n134));
  bfr _b_424(.a(_w_683),.q(n91));
  bfr _b_539(.a(_w_798),.q(_w_799));
  maj_bbi g135(.a(n130_2),.b(n134),.c(n133_0),.q(n135));
  bfr _b_426(.a(_w_685),.q(_w_686));
  maj_bbi g181(.a(n122_4),.b(n180),.c(n179_0),.q(n181));
  bfr _b_428(.a(_w_687),.q(n86));
  maj_bbi g114(.a(n111_1),.b(n112_1),.c(n110_1),.q(_w_712));
  bfr _b_432(.a(_w_691),.q(n109));
  and_bb g132(.a(in_50_),.b(in_51_),.q(n132));
  bfr _b_394(.a(_w_653),.q(_w_654));
  bfr _b_478(.a(_w_737),.q(n120));
  bfr _b_434(.a(_w_693),.q(n83));
  bfr _b_435(.a(_w_694),.q(n80));
  spl3L g189_s_0(.a(n189),.q0(n189_0),.q1(n189_1),.q2(n189_2));
  bfr _b_436(.a(_w_695),.q(_w_696));
  maj_bbi g156(.a(n155),.b(n79_4),.c(n154_0),.q(n156));
  bfr _b_446(.a(_w_705),.q(_w_706));
  bfr _b_447(.a(_w_706),.q(_w_707));
  bfr _b_448(.a(_w_707),.q(n66));
  bfr _b_401(.a(_w_660),.q(n103));
  bfr _b_528(.a(_w_787),.q(_w_788));
  bfr _b_450(.a(_w_709),.q(n93_2));
  bfr _b_454(.a(_w_713),.q(n198));
  bfr _b_455(.a(_w_714),.q(n77));
  bfr _b_464(.a(_w_723),.q(_w_724));
  bfr _b_457(.a(_w_716),.q(_w_717));
  bfr _b_463(.a(_w_722),.q(n154_1));
  spl2 g190_s_0(.a(n190),.q0(n190_0),.q1(n190_1));
  bfr _b_465(.a(_w_724),.q(_w_725));
  bfr _b_467(.a(_w_726),.q(_w_727));
  bfr _b_504(.a(_w_763),.q(n90_3));
  bfr _b_468(.a(_w_727),.q(n86_2));
  bfr _b_404(.a(_w_663),.q(_w_664));
  bfr _b_469(.a(_w_728),.q(_w_729));
  bfr _b_470(.a(_w_729),.q(_w_730));
  bfr _b_473(.a(_w_732),.q(_w_733));
  bfr _b_476(.a(_w_735),.q(n108));
  bfr _b_477(.a(_w_736),.q(n166));
  or_bb g149(.a(n127_1),.b(n147_1),.q(_w_715));
  bfr _b_445(.a(_w_704),.q(_w_705));
  bfr _b_480(.a(_w_739),.q(n70_3));
  bfr _b_513(.a(_w_772),.q(_w_773));
  bfr _b_481(.a(_w_740),.q(n196));
  bfr _b_392(.a(_w_651),.q(_w_652));
  bfr _b_482(.a(_w_741),.q(n139_3));
  bfr _b_353(.a(_w_612),.q(_w_613));
  spl3L g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1),.q2(n172_2));
  bfr _b_483(.a(_w_742),.q(_w_743));
  bfr _b_484(.a(_w_743),.q(_w_744));
  bfr _b_485(.a(_w_744),.q(n161_1));
  spl3L g158_s_1(.a(n158_1),.q0(n158_2),.q1(n158_3),.q2(_w_745));
  bfr _b_486(.a(_w_745),.q(_w_746));
  bfr _b_366(.a(_w_625),.q(n175_1));
  bfr _b_488(.a(_w_747),.q(n158_4));
  bfr _b_514(.a(_w_773),.q(n113_1));
  bfr _b_489(.a(_w_748),.q(_w_749));
  bfr _b_490(.a(_w_749),.q(_w_750));
  bfr _b_494(.a(_w_753),.q(out_4_));
  bfr _b_402(.a(_w_661),.q(n152));
  bfr _b_495(.a(_w_754),.q(n119_3));
  bfr _b_499(.a(_w_758),.q(n179_1));
  bfr _b_510(.a(_w_769),.q(_w_770));
  and_bb g93(.a(in_26_),.b(in_27_),.q(n93));
  bfr _b_508(.a(_w_767),.q(n76_1));
  bfr _b_414(.a(_w_673),.q(n128));
  bfr _b_511(.a(_w_770),.q(n119_1));
  bfr _b_517(.a(_w_776),.q(n105_2));
  bfr _b_519(.a(_w_778),.q(_w_779));
  bfr _b_520(.a(_w_779),.q(n186_1));
  bfr _b_433(.a(_w_692),.q(n143));
  bfr _b_522(.a(_w_781),.q(n87_2));
  bfr _b_523(.a(_w_782),.q(_w_783));
  bfr _b_524(.a(_w_783),.q(_w_784));
  bfr _b_526(.a(_w_785),.q(_w_786));
  bfr _b_530(.a(_w_789),.q(n85));
  bfr _b_532(.a(_w_791),.q(n116_2));
  bfr _b_534(.a(_w_793),.q(n73_2));
  or_bb g191(.a(n186_3),.b(n189_2),.q(_w_738));
  and_bb g182(.a(n125_1),.b(n181_0),.q(n182));
  bfr _b_535(.a(_w_794),.q(n76_3));
  maj_bbi g97(.a(n94_1),.b(n95_1),.c(n93_1),.q(_w_764));
  bfr _b_536(.a(_w_795),.q(_w_796));
  bfr _b_537(.a(_w_796),.q(_w_797));
  bfr _b_538(.a(_w_797),.q(n70_1));
  assign out_0_ = 1'b0;
endmodule
