module c880 (N1,N101,N106,N111,N116,N121,N126,N13,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N17,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N26,N260,N261,N267,N268,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N8,N80,N85,N86,N87,N88,N89,N90,N91,N96,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880);
  input N1,N101,N106,N111,N116,N121,N126,N13,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N17,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N26,N260,N261,N267,N268,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N8,N80,N85,N86,N87,N88,N89,N90,N91,N96;
  output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880;
  wire _w_2172,_w_2171,_w_2168,_w_2167,_w_2166,_w_2161,_w_2158,_w_2156,_w_2147,_w_2146,_w_2145,_w_2140,_w_2135,_w_2133,_w_2131,_w_2125,_w_2124,_w_2121,_w_2120,_w_2115,_w_2111,_w_2109,_w_2105,_w_2103,_w_2101,_w_2100,_w_2099,_w_2096,_w_2095,_w_2094,_w_2092,_w_2090,_w_2088,_w_2086,_w_2084,_w_2162,_w_2083,_w_2080,_w_2173,_w_2106,_w_2078,_w_2073,_w_2072,_w_2071,_w_2070,_w_2067,_w_2066,_w_2054,_w_2050,_w_2049,_w_2043,_w_2042,_w_2041,_w_2039,_w_2036,_w_2033,_w_2031,_w_2028,_w_2026,_w_2024,_w_2020,_w_2016,_w_2015,_w_2014,_w_2013,_w_2009,_w_2008,_w_2007,_w_2006,_w_2005,_w_2004,_w_2000,_w_1999,_w_1996,_w_1994,_w_1993,_w_1991,_w_1989,_w_1986,_w_1983,_w_1981,_w_1980,_w_1975,_w_1973,_w_1972,_w_1967,_w_1964,_w_1960,_w_1959,_w_1958,_w_1957,_w_1954,_w_1952,_w_1951,_w_1948,_w_1946,_w_1945,_w_1941,_w_1940,_w_1971,_w_1939,_w_1936,_w_1935,_w_1934,_w_1933,_w_1925,_w_1924,_w_1923,_w_1921,_w_1916,_w_1915,_w_1913,_w_1912,_w_1909,_w_2089,_w_1906,_w_1904,_w_1903,_w_1902,_w_1899,_w_1898,_w_1897,_w_1895,_w_1886,_w_1885,_w_1882,_w_1881,_w_1879,_w_1877,_w_1875,_w_1874,_w_1872,_w_1920,_w_1870,_w_1869,_w_2142,_w_1867,_w_1865,_w_2068,_w_1862,_w_1861,_w_1860,_w_1859,_w_1856,_w_1851,_w_1850,_w_1849,_w_2055,_w_1848,_w_1846,_w_1844,_w_1842,_w_1840,_w_1839,_w_1838,_w_1836,_w_1828,_w_1827,_w_1826,_w_1825,_w_1823,_w_1820,_w_1819,_w_1818,_w_1816,_w_1810,_w_1805,_w_1835,_w_1803,_w_1802,_w_1799,_w_1794,_w_1793,_w_1792,_w_1791,_w_1789,_w_1787,_w_1785,_w_1873,_w_1853,_w_1784,_w_1781,_w_1780,_w_1779,_w_2069,_w_1777,_w_1776,_w_1775,_w_1772,_w_1771,_w_1770,_w_2087,_w_1768,_w_1766,_w_1765,_w_1764,_w_1763,_w_1762,_w_1760,_w_1759,_w_1758,_w_1757,_w_1756,_w_1876,_w_1755,_w_1752,_w_1749,_w_1747,_w_1963,_w_1745,_w_1744,_w_1738,_w_1737,_w_1893,_w_1733,_w_1731,_w_1938,_w_1726,_w_1724,_w_1722,_w_1721,_w_1720,_w_1719,_w_1718,_w_1717,_w_1716,_w_1710,_w_1707,_w_2107,_w_1704,_w_1701,_w_1700,_w_1698,_w_1696,_w_1695,_w_2129,_w_1694,_w_2023,_w_1691,_w_1686,_w_1685,_w_1684,_w_1681,_w_1680,_w_1675,_w_1673,_w_1668,_w_1666,_w_2012,_w_1665,_w_1660,_w_1814,_w_1658,_w_1657,_w_1655,_w_2134,_w_2119,_w_1654,_w_1653,_w_1652,_w_1651,_w_1650,_w_1647,_w_1644,_w_1643,_w_1642,_w_2038,_w_1639,_w_1832,_w_1638,_w_1634,_w_2082,_w_1630,_w_1623,_w_1622,_w_2017,_w_1621,_w_1997,_w_1612,_w_1611,_w_1627,_w_1610,_w_1609,_w_1607,_w_1606,_w_1605,_w_1603,_w_1599,_w_1597,_w_1595,_w_1592,_w_1590,_w_1589,_w_1976,_w_1588,_w_1927,_w_1587,_w_1833,_w_1584,_w_1583,_w_1582,_w_1581,_w_2037,_w_1579,_w_1837,_w_1576,_w_1575,_w_1574,_w_1572,_w_1570,_w_1568,_w_1567,_w_1565,_w_1562,_w_1561,_w_2058,_w_1559,_w_1558,_w_1557,_w_1556,_w_1552,_w_1550,_w_1543,_w_2170,_w_1542,_w_1541,_w_1538,_w_1555,_w_1537,_w_1536,_w_1535,_w_1544,_w_1533,_w_1532,_w_1528,_w_2021,_w_1693,_w_1560,_w_1527,_w_1831,_w_1522,_w_1520,_w_1518,_w_1513,_w_1640,_w_1512,_w_2085,_w_1511,_w_1510,_w_1507,_w_1505,_w_1504,_w_1502,_w_1499,_w_1495,_w_1761,_w_1493,_w_1491,_w_1490,_w_1806,_w_1486,_w_1484,_w_1482,_w_1481,_w_1809,_w_1479,_w_1476,_w_1474,_w_1472,_w_1470,_w_1467,_w_1600,_w_1466,_w_1930,_w_1628,_w_1465,_w_1463,_w_2076,_w_1460,_w_1457,_w_1456,_w_1821,_w_1453,_w_1451,_w_1448,_w_1447,_w_1446,_w_1444,_w_1855,_w_1443,_w_1442,_w_1441,_w_2077,_w_2061,_w_1440,_w_1439,_w_1648,_w_1438,_w_1434,_w_1427,_w_1425,_w_1424,_w_1667,_w_1422,_w_1421,_w_1496,_w_1420,_w_1415,_w_1414,_w_1413,_w_1754,_w_1732,_w_1437,_w_1412,_w_1868,_w_1410,_w_1406,_w_1402,_w_1401,_w_1400,_w_1399,_w_1398,_w_2108,_w_1394,_w_1616,_w_1392,_w_1995,_w_1515,_w_1391,_w_1390,_w_1388,_w_1387,_w_1384,_w_1383,_w_1382,_w_1547,_w_1381,_w_1564,_w_1380,_w_1379,_w_2027,_w_1378,_w_1678,_w_1376,_w_1375,_w_1373,_w_1371,_w_1369,_w_1713,_w_1368,_w_1365,_w_1364,_w_1950,_w_1362,_w_1360,_w_2001,_w_1358,_w_1356,_w_1355,_w_1677,_w_1353,_w_1351,_w_1350,_w_1348,_w_1345,_w_2010,_w_1342,_w_1430,_w_1339,_w_2059,_w_1807,_w_1337,_w_1334,_w_1598,_w_1344,_w_1333,_w_2152,_w_1332,_w_1330,_w_2153,_w_1699,_w_1329,_w_1323,_w_2112,_w_1322,_w_1321,_w_2136,_w_2132,_w_1320,_w_1319,_w_1937,_w_1315,_w_1314,_w_1312,_w_1311,_w_1813,_w_1540,_w_1309,_w_1308,_w_2141,_w_1307,_w_2169,_w_1306,_w_2045,_w_1303,_w_1301,_w_1300,_w_1297,_w_1296,_w_1689,_w_1294,_w_1293,_w_1292,_w_1291,_w_1289,_w_1546,_w_1287,_w_1521,_w_1286,_w_1349,_w_1284,_w_1283,_w_1282,_w_1619,_w_1281,_w_1955,_w_1280,_w_1279,_w_1277,_w_1276,_w_1275,_w_1662,_w_1273,_w_1272,_w_1485,_w_1270,_w_1468,_w_1267,_w_1264,_w_1263,_w_1261,_w_1259,_w_1847,_w_1258,_w_1688,_w_1257,_w_1256,_w_1255,_w_1253,_w_1636,_w_1252,_w_1459,_w_1251,_w_1250,_w_1340,_w_1249,_w_1248,_w_1594,_w_1245,_w_1242,_w_1241,_w_1238,_w_1237,_w_1596,_w_1233,_w_1232,_w_1230,_w_1372,_w_1223,_w_1222,_w_1428,_w_1221,_w_1409,_w_1243,_w_1220,_w_1480,_w_1217,_w_1900,_w_1735,_w_1215,_w_1214,_w_1213,_w_1211,_w_1210,_w_1208,_w_1206,_w_1204,_w_2159,_w_1203,_w_1200,_w_1199,_w_1197,_w_2062,_w_1585,_w_1194,_w_1928,_w_1730,_w_1193,_w_1191,_w_1190,_w_1817,_w_1187,_w_1186,_w_1432,_w_1184,_w_1219,_w_1183,_w_2104,_w_1182,_w_1632,_w_1181,_w_1179,_w_1176,_w_1175,_w_1174,_w_1173,_w_1171,_w_1901,_w_1767,_w_1509,_w_1169,_w_1664,_w_1166,_w_1396,_w_1163,_w_1162,_w_1159,_w_1483,_w_1158,_w_2052,_w_1157,_w_1156,_w_2138,_w_1246,_w_1155,_w_1153,_w_2144,_w_1152,_w_2046,_w_1949,_w_1150,_w_1646,_w_1149,_w_1617,_w_1146,_w_1144,_w_1890,_w_1141,_w_1138,_w_1137,_w_1134,_w_1133,_w_1132,_w_1131,_w_1129,_w_1127,_w_1126,_w_1122,_w_1120,_w_2003,_w_1753,_w_1119,_w_1118,_w_1117,_w_1216,_w_1115,_w_1114,_w_1961,_w_1435,_w_1113,_w_1112,_w_1111,_w_1464,n145_0,_w_2025,N55_2,N255_1,N268_3,_w_1477,_w_953,_w_1012,_w_1054,n92_1,_w_1235,n92_0,_w_1161,N59_1,_w_886,N59_0,_w_1626,N390_1,n302_0,_w_1450,n253,N390_0,_w_1445,_w_1423,n286_1,N17_5,_w_1539,n162_1,_w_845,N17_3,_w_2149,_w_1586,n263_0,N17_2,_w_1052,_w_1649,N17_0,_w_1894,_w_1475,_w_1417,N80_2,_w_2128,_w_864,_w_1452,n75_0,n95_0,N42_7,_w_871,_w_1703,N42_1,N42_6,_w_1709,_w_1271,N42_0,_w_1907,N130_3,_w_2164,_w_909,N106_1,N91_0,_w_1635,n296,N96_1,_w_1979,n162_3,_w_1808,n322_1,N447_1,N153_1,_w_1290,N153_0,_w_2150,n153,_w_1645,_w_1563,N68_0,_w_1288,n70_1,n270_3,n270_2,n191,_w_1748,_w_1262,n270_1,n270_0,n198_1,n73_0,n122,_w_1687,N135_1,_w_2130,_w_962,n199_2,_w_1525,n210,n110_1,_w_1679,_w_1067,n113_1,_w_1822,n235,_w_1436,n286_3,_w_1433,N101_3,n67,_w_1674,N101_1,N101_0,n263_3,n194_0,_w_925,n263_1,N17_8,_w_844,_w_2102,N42_9,n350,_w_1299,_w_889,n144,_w_1982,N13_0,n278_1,_w_1571,n202_1,_w_2139,_w_1285,n279_1,_w_861,_w_1501,n294_3,_w_2040,_w_1019,N42_5,_w_2093,_w_1812,_w_1712,n294_2,n199_1,_w_1843,n294_1,n296_1,n338,N29_2,_w_1489,N171_1,n298_0,n304_2,n281,_w_1942,_w_1473,n304_1,N237_1,n61,_w_884,_w_1317,_w_968,n337_0,_w_1519,n61_1,n364,_w_1910,_w_1201,n363,n138,n359,n207,n271_2,N219_1,n356,n355,n248,_w_1578,n349,n348,N51_0,N91_3,n345,n206_1,n343,N126_0,_w_1854,n166_1,_w_1620,_w_1045,n340,_w_954,n339,_w_1244,n162_0,n68_0,n342,n272_1,n337,n335,n334,n280_0,n151,n331,_w_1488,n330,_w_1931,n186,N189_3,_w_1947,_w_1366,n198_0,_w_902,n329,N68_1,n152_0,n328,_w_1096,n110_0,n83_1,n134_0,n325,_w_1164,n323,n320,n165_2,n319,n302_1,_w_2081,n358,_w_1830,n316,N13_1,_w_1637,_w_975,n312,_w_1154,n310,n239,_w_1188,_w_1092,n308,_w_1659,n142,_w_1260,n305,_w_1361,_w_989,n304,n199,N149_0,n341,n193_0,n301,_w_1711,N219_14,_w_1225,_w_969,n300,_w_1984,_w_1888,n303,n109,_w_1811,N210_4,_w_2047,_w_1487,_w_1236,n297,_w_2091,_w_1553,_w_1010,_w_1354,n337_1,N447_2,n289,n271_1,n128_1,n284,_w_2079,n226,n282,n277,n324,_w_1723,n302,n182,n147_3,n233,_w_1663,_w_1109,_w_908,_w_976,_w_1148,n276,_w_1254,n162_2,n272,_w_963,_w_994,_w_1714,n266,_w_1346,N29_0,n279_0,N447_0,n317,n262,_w_1834,n259,_w_978,_w_1227,_w_998,_w_1226,N17_6,n258,n300_1,_w_1234,n256,N165_1,_w_1123,_w_912,_w_1099,n254,_w_1769,n197,n124,n286,n228_1,_w_1896,_w_1192,n113,n106,n90,n111,_w_1953,n63_0,_w_1965,n228_0,_w_1001,n78_0,n150_1,n187,n249,_w_1205,_w_1198,n128,n192,_w_1304,n211,_w_2116,n103,n234,_w_1228,N447_3,n102,_w_2011,N59_2,_w_1708,_w_1269,n315,_w_1177,N143_0,n162_5,N261_1,_w_2057,n292,n194_1,n215,_w_1966,_w_1697,_w_875,n87,n195,n68,N42_3,n78,_w_1824,n347,n270,n294,n218,n332,_w_1015,n117,n94,_w_1128,n295,_w_841,_w_1032,n271,n133,_w_1871,N121_1,N210_0,_w_887,_w_1503,_w_1011,N80_3,n162_9,n174,_w_1741,n184,n293,n223,_w_1683,_w_1526,n154,n178,_w_1506,n278_3,n318,n288_0,_w_1740,_w_1079,n280,n322,N159_0,n162,_w_1841,n271_0,_w_1892,n183,n162_4,_w_1727,_w_894,n283,n268,_w_1367,n286_0,n130,_w_2163,n365,_w_952,_w_1101,_w_1864,_w_1151,N135_0,_w_1462,n245,n98_0,n247,_w_1548,n287_1,_w_1325,_w_847,_w_1970,n337_2,n93,n163,_w_862,n75,_w_1566,n131,n172,n300_2,n205,_w_2051,n131_1,N171_2,N75_1,n83_0,n307_1,n220,_w_1778,_w_965,_w_1706,N42_4,_w_1577,n228,N228_11,n229,_w_1110,_w_1458,_w_2053,N51_3,_w_2063,N171_6,n279_2,n83,n322_2,n150_0,n209,_w_1416,n285,_w_1023,_w_1601,n266_2,_w_2056,_w_1028,_w_1140,N201_1,n61_0,n278,_w_851,N91_4,_w_1880,_w_997,n112,N237_4,_w_2030,N219_2,N219_10,n147,n145,_w_921,_w_1884,n313,_w_1105,n265,_w_1108,n302_2,n113_0,n162_8,_w_1072,_w_1060,n167,_w_1266,n255,_w_1656,_w_1419,_w_1998,n101,n327,N29_1,n216,n136,_w_1676,_w_1407,_w_939,n73_1,n96,_w_1911,_w_1786,_w_984,N228_3,n278_2,n280_1,_w_2113,n134_1,N80_1,N80_4,_w_1029,N228_7,N246_3,_w_2118,_w_1914,_w_1863,_w_982,n160,_w_1932,n91,n298_1,n169,n128_0,_w_1104,_w_1545,n360,n155,n180,_w_1887,_w_1829,_w_2154,_w_1049,_w_1310,_w_1318,N165_0,N177_1,n179_5,n257,_w_1492,n311,_w_950,N268_0,n110,n333,n120,_w_1790,n147_0,_w_1962,n352,n161,_w_1038,_w_1085,n125,n196,_w_2126,n132,n129,n263_2,_w_867,_w_1147,n86_1,N17_4,_w_1524,n213_0,_w_852,_w_942,N246_10,_w_1551,n86_0,N237_8,n175,N165_3,_w_1357,n298,N143_1,n118,_w_1514,n107_0,n267,_w_1395,_w_857,n168,n344,n78_1,n326,_w_957,_w_1265,n204,_w_1728,n137,n199_0,N268_2,n100,_w_1027,_w_1135,n139,n211_0,n288,n158,_w_993,n144_0,n84,_w_1328,_w_834,n240,N96_0,n238,N189_5,_w_1671,n300_0,_w_1338,n140,n104,N96_2,n148,_w_1783,n179_2,_w_1591,_w_1508,n202,_w_896,n125_0,_w_899,_w_1359,n149,n123,_w_1374,n98_1,N390_2,N210_6,_w_1750,n266_0,n168_1,_w_1397,n152,n67_2,_w_1593,n278_0,_w_2123,n322_0,n309,N228_9,n314,n97,_w_831,_w_1580,n156,_w_1631,_w_1142,_w_1077,_w_1078,n157,_w_1385,n193,n162_7,n217,N101_2,n179_1,n228_2,_w_1549,n274,n83_2,_w_2148,_w_1268,n214,_w_1682,_w_1084,_w_1969,n194,_w_1316,N268_1,n164,n298_2,n210_1,_w_936,_w_1889,n165,_w_2160,n213_2,n166,n170,_w_1302,n206_0,n98,_w_1313,n354,n171,_w_1449,n287,_w_1065,n176,_w_2155,n82,N237_13,_w_1426,n177,N210_1,_w_1036,n179,_w_1705,_w_1454,_w_1370,N80_0,_w_1618,_w_859,_w_1178,n181,n304_0,_w_2065,_w_1944,n189,_w_2060,_w_1883,N91_2,_w_907,n70,_w_935,n208,n296_0,n202_0,_w_916,N261_2,n200,_w_1404,_w_972,n159,n75_1,n99,_w_1389,_w_1005,n203,_w_1615,_w_1107,n115,_w_973,n353,N17_1,n212,_w_1343,n213,N201_3,_w_1604,n295_0,N261_0,n204_0,n219,n162_6,n221,N101_4,N51_1,_w_2034,n225,N106_2,n134,_w_1641,N91_1,_w_1523,n230,n237,N177_6,N17_10,n86,n291,_w_1554,n246,N121_2,_w_1331,n202_2,n105,n68_1,n213_1,_w_1742,N96_3,_w_1098,_w_1008,n198,n362,_w_1327,N219_7,_w_890,n146,_w_1573,n294_0,_w_1725,_w_836,n242,n243,N1_2,_w_1074,n286_2,_w_1239,n70_0,N17_9,n71,n251,N55_1,N36_0,_w_1529,_w_854,N36_1,_w_1905,n250,N237_0,_w_1195,N29_3,n71_1,N237_2,N237_3,_w_1168,_w_835,_w_850,N237_5,_w_1773,_w_1729,N237_6,_w_1530,n352_0,_w_1091,_w_1990,_w_1025,n263,N237_7,_w_2019,_w_1804,_w_905,_w_1968,N237_9,_w_1405,N237_12,_w_1167,n167_0,_w_1231,n167_1,N111_1,_w_1471,n167_2,N219_3,N210_5,N219_5,N219_6,_w_2029,_w_1121,N219_8,_w_1469,N219_11,N42_10,_w_911,N219_12,_w_1613,N55_0,N207_0,N207_1,n101_0,N159_2,_w_1295,n101_1,N189_0,_w_1497,N189_1,N189_2,_w_1977,N189_4,_w_999,N189_6,n190,n67_0,_w_1037,N228_12,n67_1,_w_1305,n119_0,N183_1,_w_1003,n260,_w_1090,_w_1139,N183_2,N183_3,_w_943,_w_1224,N237_11,N183_4,_w_1788,_w_1143,N138_1,_w_2122,_w_1891,n114,N183_5,n236,N183_6,_w_858,N177_0,_w_855,_w_2002,N177_2,_w_2032,N177_4,_w_981,n224,N177_5,N159_5,N1_0,_w_1908,N1_1,N8_0,_w_1478,N8_1,_w_863,N165_2,N165_4,N255_0,_w_898,N165_5,_w_900,n272_0,N177_3,N165_6,_w_1569,n193_2,N121_0,N121_3,n192_0,_w_1661,_w_1429,_w_1298,n192_1,_w_1782,N210_7,n192_2,_w_958,n192_3,N138_0,_w_2151,_w_1743,N138_3,N130_0,N130_2,_w_1858,N130_4,_w_1715,_w_1070,N126_1,N126_2,n71_0,N149_1,n201,n287_0,_w_1629,N246_1,_w_1866,_w_1608,_w_1063,n287_2,N75_0,_w_2064,N111_0,_w_1013,N195_2,_w_922,N111_2,n198_2,_w_879,N111_3,_w_1240,_w_948,N106_0,_w_1278,_w_1172,_w_1071,N106_3,_w_1494,N106_4,_w_1531,_w_960,_w_1534,n288_1,N116_0,_w_881,N116_1,_w_838,n144_1,_w_1076,_w_1988,N116_2,N42_2,n141,N116_3,n119_1,_w_2127,_w_1702,_w_1018,N159_1,_w_949,N159_3,_w_1774,N219_13,N159_6,N171_0,n122_0,n122_1,_w_1196,n352_2,_w_1247,n125_1,_w_1625,n140_1,_w_874,_w_1006,_w_1633,N228_0,_w_873,N228_1,_w_1795,N228_2,_w_865,N228_4,n279,_w_986,N228_5,_w_2137,_w_1180,N228_6,_w_938,n206,_w_1094,_w_1919,N228_8,n137_0,_w_934,N228_10,n266_3,_w_1087,_w_2022,_w_1363,n168_0,N201_6,n135,n168_2,n204_1,n204_2,n241,n179_3,N138_2,_w_914,n137_1,_w_2075,N146_0,n140_0,n104_0,_w_928,n104_1,_w_2110,_w_1064,_w_1106,n147_1,_w_1922,_w_1878,_w_1136,n63_1,n152_1,n173,n131_0,n152_2,_w_1069,_w_1797,n152_3,n152_4,N171_3,_w_1845,n95_1,N171_4,N51_2,n107,_w_961,_w_1624,n165_0,_w_1670,n165_1,n166_0,_w_951,_w_945,N17_7,N210_3,_w_1614,N210_8,N210_9,n210_0,n210_2,n206_2,n210_3,n92,n179_0,n179_4,n179_7,_w_1987,N246_0,n179_8,_w_1341,n273,n307_0,_w_1145,n361,N201_0,N201_2,N201_4,N195_0,N201_5,n200_0,n200_1,_w_1498,_w_1103,n179_6,N195_1,n211_1,_w_1100,_w_1796,_w_1274,_w_995,N228_13,N195_4,N42_8,_w_1022,_w_2165,_w_1229,N195_5,_w_2074,N195_6,_w_1335,n211_2,_w_1326,_w_1189,n185,_w_1042,n212_0,_w_2098,n252,n212_1,N246_2,N246_4,N219_9,N246_5,_w_1734,_w_1352,_w_1202,n352_1,N246_6,_w_1943,N96_4,n232,N246_7,N246_8,N246_9,_w_2048,_w_1801,n295_1,N138_4,_w_918,n107_1,_w_1672,n245_0,_w_1455,_w_946,n245_1,_w_1130,n346,n245_2,_w_833,_w_1800,_w_837,_w_839,N183_0,_w_840,_w_1461,n307,_w_1000,_w_842,_w_1602,_w_843,_w_1418,_w_846,_w_1431,_w_848,_w_849,_w_944,_w_1377,_w_853,_w_856,_w_860,_w_868,_w_1393,_w_869,_w_1209,_w_872,_w_870,_w_876,_w_1852,_w_931,_w_1170,_w_1044,_w_866,_w_877,_w_1669,_w_878,_w_880,_w_1075,N171_5,_w_882,_w_883,_w_885,_w_888,_w_891,n299,_w_832,_w_892,_w_893,_w_895,_w_897,n150,_w_901,_w_990,n295_2,_w_903,n73,_w_904,_w_1956,_w_1929,_w_906,_w_910,_w_1857,_w_1082,_w_1918,n290,_w_913,_w_1324,_w_915,_w_2117,N237_10,N130_1,N55_3,_w_917,_w_919,_w_1974,_w_1386,N146_1,_w_920,_w_1009,n147_2,_w_923,_w_1124,_w_924,n266_1,_w_926,_w_927,n357,_w_929,_w_2018,_w_930,n119,_w_932,_w_933,n127,_w_937,n126,_w_940,_w_941,_w_947,N219_4,_w_955,_w_956,_w_1056,_w_1212,_w_959,_w_2035,_w_964,_w_966,_w_967,_w_1411,_w_970,_w_1690,_w_971,_w_1093,_w_1815,_w_1403,_w_1207,_w_974,_w_1517,_w_1408,N219_0,n63,_w_977,_w_1125,_w_979,_w_980,_w_2044,_w_983,_w_985,_w_1160,_w_1024,N210_2,_w_987,_w_988,_w_1917,_w_991,_w_992,_w_996,_w_1739,_w_1002,_w_1004,_w_1692,_w_1500,_w_1007,n231,_w_1014,_w_1751,_w_1165,_w_1016,_w_1798,_w_1516,_w_1017,_w_1336,_w_1020,_w_2114,_w_1021,_w_1026,_w_1030,_w_1736,_w_1347,_w_1031,n264,_w_1040,n269,_w_1033,_w_1978,_w_1746,n222,_w_1034,_w_1035,N255_2,_w_1039,N59_3,_w_1041,_w_1043,_w_1046,_w_1047,_w_1992,_w_1048,_w_1116,N195_3,_w_1050,n179_9,_w_1051,_w_2157,n145_1,N261_3,_w_1053,n198_3,_w_1055,_w_1185,_w_1057,_w_1985,n275,_w_1058,n193_1,_w_1059,_w_1061,n108,_w_1062,_w_1066,_w_1068,_w_1926,_w_1073,_w_1080,_w_2143,_w_1081,_w_1218,_w_1083,n95,_w_1086,_w_1088,_w_2097,_w_1089,_w_1095,n121,_w_1097,N159_4,_w_1102;

  bfr _b_1837(.a(_w_2169),.q(_w_2170));
  bfr _b_1836(.a(_w_2168),.q(_w_2169));
  bfr _b_1832(.a(_w_2164),.q(_w_2163));
  bfr _b_1831(.a(N90),.q(_w_2164));
  bfr _b_1829(.a(N89),.q(_w_2162));
  bfr _b_1827(.a(_w_2159),.q(_w_2160));
  bfr _b_1825(.a(_w_2157),.q(_w_2155));
  bfr _b_1824(.a(_w_2156),.q(_w_2157));
  bfr _b_1823(.a(N74),.q(_w_2156));
  bfr _b_1821(.a(N73),.q(_w_2154));
  bfr _b_1814(.a(N268),.q(_w_2147));
  bfr _b_1813(.a(N267),.q(_w_2145));
  bfr _b_1812(.a(_w_2144),.q(_w_2131));
  bfr _b_1808(.a(_w_2140),.q(_w_2141));
  bfr _b_1807(.a(_w_2139),.q(_w_2140));
  bfr _b_1805(.a(_w_2137),.q(_w_2138));
  bfr _b_1804(.a(_w_2136),.q(_w_2137));
  bfr _b_1799(.a(N261),.q(_w_2132));
  bfr _b_1796(.a(N259),.q(_w_2128));
  bfr _b_1794(.a(_w_2126),.q(_w_2127));
  bfr _b_1793(.a(_w_2125),.q(_w_2126));
  bfr _b_1792(.a(_w_2124),.q(_w_2125));
  bfr _b_1789(.a(_w_2121),.q(_w_2122));
  bfr _b_1788(.a(_w_2120),.q(_w_2121));
  bfr _b_1787(.a(_w_2119),.q(_w_2120));
  bfr _b_1786(.a(_w_2118),.q(_w_2119));
  bfr _b_1783(.a(_w_2115),.q(_w_2116));
  bfr _b_1781(.a(_w_2113),.q(_w_2114));
  bfr _b_1777(.a(_w_2109),.q(_w_2110));
  bfr _b_1774(.a(_w_2106),.q(_w_2107));
  bfr _b_1769(.a(_w_2101),.q(_w_2102));
  bfr _b_1768(.a(_w_2100),.q(_w_2101));
  bfr _b_1767(.a(_w_2099),.q(_w_2100));
  bfr _b_1765(.a(_w_2097),.q(_w_2098));
  bfr _b_1763(.a(_w_2095),.q(_w_2096));
  bfr _b_1758(.a(_w_2090),.q(_w_2091));
  bfr _b_1754(.a(_w_2086),.q(_w_2070));
  bfr _b_1752(.a(_w_2084),.q(_w_2085));
  bfr _b_1750(.a(_w_2082),.q(_w_2083));
  bfr _b_1749(.a(_w_2081),.q(_w_2082));
  bfr _b_1748(.a(_w_2080),.q(_w_2081));
  bfr _b_1747(.a(_w_2079),.q(_w_2080));
  bfr _b_1746(.a(_w_2078),.q(_w_2079));
  bfr _b_1745(.a(_w_2077),.q(_w_2078));
  bfr _b_1742(.a(_w_2074),.q(_w_2075));
  bfr _b_1740(.a(_w_2072),.q(_w_2073));
  bfr _b_1736(.a(_w_2068),.q(_w_2069));
  bfr _b_1735(.a(N207),.q(_w_2068));
  bfr _b_1732(.a(N159),.q(_w_2064));
  bfr _b_1730(.a(_w_2062),.q(_w_2055));
  bfr _b_1725(.a(_w_2057),.q(_w_2058));
  bfr _b_1724(.a(_w_2056),.q(_w_2057));
  bfr _b_1723(.a(N153),.q(_w_2056));
  bfr _b_1722(.a(N152),.q(_w_2054));
  bfr _b_1720(.a(_w_2052),.q(_w_2053));
  bfr _b_1717(.a(_w_2049),.q(_w_2050));
  bfr _b_1714(.a(N149),.q(_w_2047));
  bfr _b_1713(.a(_w_2045),.q(_w_2038));
  bfr _b_1711(.a(_w_2043),.q(_w_2044));
  bfr _b_1710(.a(_w_2042),.q(_w_2043));
  bfr _b_1738(.a(N219),.q(_w_2071));
  bfr _b_1708(.a(_w_2040),.q(_w_2041));
  bfr _b_1706(.a(N146),.q(_w_2039));
  bfr _b_1705(.a(_w_2037),.q(_w_2030));
  bfr _b_1703(.a(_w_2035),.q(_w_2036));
  bfr _b_1702(.a(_w_2034),.q(_w_2035));
  bfr _b_1701(.a(_w_2033),.q(_w_2034));
  bfr _b_1761(.a(_w_2093),.q(_w_2094));
  bfr _b_1698(.a(N143),.q(_w_2031));
  bfr _b_1697(.a(_w_2029),.q(_w_2027));
  bfr _b_1696(.a(_w_2028),.q(_w_2029));
  bfr _b_1694(.a(N13),.q(_w_2026));
  bfr _b_1692(.a(_w_2024),.q(_w_2025));
  bfr _b_1691(.a(N126),.q(_w_2024));
  bfr _b_1689(.a(_w_2021),.q(_w_2022));
  bfr _b_1688(.a(_w_2020),.q(_w_2021));
  bfr _b_1687(.a(_w_2019),.q(n210_1));
  bfr _b_1686(.a(_w_2018),.q(_w_2019));
  bfr _b_1681(.a(_w_2013),.q(n296));
  bfr _b_1680(.a(_w_2012),.q(_w_2013));
  bfr _b_1679(.a(_w_2011),.q(_w_2012));
  bfr _b_1677(.a(_w_2009),.q(_w_2010));
  bfr _b_1764(.a(_w_2096),.q(_w_2097));
  bfr _b_1675(.a(_w_2007),.q(_w_2008));
  bfr _b_1672(.a(_w_2004),.q(_w_2005));
  bfr _b_1671(.a(_w_2003),.q(_w_2004));
  bfr _b_1666(.a(_w_1998),.q(_w_1999));
  bfr _b_1664(.a(_w_1996),.q(_w_1997));
  bfr _b_1658(.a(_w_1990),.q(_w_1991));
  bfr _b_1657(.a(_w_1989),.q(_w_1990));
  bfr _b_1656(.a(_w_1988),.q(_w_1989));
  bfr _b_1651(.a(_w_1983),.q(_w_1984));
  bfr _b_1649(.a(_w_1981),.q(_w_1982));
  bfr _b_1648(.a(_w_1980),.q(_w_1981));
  bfr _b_1646(.a(_w_1978),.q(N418));
  bfr _b_1641(.a(_w_1973),.q(_w_1974));
  bfr _b_1638(.a(_w_1970),.q(_w_1971));
  bfr _b_1728(.a(_w_2060),.q(_w_2061));
  bfr _b_1634(.a(_w_1966),.q(_w_1967));
  bfr _b_1630(.a(_w_1962),.q(_w_1963));
  bfr _b_1629(.a(_w_1961),.q(_w_1962));
  bfr _b_1628(.a(_w_1960),.q(_w_1961));
  bfr _b_1637(.a(_w_1969),.q(_w_1970));
  bfr _b_1627(.a(_w_1959),.q(_w_1960));
  bfr _b_1625(.a(_w_1957),.q(_w_1958));
  bfr _b_1624(.a(_w_1956),.q(_w_1957));
  bfr _b_1623(.a(_w_1955),.q(_w_1956));
  bfr _b_1621(.a(_w_1953),.q(_w_1954));
  bfr _b_1620(.a(_w_1952),.q(_w_1953));
  bfr _b_1618(.a(_w_1950),.q(_w_1951));
  bfr _b_1614(.a(_w_1946),.q(n280));
  bfr _b_1611(.a(_w_1943),.q(_w_1944));
  bfr _b_1610(.a(_w_1942),.q(_w_1943));
  bfr _b_1609(.a(_w_1941),.q(_w_1942));
  bfr _b_1607(.a(_w_1939),.q(_w_1940));
  bfr _b_1603(.a(_w_1935),.q(_w_1936));
  bfr _b_1600(.a(_w_1932),.q(_w_1933));
  bfr _b_1599(.a(_w_1931),.q(N219_3));
  bfr _b_1596(.a(_w_1928),.q(_w_1929));
  bfr _b_1595(.a(_w_1927),.q(_w_1928));
  bfr _b_1594(.a(_w_1926),.q(_w_1927));
  bfr _b_1593(.a(_w_1925),.q(_w_1926));
  bfr _b_1591(.a(_w_1923),.q(n272));
  bfr _b_1590(.a(_w_1922),.q(_w_1923));
  bfr _b_1773(.a(_w_2105),.q(_w_2106));
  bfr _b_1587(.a(_w_1919),.q(_w_1920));
  bfr _b_1586(.a(_w_1918),.q(_w_1919));
  bfr _b_1584(.a(_w_1916),.q(_w_1917));
  bfr _b_1583(.a(_w_1915),.q(_w_1916));
  bfr _b_1582(.a(_w_1914),.q(_w_1915));
  bfr _b_1580(.a(_w_1912),.q(_w_1913));
  bfr _b_1579(.a(_w_1911),.q(_w_1912));
  bfr _b_1578(.a(_w_1910),.q(_w_1911));
  bfr _b_1577(.a(_w_1909),.q(_w_1910));
  bfr _b_1575(.a(_w_1907),.q(_w_1908));
  bfr _b_1574(.a(_w_1906),.q(_w_1907));
  bfr _b_1573(.a(_w_1905),.q(n271));
  bfr _b_1572(.a(_w_1904),.q(_w_1905));
  bfr _b_1568(.a(_w_1900),.q(_w_1901));
  bfr _b_1567(.a(_w_1899),.q(_w_1900));
  bfr _b_1566(.a(_w_1898),.q(_w_1899));
  bfr _b_1565(.a(_w_1897),.q(_w_1898));
  bfr _b_1563(.a(_w_1895),.q(_w_1896));
  bfr _b_1562(.a(_w_1894),.q(_w_1895));
  bfr _b_1652(.a(_w_1984),.q(_w_1985));
  bfr _b_1560(.a(_w_1892),.q(_w_1893));
  bfr _b_1559(.a(_w_1891),.q(_w_1892));
  bfr _b_1556(.a(_w_1888),.q(_w_1889));
  bfr _b_1555(.a(_w_1887),.q(n267));
  bfr _b_1605(.a(_w_1937),.q(_w_1938));
  bfr _b_1554(.a(_w_1886),.q(_w_1887));
  bfr _b_1841(.a(_w_2173),.q(_w_2171));
  bfr _b_1553(.a(_w_1885),.q(_w_1886));
  bfr _b_1551(.a(_w_1883),.q(_w_1884));
  bfr _b_1550(.a(_w_1882),.q(n260));
  bfr _b_1546(.a(_w_1878),.q(_w_1879));
  bfr _b_1545(.a(_w_1877),.q(_w_1878));
  bfr _b_1633(.a(_w_1965),.q(_w_1966));
  bfr _b_1544(.a(_w_1876),.q(_w_1877));
  bfr _b_1576(.a(_w_1908),.q(_w_1909));
  bfr _b_1542(.a(_w_1874),.q(_w_1875));
  bfr _b_1604(.a(_w_1936),.q(_w_1937));
  bfr _b_1539(.a(_w_1871),.q(_w_1872));
  bfr _b_1690(.a(_w_2022),.q(n199_2));
  bfr _b_1537(.a(_w_1869),.q(_w_1870));
  bfr _b_1536(.a(_w_1868),.q(_w_1869));
  bfr _b_1535(.a(_w_1867),.q(_w_1868));
  bfr _b_1533(.a(_w_1865),.q(_w_1866));
  bfr _b_1541(.a(_w_1873),.q(_w_1874));
  bfr _b_1528(.a(_w_1860),.q(_w_1861));
  bfr _b_1523(.a(_w_1855),.q(_w_1856));
  bfr _b_1522(.a(_w_1854),.q(_w_1855));
  bfr _b_1521(.a(_w_1853),.q(_w_1854));
  bfr _b_1520(.a(_w_1852),.q(_w_1853));
  bfr _b_1519(.a(_w_1851),.q(_w_1852));
  bfr _b_1516(.a(_w_1848),.q(_w_1849));
  bfr _b_1515(.a(_w_1847),.q(N864));
  bfr _b_1513(.a(_w_1845),.q(_w_1846));
  bfr _b_1512(.a(_w_1844),.q(_w_1845));
  bfr _b_1782(.a(_w_2114),.q(_w_2115));
  bfr _b_1507(.a(_w_1839),.q(_w_1840));
  bfr _b_1506(.a(_w_1838),.q(_w_1839));
  bfr _b_1504(.a(_w_1836),.q(_w_1837));
  bfr _b_1503(.a(_w_1835),.q(_w_1836));
  bfr _b_1500(.a(_w_1832),.q(n243));
  bfr _b_1499(.a(_w_1831),.q(n242));
  bfr _b_1497(.a(_w_1829),.q(_w_1830));
  bfr _b_1496(.a(_w_1828),.q(_w_1829));
  bfr _b_1495(.a(_w_1827),.q(_w_1828));
  bfr _b_1493(.a(_w_1825),.q(N143_1));
  bfr _b_1491(.a(_w_1823),.q(_w_1824));
  bfr _b_1490(.a(_w_1822),.q(N863));
  bfr _b_1489(.a(_w_1821),.q(_w_1822));
  bfr _b_1480(.a(_w_1812),.q(_w_1813));
  bfr _b_1479(.a(_w_1811),.q(_w_1812));
  bfr _b_1475(.a(_w_1807),.q(_w_1808));
  bfr _b_1474(.a(_w_1806),.q(_w_1807));
  bfr _b_1785(.a(N246),.q(_w_2118));
  bfr _b_1473(.a(_w_1805),.q(_w_1806));
  bfr _b_1472(.a(_w_1804),.q(_w_1805));
  bfr _b_1471(.a(_w_1803),.q(N261_1));
  bfr _b_1468(.a(_w_1800),.q(_w_1801));
  bfr _b_1734(.a(N177),.q(_w_2066));
  bfr _b_1466(.a(_w_1798),.q(_w_1799));
  bfr _b_1465(.a(_w_1797),.q(_w_1798));
  bfr _b_1462(.a(_w_1794),.q(_w_1795));
  bfr _b_1459(.a(_w_1791),.q(_w_1792));
  bfr _b_1458(.a(_w_1790),.q(_w_1791));
  bfr _b_1456(.a(_w_1788),.q(_w_1789));
  bfr _b_1455(.a(_w_1787),.q(_w_1788));
  bfr _b_1454(.a(_w_1786),.q(_w_1787));
  bfr _b_1756(.a(_w_2088),.q(_w_2089));
  bfr _b_1453(.a(_w_1785),.q(_w_1786));
  bfr _b_1450(.a(_w_1782),.q(_w_1783));
  bfr _b_1449(.a(_w_1781),.q(_w_1782));
  bfr _b_1445(.a(_w_1777),.q(_w_1778));
  bfr _b_1444(.a(_w_1776),.q(_w_1777));
  bfr _b_1442(.a(_w_1774),.q(_w_1775));
  bfr _b_1461(.a(_w_1793),.q(_w_1794));
  bfr _b_1441(.a(_w_1773),.q(_w_1774));
  bfr _b_1440(.a(_w_1772),.q(_w_1773));
  bfr _b_1433(.a(_w_1765),.q(_w_1766));
  bfr _b_1432(.a(_w_1764),.q(_w_1765));
  bfr _b_1585(.a(_w_1917),.q(_w_1918));
  bfr _b_1431(.a(_w_1763),.q(_w_1764));
  bfr _b_1429(.a(_w_1761),.q(_w_1762));
  bfr _b_1427(.a(_w_1759),.q(_w_1760));
  bfr _b_1426(.a(_w_1758),.q(_w_1759));
  bfr _b_1548(.a(_w_1880),.q(_w_1881));
  bfr _b_1424(.a(_w_1756),.q(_w_1757));
  bfr _b_1423(.a(_w_1755),.q(_w_1756));
  bfr _b_1422(.a(_w_1754),.q(n71));
  bfr _b_1673(.a(_w_2005),.q(n67_2));
  bfr _b_1420(.a(_w_1752),.q(_w_1753));
  bfr _b_1419(.a(_w_1751),.q(_w_1752));
  bfr _b_1418(.a(_w_1750),.q(_w_1751));
  bfr _b_1417(.a(_w_1749),.q(_w_1750));
  bfr _b_1571(.a(_w_1903),.q(_w_1904));
  bfr _b_1412(.a(_w_1744),.q(_w_1745));
  bfr _b_1410(.a(_w_1742),.q(_w_1743));
  bfr _b_1409(.a(_w_1741),.q(_w_1742));
  bfr _b_1408(.a(_w_1740),.q(_w_1741));
  bfr _b_1407(.a(_w_1739),.q(_w_1740));
  bfr _b_1406(.a(_w_1738),.q(_w_1739));
  bfr _b_1795(.a(_w_2127),.q(_w_2117));
  bfr _b_1405(.a(_w_1737),.q(_w_1738));
  bfr _b_1635(.a(_w_1967),.q(_w_1968));
  bfr _b_1404(.a(_w_1736),.q(_w_1737));
  bfr _b_1403(.a(_w_1735),.q(_w_1736));
  bfr _b_1402(.a(_w_1734),.q(_w_1735));
  bfr _b_1398(.a(_w_1730),.q(_w_1731));
  bfr _b_1396(.a(_w_1728),.q(_w_1729));
  bfr _b_1394(.a(_w_1726),.q(n258));
  bfr _b_1391(.a(_w_1723),.q(N17_1));
  bfr _b_1700(.a(_w_2032),.q(_w_2033));
  bfr _b_1388(.a(_w_1720),.q(_w_1721));
  bfr _b_1384(.a(_w_1716),.q(_w_1717));
  bfr _b_1381(.a(_w_1713),.q(_w_1714));
  bfr _b_1380(.a(_w_1712),.q(_w_1713));
  bfr _b_1379(.a(_w_1711),.q(_w_1712));
  bfr _b_1378(.a(_w_1710),.q(_w_1711));
  bfr _b_1377(.a(_w_1709),.q(_w_1710));
  bfr _b_1413(.a(_w_1745),.q(_w_1746));
  bfr _b_1375(.a(_w_1707),.q(_w_1708));
  bfr _b_1374(.a(_w_1706),.q(_w_1707));
  bfr _b_1373(.a(_w_1705),.q(_w_1706));
  bfr _b_1371(.a(_w_1703),.q(_w_1704));
  bfr _b_1707(.a(_w_2039),.q(_w_2040));
  bfr _b_1369(.a(_w_1701),.q(_w_1702));
  bfr _b_1639(.a(_w_1971),.q(_w_1972));
  bfr _b_1366(.a(_w_1698),.q(_w_1699));
  bfr _b_1364(.a(_w_1696),.q(_w_1697));
  bfr _b_1360(.a(_w_1692),.q(_w_1693));
  bfr _b_1834(.a(_w_2166),.q(_w_2167));
  bfr _b_1359(.a(_w_1691),.q(_w_1692));
  bfr _b_1357(.a(_w_1689),.q(_w_1690));
  bfr _b_1356(.a(_w_1688),.q(_w_1689));
  bfr _b_1660(.a(_w_1992),.q(_w_1993));
  bfr _b_1355(.a(_w_1687),.q(_w_1688));
  bfr _b_1354(.a(_w_1686),.q(_w_1687));
  bfr _b_1351(.a(_w_1683),.q(N228_5));
  bfr _b_1350(.a(_w_1682),.q(_w_1683));
  bfr _b_1349(.a(_w_1681),.q(n189));
  bfr _b_1348(.a(_w_1680),.q(n241));
  bfr _b_1347(.a(_w_1679),.q(_w_1680));
  bfr _b_1460(.a(_w_1792),.q(_w_1793));
  bfr _b_1345(.a(_w_1677),.q(_w_1678));
  bfr _b_1626(.a(_w_1958),.q(_w_1959));
  bfr _b_1341(.a(_w_1673),.q(_w_1674));
  bfr _b_1338(.a(_w_1670),.q(_w_1671));
  bfr _b_1337(.a(_w_1669),.q(_w_1670));
  bfr _b_1336(.a(_w_1668),.q(_w_1669));
  bfr _b_1335(.a(_w_1667),.q(_w_1668));
  bfr _b_1334(.a(_w_1666),.q(_w_1667));
  bfr _b_1330(.a(_w_1662),.q(_w_1663));
  bfr _b_1329(.a(_w_1661),.q(_w_1662));
  bfr _b_1328(.a(_w_1660),.q(_w_1661));
  bfr _b_1325(.a(_w_1657),.q(n75));
  bfr _b_1810(.a(_w_2142),.q(_w_2143));
  bfr _b_1669(.a(_w_2001),.q(_w_2002));
  bfr _b_1332(.a(_w_1664),.q(_w_1665));
  bfr _b_1322(.a(_w_1654),.q(_w_1655));
  bfr _b_1321(.a(_w_1653),.q(n200_1));
  bfr _b_1320(.a(_w_1652),.q(_w_1653));
  bfr _b_1525(.a(_w_1857),.q(N106_2));
  bfr _b_1319(.a(_w_1651),.q(n256));
  bfr _b_1317(.a(_w_1649),.q(_w_1650));
  bfr _b_1314(.a(_w_1646),.q(_w_1647));
  bfr _b_1312(.a(_w_1644),.q(_w_1645));
  bfr _b_1397(.a(_w_1729),.q(_w_1730));
  bfr _b_1311(.a(_w_1643),.q(_w_1644));
  bfr _b_1307(.a(_w_1639),.q(N447));
  bfr _b_1306(.a(_w_1638),.q(_w_1639));
  bfr _b_1305(.a(_w_1637),.q(_w_1638));
  bfr _b_1304(.a(_w_1636),.q(_w_1637));
  bfr _b_1303(.a(_w_1635),.q(_w_1636));
  bfr _b_1302(.a(_w_1634),.q(_w_1635));
  bfr _b_1301(.a(_w_1633),.q(_w_1634));
  bfr _b_1300(.a(_w_1632),.q(_w_1633));
  bfr _b_1818(.a(N51),.q(_w_2150));
  bfr _b_1298(.a(_w_1630),.q(_w_1631));
  bfr _b_1297(.a(_w_1629),.q(_w_1630));
  bfr _b_1295(.a(_w_1627),.q(_w_1628));
  bfr _b_1294(.a(_w_1626),.q(_w_1627));
  bfr _b_1654(.a(_w_1986),.q(_w_1987));
  bfr _b_1291(.a(_w_1623),.q(_w_1624));
  bfr _b_1290(.a(_w_1622),.q(_w_1623));
  bfr _b_1289(.a(_w_1621),.q(_w_1622));
  bfr _b_1514(.a(_w_1846),.q(_w_1847));
  bfr _b_1287(.a(_w_1619),.q(_w_1620));
  bfr _b_1283(.a(_w_1615),.q(_w_1616));
  bfr _b_1282(.a(_w_1614),.q(_w_1615));
  bfr _b_1327(.a(_w_1659),.q(_w_1660));
  bfr _b_1280(.a(_w_1612),.q(_w_1613));
  bfr _b_1279(.a(_w_1611),.q(_w_1612));
  bfr _b_1276(.a(_w_1608),.q(_w_1609));
  bfr _b_1275(.a(_w_1607),.q(_w_1608));
  bfr _b_1274(.a(_w_1606),.q(_w_1607));
  bfr _b_1278(.a(_w_1610),.q(_w_1611));
  bfr _b_1272(.a(_w_1604),.q(N422));
  bfr _b_1683(.a(_w_2015),.q(_w_2016));
  bfr _b_1268(.a(_w_1600),.q(_w_1601));
  bfr _b_1277(.a(_w_1609),.q(_w_1610));
  bfr _b_1267(.a(_w_1599),.q(_w_1600));
  bfr _b_1264(.a(_w_1596),.q(_w_1597));
  bfr _b_1299(.a(_w_1631),.q(_w_1632));
  bfr _b_1262(.a(_w_1594),.q(_w_1595));
  bfr _b_1260(.a(_w_1592),.q(_w_1593));
  bfr _b_1259(.a(_w_1591),.q(_w_1592));
  bfr _b_1254(.a(_w_1586),.q(_w_1587));
  bfr _b_1253(.a(_w_1585),.q(_w_1586));
  bfr _b_1250(.a(_w_1582),.q(_w_1583));
  bfr _b_1249(.a(_w_1581),.q(_w_1582));
  bfr _b_1248(.a(_w_1580),.q(_w_1581));
  bfr _b_1771(.a(N237),.q(_w_2104));
  bfr _b_1372(.a(_w_1704),.q(_w_1705));
  bfr _b_1246(.a(_w_1578),.q(_w_1579));
  bfr _b_1245(.a(_w_1577),.q(_w_1578));
  bfr _b_1242(.a(_w_1574),.q(_w_1575));
  bfr _b_1241(.a(_w_1573),.q(_w_1574));
  bfr _b_1240(.a(_w_1572),.q(_w_1573));
  bfr _b_1324(.a(_w_1656),.q(_w_1657));
  bfr _b_1235(.a(_w_1567),.q(N420));
  bfr _b_1234(.a(_w_1566),.q(_w_1567));
  bfr _b_1233(.a(_w_1565),.q(_w_1566));
  bfr _b_1361(.a(_w_1693),.q(_w_1694));
  bfr _b_1232(.a(_w_1564),.q(_w_1565));
  bfr _b_1230(.a(_w_1562),.q(_w_1563));
  bfr _b_1229(.a(_w_1561),.q(_w_1562));
  bfr _b_1228(.a(_w_1560),.q(_w_1561));
  bfr _b_1227(.a(_w_1559),.q(_w_1560));
  bfr _b_1370(.a(_w_1702),.q(_w_1703));
  bfr _b_1323(.a(_w_1655),.q(N268_3));
  bfr _b_1226(.a(_w_1558),.q(_w_1559));
  bfr _b_1224(.a(_w_1556),.q(_w_1557));
  bfr _b_1222(.a(_w_1554),.q(_w_1555));
  bfr _b_1221(.a(_w_1553),.q(_w_1554));
  bfr _b_1806(.a(_w_2138),.q(_w_2139));
  bfr _b_1598(.a(_w_1930),.q(_w_1931));
  bfr _b_1270(.a(_w_1602),.q(_w_1603));
  bfr _b_1263(.a(_w_1595),.q(_w_1596));
  bfr _b_1220(.a(_w_1552),.q(_w_1553));
  bfr _b_1219(.a(_w_1551),.q(_w_1552));
  bfr _b_1443(.a(_w_1775),.q(_w_1776));
  bfr _b_1216(.a(_w_1548),.q(_w_1549));
  bfr _b_1362(.a(_w_1694),.q(_w_1695));
  bfr _b_1215(.a(_w_1547),.q(_w_1548));
  bfr _b_1214(.a(_w_1546),.q(_w_1547));
  bfr _b_1213(.a(_w_1545),.q(_w_1546));
  bfr _b_1211(.a(_w_1543),.q(_w_1544));
  bfr _b_1207(.a(_w_1539),.q(_w_1540));
  bfr _b_1206(.a(_w_1538),.q(_w_1539));
  bfr _b_1205(.a(_w_1537),.q(_w_1538));
  bfr _b_1204(.a(_w_1536),.q(_w_1537));
  bfr _b_1201(.a(_w_1533),.q(n283));
  bfr _b_1615(.a(_w_1947),.q(_w_1948));
  bfr _b_1200(.a(_w_1532),.q(N390));
  bfr _b_1549(.a(_w_1881),.q(n183));
  bfr _b_1199(.a(_w_1531),.q(n169));
  bfr _b_1198(.a(_w_1530),.q(n239));
  bfr _b_1196(.a(_w_1528),.q(_w_1529));
  bfr _b_1194(.a(_w_1526),.q(_w_1527));
  bfr _b_1192(.a(_w_1524),.q(N391));
  bfr _b_1191(.a(_w_1523),.q(_w_1524));
  bfr _b_1190(.a(_w_1522),.q(_w_1523));
  bfr _b_1189(.a(_w_1521),.q(_w_1522));
  bfr _b_1790(.a(_w_2122),.q(_w_2123));
  bfr _b_1188(.a(_w_1520),.q(_w_1521));
  bfr _b_1187(.a(_w_1519),.q(_w_1520));
  bfr _b_1822(.a(_w_2154),.q(_w_2153));
  bfr _b_1186(.a(_w_1518),.q(_w_1519));
  bfr _b_1389(.a(_w_1721),.q(_w_1722));
  bfr _b_1183(.a(_w_1515),.q(_w_1516));
  bfr _b_1180(.a(_w_1512),.q(_w_1513));
  bfr _b_1798(.a(N260),.q(_w_2130));
  bfr _b_1179(.a(_w_1511),.q(_w_1512));
  bfr _b_1178(.a(_w_1510),.q(_w_1511));
  bfr _b_1177(.a(_w_1509),.q(_w_1510));
  bfr _b_1176(.a(_w_1508),.q(_w_1509));
  bfr _b_1174(.a(_w_1506),.q(_w_1507));
  bfr _b_1173(.a(_w_1505),.q(_w_1506));
  bfr _b_1838(.a(_w_2170),.q(_w_2165));
  bfr _b_1266(.a(_w_1598),.q(_w_1599));
  bfr _b_1172(.a(_w_1504),.q(_w_1505));
  bfr _b_1171(.a(_w_1503),.q(_w_1504));
  bfr _b_1751(.a(_w_2083),.q(_w_2084));
  bfr _b_1170(.a(_w_1502),.q(_w_1503));
  bfr _b_1169(.a(_w_1501),.q(_w_1502));
  bfr _b_1168(.a(_w_1500),.q(_w_1501));
  bfr _b_1167(.a(_w_1499),.q(_w_1500));
  bfr _b_1166(.a(_w_1498),.q(_w_1499));
  bfr _b_1163(.a(_w_1495),.q(_w_1496));
  bfr _b_1716(.a(_w_2048),.q(_w_2049));
  bfr _b_1162(.a(_w_1494),.q(_w_1495));
  bfr _b_1161(.a(_w_1493),.q(_w_1494));
  bfr _b_1159(.a(_w_1491),.q(_w_1492));
  bfr _b_1158(.a(_w_1490),.q(_w_1491));
  bfr _b_1157(.a(_w_1489),.q(_w_1490));
  bfr _b_1156(.a(_w_1488),.q(_w_1489));
  bfr _b_1154(.a(_w_1486),.q(_w_1487));
  bfr _b_1153(.a(_w_1485),.q(n61_1));
  bfr _b_1152(.a(_w_1484),.q(_w_1485));
  bfr _b_1148(.a(_w_1480),.q(_w_1481));
  bfr _b_1147(.a(_w_1479),.q(_w_1480));
  bfr _b_1146(.a(_w_1478),.q(_w_1479));
  bfr _b_1141(.a(_w_1473),.q(_w_1474));
  bfr _b_1140(.a(_w_1472),.q(_w_1473));
  bfr _b_1138(.a(_w_1470),.q(_w_1471));
  bfr _b_1137(.a(_w_1469),.q(_w_1470));
  bfr _b_1136(.a(_w_1468),.q(_w_1469));
  bfr _b_1134(.a(_w_1466),.q(_w_1467));
  bfr _b_1133(.a(_w_1465),.q(_w_1466));
  bfr _b_1132(.a(_w_1464),.q(_w_1465));
  bfr _b_1293(.a(_w_1625),.q(_w_1626));
  bfr _b_1131(.a(_w_1463),.q(_w_1464));
  bfr _b_1129(.a(_w_1461),.q(_w_1462));
  bfr _b_1128(.a(_w_1460),.q(_w_1461));
  bfr _b_1127(.a(_w_1459),.q(_w_1460));
  bfr _b_1125(.a(_w_1457),.q(_w_1458));
  bfr _b_1124(.a(_w_1456),.q(_w_1457));
  bfr _b_1160(.a(_w_1492),.q(_w_1493));
  bfr _b_1122(.a(_w_1454),.q(_w_1455));
  bfr _b_1120(.a(_w_1452),.q(_w_1453));
  bfr _b_1118(.a(_w_1450),.q(_w_1451));
  bfr _b_1114(.a(_w_1446),.q(_w_1447));
  bfr _b_1113(.a(_w_1445),.q(_w_1446));
  bfr _b_1111(.a(_w_1443),.q(N177_4));
  bfr _b_1110(.a(_w_1442),.q(_w_1443));
  bfr _b_1109(.a(_w_1441),.q(_w_1442));
  bfr _b_538(.a(_w_870),.q(_w_871));
  bfr _b_536(.a(_w_868),.q(_w_869));
  and_bb g97(.a(N121_1),.b(N135_1),.q(n97));
  bfr _b_656(.a(_w_988),.q(_w_989));
  bfr _b_530(.a(_w_862),.q(N210_3));
  bfr _b_523(.a(_w_855),.q(N201_2));
  bfr _b_522(.a(_w_854),.q(_w_855));
  bfr _b_517(.a(_w_849),.q(N201_4));
  bfr _b_513(.a(_w_845),.q(N195_2));
  and_bb g271(.a(N159_5),.b(n270_2),.q(_w_1888));
  bfr _b_511(.a(_w_843),.q(_w_844));
  bfr _b_508(.a(_w_840),.q(_w_841));
  bfr _b_1310(.a(_w_1642),.q(n362));
  and_bb g93(.a(N91_0),.b(n92_0),.q(n93));
  bfr _b_562(.a(_w_894),.q(_w_895));
  bfr _b_1640(.a(_w_1972),.q(_w_1973));
  bfr _b_504(.a(_w_836),.q(_w_837));
  bfr _b_1816(.a(_w_2148),.q(_w_2149));
  and_bb g253(.a(N195_3),.b(n179_2),.q(n253));
  bfr _b_1650(.a(_w_1982),.q(_w_1983));
  spl3L g228_s_0(.a(n228),.q0(n228_0),.q1(n228_1),.q2(n228_2));
  spl3L g295_s_0(.a(n295),.q0(n295_0),.q1(n295_1),.q2(_w_831));
  bfr _b_789(.a(_w_1121),.q(_w_1122));
  spl3L N246_s_1(.a(N246_0),.q0(N246_2),.q1(N246_3),.q2(N246_4));
  spl2 N195_s_1(.a(N195_2),.q0(N195_3),.q1(_w_835));
  bfr _b_1483(.a(_w_1815),.q(_w_1816));
  bfr _b_737(.a(_w_1069),.q(_w_1070));
  bfr _b_1820(.a(N72),.q(_w_2152));
  spl3L N195_s_0(.a(N195),.q0(N195_0),.q1(N195_1),.q2(_w_840));
  spl2 N201_s_1(.a(N201_2),.q0(N201_3),.q1(_w_846));
  or_bb g185(.a(n175),.b(n184),.q(_w_1105));
  spl3L N201_s_0(.a(N201),.q0(N201_0),.q1(N201_1),.q2(_w_850));
  bfr _b_934(.a(_w_1266),.q(_w_1267));
  bfr _b_1470(.a(_w_1802),.q(n223));
  spl2 g179_s_1(.a(n179_3),.q0(n179_4),.q1(n179_5));
  spl2 g210_s_1(.a(n210_1),.q0(n210_2),.q1(n210_3));
  bfr _b_1117(.a(_w_1449),.q(_w_1450));
  or_bb g187(.a(n173),.b(n186),.q(_w_1225));
  spl4L N210_s_0(.a(N210),.q0(N210_0),.q1(N210_1),.q2(N210_2),.q3(_w_856));
  spl2 g166_s_0(.a(n166),.q0(n166_0),.q1(_w_863));
  or_bb g197(.a(n152_1),.b(n196),.q(n197));
  spl2 g286_s_1(.a(n286_1),.q0(n286_2),.q1(n286_3));
  bfr _b_820(.a(_w_1152),.q(_w_1153));
  bfr _b_1485(.a(_w_1817),.q(_w_1818));
  spl2 g134_s_0(.a(n134),.q0(n134_0),.q1(n134_1));
  spl2 N51_s_1(.a(N51_1),.q0(N51_2),.q1(N51_3));
  spl2 g198_s_0(.a(n198),.q0(n198_0),.q1(n198_1));
  bfr _b_1809(.a(_w_2141),.q(_w_2142));
  bfr _b_1663(.a(_w_1995),.q(_w_1996));
  spl2 g152_s_1(.a(n152_2),.q0(n152_3),.q1(_w_867));
  bfr _b_541(.a(_w_873),.q(_w_874));
  spl2 g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1));
  spl4L g147_s_0(.a(n147),.q0(n147_0),.q1(n147_1),.q2(n147_2),.q3(n147_3));
  spl2 g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1));
  bfr _b_1237(.a(_w_1569),.q(_w_1570));
  bfr _b_713(.a(_w_1045),.q(_w_1046));
  and_bb g203(.a(n200_1),.b(n202_0),.q(n203));
  or_bb g105(.a(N111_0),.b(N116_0),.q(n105));
  bfr _b_1826(.a(N80),.q(_w_2159));
  bfr _b_1463(.a(_w_1795),.q(_w_1796));
  spl2 N189_s_1(.a(N189_2),.q0(N189_3),.q1(_w_925));
  and_bb g281(.a(N101_3),.b(n162_8),.q(n281));
  bfr _b_1428(.a(_w_1760),.q(_w_1761));
  bfr _b_1376(.a(_w_1708),.q(_w_1709));
  bfr _b_1039(.a(_w_1371),.q(_w_1372));
  spl2 N228_s_3(.a(N228_5),.q0(N228_6),.q1(_w_870));
  and_bb g169(.a(N261_3),.b(n168_2),.q(_w_1531));
  spl2 N171_s_1(.a(N171_2),.q0(N171_3),.q1(_w_1568));
  bfr _b_525(.a(_w_857),.q(_w_858));
  spl2 g122_s_0(.a(n122),.q0(n122_0),.q1(n122_1));
  and_bi g141(.a(n122_0),.b(n140_0),.q(n141));
  bfr _b_510(.a(_w_842),.q(_w_843));
  spl2 N159_s_2(.a(N159_4),.q0(N159_5),.q1(N159_6));
  spl2 N159_s_1(.a(N159_2),.q0(N159_3),.q1(_w_873));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(n119_1));
  bfr _b_750(.a(_w_1082),.q(N219_10));
  bfr _b_1368(.a(_w_1700),.q(_w_1701));
  bfr _b_658(.a(_w_990),.q(_w_991));
  spl2 N13_s_0(.a(_w_2026),.q0(N13_0),.q1(_w_876));
  spl4L N111_s_0(.a(N111),.q0(N111_0),.q1(N111_1),.q2(N111_2),.q3(_w_881));
  spl3L g287_s_0(.a(n287),.q0(n287_0),.q1(n287_1),.q2(_w_890));
  and_bi g129(.a(N201_0),.b(N165_0),.q(n129));
  spl2 N149_s_0(.a(_w_2046),.q0(N149_0),.q1(_w_893));
  bfr _b_1524(.a(_w_1856),.q(_w_1857));
  spl3L N126_s_0(.a(_w_2023),.q0(N126_0),.q1(N126_1),.q2(_w_894));
  bfr _b_1721(.a(_w_2053),.q(_w_2046));
  bfr _b_577(.a(_w_909),.q(_w_910));
  spl2 g144_s_0(.a(n144),.q0(n144_0),.q1(n144_1));
  spl2 N195_s_2(.a(N195_4),.q0(N195_5),.q1(N195_6));
  bfr _b_1042(.a(_w_1374),.q(_w_1375));
  bfr _b_1043(.a(_w_1375),.q(_w_1376));
  bfr _b_1715(.a(_w_2047),.q(_w_2048));
  or_bb g111(.a(n101_0),.b(n110_0),.q(n111));
  spl2 N165_s_2(.a(N165_4),.q0(N165_5),.q1(N165_6));
  bfr _b_716(.a(_w_1048),.q(_w_1049));
  spl2 N165_s_1(.a(N165_2),.q0(N165_3),.q1(_w_903));
  bfr _b_524(.a(_w_856),.q(_w_857));
  bfr _b_745(.a(_w_1077),.q(n320));
  bfr _b_528(.a(_w_860),.q(_w_861));
  or_bb g276(.a(n266_1),.b(n275),.q(n276));
  spl4L N121_s_0(.a(N121),.q0(N121_0),.q1(N121_1),.q2(N121_2),.q3(_w_908));
  bfr _b_1352(.a(_w_1684),.q(_w_1685));
  spl2 N210_s_1(.a(N210_3),.q0(N210_4),.q1(N210_5));
  bfr _b_1251(.a(_w_1583),.q(_w_1584));
  bfr _b_587(.a(_w_919),.q(_w_920));
  bfr _b_1098(.a(_w_1430),.q(_w_1431));
  spl2 N183_s_1(.a(N183_2),.q0(N183_3),.q1(_w_916));
  spl3L g206_s_0(.a(n206),.q0(n206_0),.q1(n206_1),.q2(n206_2));
  bfr _b_932(.a(_w_1264),.q(_w_1265));
  bfr _b_1339(.a(_w_1671),.q(_w_1672));
  spl2 N189_s_2(.a(N189_4),.q0(N189_5),.q1(N189_6));
  spl2 N17_s_4(.a(N17_8),.q0(N17_9),.q1(N17_10));
  bfr _b_1144(.a(_w_1476),.q(_w_1477));
  spl2 N183_s_2(.a(N183_4),.q0(N183_5),.q1(N183_6));
  spl2 N246_s_3(.a(N246_8),.q0(N246_9),.q1(N246_10));
  bfr _b_1115(.a(_w_1447),.q(_w_1448));
  spl2 g73_s_0(.a(n73),.q0(n73_0),.q1(_w_974));
  and_bi g102(.a(N101_0),.b(N106_0),.q(n102));
  bfr _b_1150(.a(_w_1482),.q(_w_1483));
  spl3L N189_s_0(.a(N189),.q0(N189_0),.q1(N189_1),.q2(_w_931));
  and_bb g234(.a(N237_4),.b(n193_1),.q(n234));
  bfr _b_515(.a(_w_847),.q(_w_848));
  bfr _b_1709(.a(_w_2041),.q(_w_2042));
  spl2 g125_s_0(.a(n125),.q0(n125_0),.q1(n125_1));
  spl2 g101_s_0(.a(n101),.q0(n101_0),.q1(n101_1));
  bfr _b_514(.a(_w_846),.q(_w_847));
  spl2 g71_s_0(.a(n71),.q0(n71_0),.q1(n71_1));
  bfr _b_1775(.a(_w_2107),.q(_w_2108));
  bfr _b_1193(.a(_w_1525),.q(_w_1526));
  spl2 N219_s_6(.a(N219_12),.q0(N219_13),.q1(_w_937));
  spl2 N219_s_5(.a(N219_10),.q0(N219_11),.q1(_w_940));
  spl2 g110_s_0(.a(n110),.q0(n110_0),.q1(n110_1));
  spl2 N228_s_1(.a(N228_1),.q0(N228_2),.q1(_w_942));
  spl2 N219_s_2(.a(N219_3),.q0(N219_4),.q1(_w_944));
  and_bb g295(.a(N177_5),.b(n294_2),.q(_w_1992));
  bfr _b_1083(.a(_w_1415),.q(_w_1416));
  spl2 N237_s_5(.a(N237_9),.q0(N237_10),.q1(_w_949));
  spl2 N237_s_2(.a(N237_3),.q0(N237_4),.q1(_w_952));
  bfr _b_1488(.a(_w_1820),.q(_w_1821));
  bfr _b_1333(.a(_w_1665),.q(_w_1666));
  bfr _b_589(.a(_w_921),.q(_w_922));
  bfr _b_712(.a(_w_1044),.q(_w_1045));
  spl2 N237_s_0(.a(_w_2103),.q0(N237_0),.q1(N237_1));
  bfr _b_1784(.a(_w_2116),.q(_w_2103));
  and_bb g251(.a(N237_2),.b(n199_1),.q(n251));
  spl2 N55_s_1(.a(N55_1),.q0(N55_2),.q1(N55_3));
  bfr _b_1387(.a(_w_1719),.q(_w_1720));
  spl2 N55_s_0(.a(_w_2151),.q0(N55_0),.q1(_w_956));
  spl2 g145_s_0(.a(n145),.q0(n145_0),.q1(n145_1));
  spl3L N255_s_0(.a(N255),.q0(N255_0),.q1(N255_1),.q2(N255_2));
  spl2 N68_s_0(.a(N68),.q0(N68_0),.q1(_w_960));
  spl3L N91_s_0(.a(_w_2165),.q0(N91_0),.q1(N91_1),.q2(_w_961));
  spl2 N153_s_0(.a(_w_2055),.q0(N153_0),.q1(_w_1924));
  spl2 N17_s_3(.a(N17_6),.q0(_w_963),.q1(N17_8));
  bfr _b_785(.a(_w_1117),.q(N1_2));
  bfr _b_815(.a(_w_1147),.q(_w_1148));
  bfr _b_1055(.a(_w_1387),.q(_w_1388));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(_w_964));
  spl2 g192_s_1(.a(n192_1),.q0(n192_2),.q1(n192_3));
  spl3L N42_s_2(.a(N42_3),.q0(N42_4),.q1(N42_5),.q2(N42_6));
  bfr _b_1236(.a(_w_1568),.q(_w_1569));
  and_bb g67(.a(N1_0),.b(N8_0),.q(n67));
  bfr _b_1833(.a(N91),.q(_w_2166));
  spl2 N237_s_4(.a(N237_7),.q0(N237_8),.q1(_w_1108));
  bfr _b_1606(.a(_w_1938),.q(_w_1939));
  bfr _b_1447(.a(_w_1779),.q(_w_1780));
  bfr _b_1073(.a(_w_1405),.q(_w_1406));
  bfr _b_1399(.a(_w_1731),.q(_w_1732));
  spl2 N228_s_6(.a(N228_11),.q0(N228_12),.q1(_w_965));
  bfr _b_1411(.a(_w_1743),.q(_w_1744));
  bfr _b_843(.a(_w_1175),.q(N390_0));
  bfr _b_1662(.a(_w_1994),.q(_w_1995));
  spl3L N96_s_0(.a(_w_2171),.q0(N96_0),.q1(N96_1),.q2(_w_969));
  bfr _b_1484(.a(_w_1816),.q(_w_1817));
  or_bb g294(.a(n289),.b(n293),.q(n294));
  bfr _b_1759(.a(_w_2091),.q(_w_2092));
  spl2 g162_s_1(.a(n162_2),.q0(n162_4),.q1(n162_5));
  bfr _b_516(.a(_w_848),.q(_w_849));
  bfr _b_507(.a(_w_839),.q(N195_4));
  spl2 g70_s_0(.a(n70),.q0(n70_0),.q1(_w_979));
  spl2 N237_s_1(.a(N237_1),.q0(N237_2),.q1(_w_954));
  bfr _b_821(.a(_w_1153),.q(_w_1154));
  spl2 N80_s_0(.a(_w_2158),.q0(N80_0),.q1(N80_1));
  bfr _b_1487(.a(_w_1819),.q(_w_1820));
  bfr _b_1012(.a(_w_1344),.q(_w_1345));
  bfr _b_1561(.a(_w_1893),.q(_w_1894));
  bfr _b_730(.a(_w_1062),.q(_w_1063));
  bfr _b_1256(.a(_w_1588),.q(_w_1589));
  bfr _b_765(.a(_w_1097),.q(_w_1098));
  spl2 g95_s_0(.a(n95),.q0(n95_0),.q1(n95_1));
  bfr _b_1126(.a(_w_1458),.q(_w_1459));
  spl3L N101_s_0(.a(N101),.q0(N101_0),.q1(N101_1),.q2(_w_987));
  spl4L N246_s_2(.a(N246_1),.q0(N246_5),.q1(N246_6),.q2(N246_7),.q3(N246_8));
  or_bb g137(.a(n135),.b(n136),.q(n137));
  spl2 N171_s_2(.a(N171_4),.q0(N171_5),.q1(N171_6));
  bfr _b_1030(.a(_w_1362),.q(_w_1363));
  bfr _b_1119(.a(_w_1451),.q(_w_1452));
  spl2 N130_s_1(.a(N130_2),.q0(N130_3),.q1(N130_4));
  spl2 N228_s_0(.a(_w_2087),.q0(N228_0),.q1(N228_1));
  bfr _b_748(.a(_w_1080),.q(_w_1081));
  bfr _b_1597(.a(_w_1929),.q(n275));
  bfr _b_537(.a(_w_869),.q(N228_11));
  spl2 N246_s_0(.a(_w_2117),.q0(N246_0),.q1(N246_1));
  bfr _b_1526(.a(_w_1858),.q(_w_1859));
  spl2 N42_s_3(.a(N42_6),.q0(N42_7),.q1(N42_8));
  or_bb g288(.a(N171_6),.b(n286_3),.q(_w_1755));
  spl2 g272_s_0(.a(n272),.q0(n272_0),.q1(_w_994));
  spl3L g279_s_0(.a(n279),.q0(n279_0),.q1(n279_1),.q2(_w_996));
  bfr _b_1316(.a(_w_1648),.q(_w_1649));
  and_bi g195(.a(N149_1),.b(n147_1),.q(n195));
  bfr _b_1451(.a(_w_1783),.q(_w_1784));
  bfr _b_1393(.a(_w_1725),.q(_w_1726));
  bfr _b_1343(.a(_w_1675),.q(_w_1676));
  bfr _b_795(.a(_w_1127),.q(_w_1128));
  spl4L g266_s_0(.a(n266),.q0(n266_0),.q1(n266_1),.q2(n266_2),.q3(n266_3));
  spl2 g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1));
  bfr _b_586(.a(_w_918),.q(_w_919));
  bfr _b_782(.a(_w_1114),.q(_w_1115));
  spl2 g212_s_0(.a(n212),.q0(n212_0),.q1(_w_1002));
  bfr _b_800(.a(_w_1132),.q(_w_1133));
  bfr _b_1026(.a(_w_1358),.q(N450));
  spl3L g337_s_0(.a(n337),.q0(n337_0),.q1(n337_1),.q2(n337_2));
  bfr _b_1342(.a(_w_1674),.q(_w_1675));
  or_bb g365(.a(n357),.b(n364),.q(_w_1004));
  or_bb g364(.a(n358),.b(n363),.q(_w_1005));
  bfr _b_532(.a(_w_864),.q(_w_865));
  or_bb g272(.a(N159_6),.b(n270_3),.q(_w_1906));
  bfr _b_1557(.a(_w_1889),.q(_w_1890));
  bfr _b_616(.a(_w_948),.q(N237_13));
  and_bb g359(.a(N246_7),.b(n286_0),.q(n359));
  bfr _b_1255(.a(_w_1587),.q(_w_1588));
  spl2 N207_s_0(.a(_w_2067),.q0(N207_0),.q1(N207_1));
  bfr _b_655(.a(_w_987),.q(_w_988));
  bfr _b_818(.a(_w_1150),.q(_w_1151));
  bfr _b_1552(.a(_w_1884),.q(_w_1885));
  bfr _b_637(.a(_w_969),.q(_w_970));
  bfr _b_981(.a(_w_1313),.q(_w_1314));
  bfr _b_1601(.a(_w_1933),.q(_w_1934));
  spl3L N159_s_0(.a(_w_2064),.q0(N159_0),.q1(N159_1),.q2(_w_1226));
  and_bb g355(.a(N219_11),.b(n354),.q(n355));
  and_bi g121(.a(n119_1),.b(N130_4),.q(n121));
  spl2 N42_s_0(.a(N42),.q0(N42_0),.q1(_w_968));
  or_bb g354(.a(n300_1),.b(n352_0),.q(n354));
  and_bb g326(.a(n323),.b(n325),.q(n326));
  and_bb g283(.a(N138_4),.b(N17_9),.q(_w_1533));
  and_bi g352(.a(n288_0),.b(n287_0),.q(n352));
  spl2 g307_s_0(.a(n307),.q0(n307_0),.q1(_w_1006));
  bfr _b_770(.a(_w_1102),.q(_w_1103));
  bfr _b_940(.a(_w_1272),.q(_w_1273));
  or_bb g349(.a(n343),.b(n348),.q(_w_1013));
  or_bb g183(.a(n181),.b(n182),.q(_w_1876));
  spl4L g162_s_2(.a(n162_3),.q0(n162_6),.q1(n162_7),.q2(n162_8),.q3(n162_9));
  or_bb g347(.a(n345),.b(n346),.q(_w_1031));
  or_bb g246(.a(n202_1),.b(n245_0),.q(n246));
  bfr _b_1121(.a(_w_1453),.q(_w_1454));
  bfr _b_695(.a(_w_1027),.q(_w_1028));
  spl3L g213_s_0(.a(n213),.q0(n213_0),.q1(n213_1),.q2(n213_2));
  and_bb g343(.a(N237_12),.b(n279_1),.q(n343));
  bfr _b_1655(.a(_w_1987),.q(_w_1988));
  and_bb g83(.a(n67_0),.b(n82),.q(n83));
  bfr _b_1467(.a(_w_1799),.q(N767));
  bfr _b_643(.a(_w_975),.q(n73_1));
  and_bb g342(.a(N228_12),.b(n337_1),.q(n342));
  bfr _b_535(.a(_w_867),.q(n152_4));
  and_bb g182(.a(N121_2),.b(N210_0),.q(n182));
  or_bb g191(.a(n152_3),.b(n190),.q(n191));
  bfr _b_690(.a(_w_1022),.q(_w_1023));
  and_bb g338(.a(n302_2),.b(n337_2),.q(_w_1033));
  or_bb g336(.a(n326),.b(n335),.q(N878));
  spl3L N106_s_0(.a(N106),.q0(N106_0),.q1(N106_1),.q2(_w_1850));
  or_bb g335(.a(n327),.b(n334),.q(_w_1034));
  bfr _b_1269(.a(_w_1601),.q(_w_1602));
  bfr _b_1087(.a(_w_1419),.q(_w_1420));
  bfr _b_1501(.a(_w_1833),.q(_w_1834));
  or_bb g334(.a(n328),.b(n333),.q(_w_1035));
  or_bb g333(.a(n329),.b(n332),.q(_w_1036));
  spl2 N177_s_2(.a(N177_4),.q0(N177_5),.q1(N177_6));
  or_bb g184(.a(n180),.b(n183),.q(_w_1083));
  bfr _b_1040(.a(_w_1372),.q(n363));
  or_bb g332(.a(n330),.b(n331),.q(_w_1056));
  spl4L N210_s_2(.a(N210_5),.q0(N210_6),.q1(N210_7),.q2(N210_8),.q3(N210_9));
  bfr _b_916(.a(_w_1248),.q(_w_1249));
  and_bb g330(.a(N159_3),.b(n179_6),.q(n330));
  bfr _b_1210(.a(_w_1542),.q(_w_1543));
  bfr _b_898(.a(_w_1230),.q(_w_1231));
  and_bb g328(.a(N237_13),.b(n271_1),.q(n328));
  spl2 N138_s_0(.a(N138),.q0(N138_0),.q1(_w_1066));
  bfr _b_969(.a(_w_1301),.q(_w_1302));
  bfr _b_1243(.a(_w_1575),.q(_w_1576));
  spl2 N237_s_3(.a(N237_5),.q0(N237_6),.q1(_w_951));
  and_bb g324(.a(n304_1),.b(n322_0),.q(n324));
  spl3L g245_s_0(.a(n245),.q0(n245_0),.q1(n245_1),.q2(n245_2));
  and_bi g337(.a(n280_0),.b(n279_0),.q(n337));
  and_bb g327(.a(N228_13),.b(n322_1),.q(n327));
  bfr _b_1092(.a(_w_1424),.q(_w_1425));
  and_bi g322(.a(n272_0),.b(n271_0),.q(n322));
  spl3L g302_s_0(.a(n302),.q0(n302_0),.q1(n302_1),.q2(n302_2));
  bfr _b_1815(.a(_w_2147),.q(_w_2148));
  bfr _b_1217(.a(_w_1549),.q(_w_1550));
  and_bb g361(.a(N171_3),.b(n179_8),.q(n361));
  or_bb g320(.a(n312),.b(n319),.q(_w_1077));
  bfr _b_1143(.a(_w_1475),.q(_w_1476));
  or_bb g319(.a(n313),.b(n318),.q(_w_1078));
  bfr _b_1670(.a(_w_2002),.q(_w_2003));
  bfr _b_505(.a(_w_837),.q(_w_838));
  spl2 N219_s_4(.a(N219_8),.q0(N219_9),.q1(_w_1080));
  bfr _b_602(.a(_w_934),.q(_w_935));
  or_bb g90(.a(N130_0),.b(N96_0),.q(n90));
  bfr _b_1517(.a(_w_1849),.q(n280_1));
  and_bb g264(.a(N143_0),.b(n263_0),.q(n264));
  bfr _b_1434(.a(_w_1766),.q(n288));
  spl2 g98_s_0(.a(n98),.q0(n98_0),.q1(n98_1));
  or_bb g186(.a(n174),.b(n185),.q(_w_1087));
  spl3L g168_s_0(.a(n168),.q0(n168_0),.q1(n168_1),.q2(n168_2));
  and_bb g358(.a(N237_10),.b(n287_1),.q(n358));
  and_bb g287(.a(N171_5),.b(n286_2),.q(_w_1088));
  or_bb g269(.a(n264),.b(n268),.q(n269));
  bfr _b_650(.a(_w_982),.q(_w_983));
  or_bb g257(.a(n253),.b(n256),.q(_w_1100));
  bfr _b_915(.a(_w_1247),.q(_w_1248));
  and_bi g110(.a(n108),.b(n109),.q(n110));
  bfr _b_605(.a(_w_937),.q(_w_938));
  bfr _b_1340(.a(_w_1672),.q(_w_1673));
  and_bb g173(.a(N228_0),.b(n168_1),.q(n173));
  bfr _b_1257(.a(_w_1589),.q(_w_1590));
  and_bb g252(.a(N246_3),.b(n198_0),.q(n252));
  or_bb g350(.a(n342),.b(n349),.q(_w_1012));
  bfr _b_527(.a(_w_859),.q(_w_860));
  bfr _b_1437(.a(_w_1769),.q(n225));
  spl3L g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1),.q2(n152_2));
  and_bb g171(.a(N219_0),.b(n170),.q(n171));
  bfr _b_1632(.a(_w_1964),.q(_w_1965));
  bfr _b_502(.a(_w_834),.q(n295_2));
  bfr _b_1540(.a(_w_1872),.q(_w_1873));
  bfr _b_681(.a(_w_1013),.q(n349));
  and_bb g176(.a(N42_0),.b(_w_2152),.q(n176));
  or_bb g170(.a(N261_2),.b(n168_0),.q(n170));
  and_bb g167(.a(N201_6),.b(n165_1),.q(n167));
  bfr _b_1045(.a(_w_1377),.q(_w_1378));
  bfr _b_521(.a(_w_853),.q(_w_854));
  bfr _b_841(.a(_w_1173),.q(_w_1174));
  and_bb g179(.a(n178),.b(n83_2),.q(_w_1104));
  or_bb g302(.a(n287_2),.b(n301),.q(n302));
  bfr _b_733(.a(_w_1065),.q(N165_2));
  or_bb g162(.a(n157),.b(n161),.q(n162));
  bfr _b_1395(.a(_w_1727),.q(_w_1728));
  bfr _b_1151(.a(_w_1483),.q(N177_2));
  bfr _b_1139(.a(_w_1471),.q(_w_1472));
  and_bb g219(.a(N237_6),.b(n211_1),.q(n219));
  bfr _b_1674(.a(_w_2006),.q(_w_2007));
  bfr _b_1530(.a(_w_1862),.q(_w_1863));
  bfr _b_1401(.a(_w_1733),.q(_w_1734));
  bfr _b_692(.a(_w_1024),.q(_w_1025));
  bfr _b_1063(.a(_w_1395),.q(_w_1396));
  and_bb g158(.a(N42_2),.b(n73_0),.q(n158));
  bfr _b_580(.a(_w_912),.q(_w_913));
  bfr _b_797(.a(_w_1129),.q(_w_1130));
  and_bb g190(.a(N116_3),.b(n162_4),.q(n190));
  bfr _b_1386(.a(_w_1718),.q(_w_1719));
  bfr _b_1244(.a(_w_1576),.q(_w_1577));
  bfr _b_873(.a(_w_1205),.q(_w_1206));
  or_bb g155(.a(n153),.b(n154),.q(n155));
  bfr _b_512(.a(_w_844),.q(_w_845));
  bfr _b_503(.a(_w_835),.q(_w_836));
  spl3L g167_s_0(.a(n167),.q0(n167_0),.q1(n167_1),.q2(n167_2));
  spl2 N219_s_0(.a(_w_2070),.q0(N219_0),.q1(_w_1119));
  and_bb g289(.a(N106_3),.b(n162_9),.q(n289));
  bfr _b_874(.a(_w_1206),.q(_w_1207));
  spl4L N116_s_0(.a(N116),.q0(N116_0),.q1(N116_1),.q2(N116_2),.q3(_w_1135));
  bfr _b_1733(.a(N17),.q(_w_2065));
  and_bi g147(.a(N1_2),.b(n146),.q(n147));
  or_bb g240(.a(n236),.b(n239),.q(_w_1826));
  and_bb g163(.a(N126_2),.b(n162_0),.q(n163));
  and_bb g65(.a(N42_7),.b(n63_0),.q(_w_1144));
  bfr _b_1145(.a(_w_1477),.q(N389));
  and_bb g151(.a(N55_2),.b(n150_0),.q(n151));
  or_bb g318(.a(n314),.b(n317),.q(_w_1176));
  bfr _b_880(.a(_w_1212),.q(_w_1213));
  bfr _b_1778(.a(_w_2110),.q(_w_2111));
  bfr _b_1130(.a(_w_1462),.q(_w_1463));
  bfr _b_890(.a(_w_1222),.q(N449));
  and_bb g312(.a(n298_2),.b(n311),.q(n312));
  spl2 N146_s_0(.a(_w_2038),.q0(N146_0),.q1(_w_1188));
  or_bb g140(.a(n138),.b(n139),.q(n140));
  spl2 g104_s_0(.a(n104),.q0(n104_0),.q1(n104_1));
  and_bi g138(.a(n137_0),.b(n128_0),.q(n138));
  bfr _b_518(.a(_w_850),.q(_w_851));
  and_bb g329(.a(N246_5),.b(n270_0),.q(n329));
  and_bb g88(.a(n83_1),.b(n87),.q(_w_1189));
  and_bi g154(.a(N42_5),.b(N17_3),.q(n154));
  and_bb g353(.a(n300_2),.b(n352_2),.q(_w_1223));
  bfr _b_1616(.a(_w_1948),.q(n194_1));
  bfr _b_794(.a(_w_1126),.q(_w_1127));
  bfr _b_1028(.a(_w_1360),.q(_w_1361));
  or_bb g200(.a(N195_6),.b(n198_3),.q(n200));
  bfr _b_1811(.a(_w_2143),.q(_w_2144));
  and_bi g95(.a(n94),.b(n93),.q(n95));
  spl2 N29_s_0(.a(N29),.q0(N29_0),.q1(N29_1));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(n140_1));
  or_bb g209(.a(n207),.b(n208),.q(n209));
  and_bb g174(.a(N237_0),.b(n167_1),.q(n174));
  bfr _b_1273(.a(_w_1605),.q(_w_1606));
  bfr _b_861(.a(_w_1193),.q(_w_1194));
  bfr _b_1762(.a(_w_2094),.q(_w_2095));
  and_bi g135(.a(n131_0),.b(n134_0),.q(n135));
  bfr _b_1430(.a(_w_1762),.q(_w_1763));
  spl2 N96_s_1(.a(N96_2),.q0(N96_3),.q1(N96_4));
  bfr _b_780(.a(_w_1112),.q(_w_1113));
  bfr _b_539(.a(_w_871),.q(_w_872));
  and_bb g250(.a(N228_2),.b(n245_2),.q(n250));
  bfr _b_853(.a(_w_1185),.q(n318));
  bfr _b_1760(.a(_w_2092),.q(_w_2093));
  bfr _b_1589(.a(_w_1921),.q(_w_1922));
  and_bb g160(.a(n159),.b(n67_1),.q(n160));
  and_bb g254(.a(N255_2),.b(_w_2130),.q(n254));
  and_bi g152(.a(n151),.b(N268_2),.q(n152));
  bfr _b_631(.a(_w_963),.q(N17_7));
  bfr _b_967(.a(_w_1299),.q(_w_1300));
  bfr _b_1613(.a(_w_1945),.q(_w_1946));
  and_bb g61(.a(N29_0),.b(N75_1),.q(_w_1224));
  or_bb g242(.a(n234),.b(n241),.q(_w_1831));
  bfr _b_957(.a(_w_1289),.q(_w_1290));
  and_bi g248(.a(n246),.b(n247),.q(n248));
  bfr _b_1617(.a(_w_1949),.q(_w_1950));
  or_bb g128(.a(n126),.b(n127),.q(n128));
  and_bb g193(.a(N189_5),.b(n192_2),.q(_w_1684));
  bfr _b_926(.a(_w_1258),.q(_w_1259));
  and_bi g127(.a(n125_1),.b(N207_1),.q(n127));
  bfr _b_1281(.a(_w_1613),.q(_w_1614));
  and_bi g311(.a(N219_7),.b(n307_0),.q(n311));
  and_bi g126(.a(N207_0),.b(n125_0),.q(n126));
  spl4L N59_s_0(.a(N59),.q0(N59_0),.q1(N59_1),.q2(N59_2),.q3(N59_3));
  spl2 N42_s_4(.a(N42_8),.q0(N42_9),.q1(N42_10));
  spl2 g131_s_0(.a(n131),.q0(n131_0),.q1(n131_1));
  spl4L g162_s_0(.a(n162),.q0(n162_0),.q1(n162_1),.q2(n162_2),.q3(n162_3));
  or_bb g226(.a(n218),.b(n225),.q(_w_1724));
  bfr _b_1531(.a(_w_1863),.q(_w_1864));
  and_bi g125(.a(n123),.b(n124),.q(n125));
  bfr _b_554(.a(_w_886),.q(_w_887));
  bfr _b_696(.a(_w_1028),.q(_w_1029));
  bfr _b_1202(.a(_w_1534),.q(_w_1535));
  bfr _b_672(.a(_w_1004),.q(n365));
  and_bb g124(.a(N189_1),.b(N195_1),.q(n124));
  spl2 N228_s_4(.a(N228_7),.q0(N228_8),.q1(_w_1235));
  or_bb g96(.a(N121_0),.b(N135_0),.q(n96));
  or_bb g123(.a(N189_0),.b(N195_0),.q(n123));
  and_bi g325(.a(N219_14),.b(n324),.q(n325));
  or_bb g166(.a(N201_5),.b(n165_0),.q(n166));
  bfr _b_959(.a(_w_1291),.q(_w_1292));
  bfr _b_1457(.a(_w_1789),.q(_w_1790));
  or_bb g122(.a(n120),.b(n121),.q(_w_1236));
  and_bb g86(.a(N59_1),.b(N68_0),.q(n86));
  and_bb g310(.a(n307_1),.b(n309),.q(n310));
  bfr _b_1123(.a(_w_1455),.q(_w_1456));
  and_bb g196(.a(N121_3),.b(n162_1),.q(n196));
  bfr _b_756(.a(_w_1088),.q(_w_1089));
  spl3L N171_s_0(.a(N171),.q0(N171_0),.q1(N171_1),.q2(_w_1238));
  and_bb g85(.a(n83_0),.b(n84),.q(_w_1246));
  or_bb g261(.a(n249),.b(n260),.q(_w_1858));
  bfr _b_1631(.a(_w_1963),.q(_w_1964));
  bfr _b_533(.a(_w_865),.q(_w_866));
  bfr _b_1529(.a(_w_1861),.q(_w_1862));
  spl2 g92_s_0(.a(n92),.q0(n92_0),.q1(n92_1));
  and_bb g340(.a(N219_13),.b(n339),.q(n340));
  bfr _b_964(.a(_w_1296),.q(_w_1297));
  or_bb g143(.a(n141),.b(n142),.q(_w_1288));
  bfr _b_1181(.a(_w_1513),.q(_w_1514));
  bfr _b_1103(.a(_w_1435),.q(_w_1436));
  and_bi g114(.a(n113_0),.b(n95_0),.q(n114));
  bfr _b_551(.a(_w_883),.q(_w_884));
  spl3L g211_s_0(.a(n211),.q0(n211_0),.q1(n211_1),.q2(_w_1316));
  and_bb g84(.a(N29_2),.b(N68_1),.q(_w_1319));
  bfr _b_668(.a(_w_1000),.q(_w_1001));
  or_bb g134(.a(n132),.b(n133),.q(n134));
  and_bb g89(.a(_w_2161),.b(n78_1),.q(_w_1322));
  bfr _b_652(.a(_w_984),.q(n70_1));
  bfr _b_1218(.a(_w_1550),.q(_w_1551));
  or_bb g285(.a(n282),.b(n284),.q(n285));
  and_bb g290(.a(N153_0),.b(n263_3),.q(n290));
  or_bb g363(.a(n359),.b(n362),.q(_w_1359));
  or_ii g76(.a(N80_4),.b(n75_0),.q(_w_1373));
  bfr _b_1271(.a(_w_1603),.q(_w_1604));
  and_bi g107(.a(n105),.b(n106),.q(n107));
  bfr _b_666(.a(_w_998),.q(n279_2));
  bfr _b_832(.a(_w_1164),.q(_w_1165));
  and_bb g62(.a(N42_9),.b(n61_1),.q(_w_1407));
  bfr _b_1695(.a(N130),.q(_w_2028));
  bfr _b_1077(.a(_w_1409),.q(_w_1410));
  or_bb g194(.a(N189_6),.b(n192_3),.q(_w_1233));
  spl2 N177_s_1(.a(N177_2),.q0(N177_3),.q1(_w_1440));
  spl2 g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1));
  and_bb g64(.a(N80_2),.b(n63_1),.q(_w_1444));
  spl4L g263_s_0(.a(n263),.q0(n263_0),.q1(n263_1),.q2(n263_2),.q3(n263_3));
  and_bb g217(.a(N219_6),.b(n216),.q(n217));
  bfr _b_1564(.a(_w_1896),.q(_w_1897));
  bfr _b_1414(.a(_w_1746),.q(_w_1747));
  and_bb g73(.a(N59_0),.b(N75_0),.q(n73));
  bfr _b_1739(.a(_w_2071),.q(_w_2072));
  bfr _b_777(.a(_w_1109),.q(_w_1110));
  bfr _b_1678(.a(_w_2010),.q(_w_2011));
  and_bb g346(.a(N165_3),.b(n179_7),.q(n346));
  spl3L N177_s_0(.a(_w_2066),.q0(N177_0),.q1(N177_1),.q2(_w_1478));
  bfr _b_593(.a(_w_925),.q(_w_926));
  bfr _b_955(.a(_w_1287),.q(N183_2));
  spl2 g61_s_0(.a(n61),.q0(n61_0),.q1(_w_1484));
  and_bb g299(.a(n296_1),.b(n298_0),.q(n299));
  and_bb g66(.a(N85),.b(N86),.q(_w_1486));
  or_bb g210(.a(n152_4),.b(n209),.q(n210));
  or_ii g74(.a(N80_3),.b(n73_1),.q(_w_1534));
  and_bb g222(.a(N106_4),.b(N210_9),.q(n222));
  bfr _b_1622(.a(_w_1954),.q(_w_1955));
  and_bb g220(.a(N246_9),.b(n210_0),.q(n220));
  bfr _b_1839(.a(N96),.q(_w_2172));
  bfr _b_1741(.a(_w_2073),.q(_w_2074));
  bfr _b_547(.a(_w_879),.q(_w_880));
  spl2 g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1));
  spl2 g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1));
  bfr _b_1165(.a(_w_1497),.q(_w_1498));
  and_bb g218(.a(N228_6),.b(n213_2),.q(n218));
  bfr _b_767(.a(_w_1099),.q(n287));
  bfr _b_751(.a(_w_1083),.q(_w_1084));
  and_bb g146(.a(N17_7),.b(n145_0),.q(n146));
  bfr _b_1608(.a(_w_1940),.q(_w_1941));
  bfr _b_1231(.a(_w_1563),.q(_w_1564));
  bfr _b_647(.a(_w_979),.q(_w_980));
  spl3L g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1),.q2(n165_2));
  bfr _b_1452(.a(_w_1784),.q(_w_1785));
  bfr _b_1051(.a(_w_1383),.q(_w_1384));
  bfr _b_1744(.a(_w_2076),.q(_w_2077));
  and_bb g63(.a(N29_3),.b(N36_0),.q(_w_1571));
  and_bb g150(.a(N447_2),.b(n149),.q(n150));
  or_ii g77(.a(N42_10),.b(n75_1),.q(_w_1572));
  bfr _b_1149(.a(_w_1481),.q(_w_1482));
  bfr _b_1086(.a(_w_1418),.q(_w_1419));
  and_bi g92(.a(n90),.b(n91),.q(n92));
  or_bb g300(.a(n295_2),.b(n299),.q(n300));
  bfr _b_1023(.a(_w_1355),.q(_w_1356));
  bfr _b_867(.a(_w_1199),.q(_w_1200));
  and_bi g103(.a(N106_1),.b(N101_1),.q(n103));
  or_bi g72(.a(N390_1),.b(n71_0),.q(N419));
  or_bb g260(.a(n250),.b(n259),.q(_w_1882));
  or_bb g101(.a(n100),.b(n99),.q(n101));
  bfr _b_1344(.a(_w_1676),.q(N850));
  or_bb g317(.a(n315),.b(n316),.q(_w_1643));
  and_bi g99(.a(N126_0),.b(n98_0),.q(n99));
  bfr _b_1727(.a(_w_2059),.q(_w_2060));
  bfr _b_595(.a(_w_927),.q(_w_928));
  bfr _b_1052(.a(_w_1384),.q(_w_1385));
  bfr _b_1645(.a(_w_1977),.q(_w_1978));
  spl3L N165_s_0(.a(N165),.q0(N165_0),.q1(N165_1),.q2(_w_1058));
  spl3L N130_s_0(.a(_w_2027),.q0(N130_0),.q1(N130_1),.q2(N130_2));
  spl2 g286_s_0(.a(n286),.q0(n286_0),.q1(n286_1));
  and_bi g208(.a(N143_1),.b(n147_2),.q(n208));
  spl2 g294_s_1(.a(n294_1),.q0(n294_2),.q1(n294_3));
  and_bi g213(.a(n212_0),.b(n211_0),.q(n213));
  and_bi g119(.a(n117),.b(n118),.q(n119));
  bfr _b_844(.a(_w_1176),.q(_w_1177));
  bfr _b_1318(.a(_w_1650),.q(_w_1651));
  spl3L g65_s_0(.a(N390_0),.q0(N390_1),.q1(N390_2),.q2(_w_1532));
  or_bb g256(.a(n254),.b(n255),.q(_w_1646));
  bfr _b_500(.a(_w_832),.q(_w_833));
  and_bb g237(.a(N111_2),.b(N210_1),.q(n237));
  spl2 g200_s_0(.a(n200),.q0(n200_0),.q1(_w_1652));
  bfr _b_1247(.a(_w_1579),.q(_w_1580));
  and_bi g356(.a(n355),.b(n353),.q(n356));
  bfr _b_944(.a(_w_1276),.q(_w_1277));
  bfr _b_970(.a(_w_1302),.q(_w_1303));
  bfr _b_1592(.a(_w_1924),.q(N153_1));
  or_bb g164(.a(n152_0),.b(n163),.q(n164));
  and_bi g113(.a(n111),.b(n112),.q(n113));
  or_bb g201(.a(N261_0),.b(n167_2),.q(n201));
  bfr _b_1498(.a(_w_1830),.q(n240));
  and_bb g249(.a(N219_2),.b(n248),.q(n249));
  bfr _b_1482(.a(_w_1814),.q(_w_1815));
  bfr _b_1203(.a(_w_1535),.q(_w_1536));
  bfr _b_607(.a(_w_939),.q(N219_14));
  spl2 N268_s_1(.a(N268_1),.q0(N268_2),.q1(_w_1654));
  bfr _b_1085(.a(_w_1417),.q(_w_1418));
  and_bb g75(.a(N36_1),.b(N59_3),.q(_w_1656));
  or_bb g108(.a(n104_0),.b(n107_0),.q(n108));
  and_bi g216(.a(n214),.b(n215),.q(n216));
  and_bi g228(.a(n194_0),.b(n193_0),.q(n228));
  or_bb g131(.a(n129),.b(n130),.q(n131));
  spl2 N29_s_1(.a(N29_1),.q0(N29_2),.q1(N29_3));
  bfr _b_842(.a(_w_1174),.q(_w_1175));
  and_bb g118(.a(N159_1),.b(N177_1),.q(n118));
  bfr _b_1265(.a(_w_1597),.q(_w_1598));
  bfr _b_1212(.a(_w_1544),.q(_w_1545));
  bfr _b_585(.a(_w_917),.q(_w_918));
  and_bb g297(.a(n206_2),.b(n212_1),.q(n297));
  or_bb g188(.a(n172),.b(n187),.q(_w_1658));
  bfr _b_1313(.a(_w_1645),.q(n317));
  or_bb g241(.a(n235),.b(n240),.q(_w_1677));
  and_bb g291(.a(N138_0),.b(_w_2054),.q(_w_1979));
  and_bb g273(.a(N96_3),.b(n162_7),.q(n273));
  or_bb g116(.a(n114),.b(n115),.q(_w_1772));
  bfr _b_553(.a(_w_885),.q(_w_886));
  and_bb g157(.a(n155),.b(n156),.q(n157));
  and_bb g331(.a(N210_6),.b(N268_3),.q(n331));
  bfr _b_772(.a(_w_1104),.q(n179));
  or_bb g268(.a(n266_0),.b(n267),.q(n268));
  bfr _b_1737(.a(_w_2069),.q(_w_2067));
  or_bb g244(.a(n232),.b(n243),.q(_w_1833));
  and_bb g199(.a(N195_5),.b(n198_2),.q(n199));
  or_bb g292(.a(n266_3),.b(n291),.q(n292));
  bfr _b_509(.a(_w_841),.q(_w_842));
  spl2 g278_s_1(.a(n278_1),.q0(n278_2),.q1(n278_3));
  and_bb g202(.a(n166_1),.b(n201),.q(n202));
  bfr _b_1175(.a(_w_1507),.q(_w_1508));
  bfr _b_660(.a(_w_992),.q(_w_993));
  or_bb g204(.a(n199_2),.b(n203),.q(n204));
  bfr _b_1532(.a(_w_1864),.q(_w_1865));
  bfr _b_1464(.a(_w_1796),.q(_w_1797));
  bfr _b_1309(.a(_w_1641),.q(_w_1642));
  spl3L N219_s_3(.a(N219_5),.q0(N219_6),.q1(N219_7),.q2(N219_8));
  and_bb g82(.a(N13_0),.b(N55_0),.q(n82));
  and_bb g301(.a(n288_1),.b(n300_0),.q(n301));
  bfr _b_943(.a(_w_1275),.q(_w_1276));
  spl4L g81_s_0(.a(N447_0),.q0(N447_1),.q1(N447_2),.q2(N447_3),.q3(_w_1605));
  or_bb g258(.a(n252),.b(n257),.q(_w_1725));
  and_bb g71(.a(n68_0),.b(n70_1),.q(_w_1727));
  bfr _b_1112(.a(_w_1444),.q(_w_1445));
  or_bb g206(.a(n193_2),.b(n205),.q(n206));
  bfr _b_594(.a(_w_926),.q(_w_927));
  and_bb g106(.a(N111_1),.b(N116_1),.q(n106));
  and_bi g115(.a(n95_1),.b(n113_1),.q(n115));
  and_bi g265(.a(N17_5),.b(N268_0),.q(_w_1118));
  and_bb g207(.a(N111_3),.b(n162_5),.q(n207));
  and_bb g360(.a(N210_8),.b(N96_4),.q(n360));
  bfr _b_769(.a(_w_1101),.q(_w_1102));
  and_bb g211(.a(N183_5),.b(n210_2),.q(n211));
  bfr _b_1358(.a(_w_1690),.q(_w_1691));
  bfr _b_706(.a(_w_1038),.q(_w_1039));
  bfr _b_1543(.a(_w_1875),.q(N865));
  spl2 g278_s_0(.a(n278),.q0(n278_0),.q1(n278_1));
  and_bb g70(.a(N1_1),.b(_w_2129),.q(n70));
  bfr _b_1435(.a(_w_1767),.q(_w_1768));
  spl2 g150_s_0(.a(n150),.q0(n150_0),.q1(n150_1));
  and_bi g133(.a(N183_1),.b(N171_1),.q(n133));
  bfr _b_1057(.a(_w_1389),.q(_w_1390));
  spl2 g288_s_0(.a(n288),.q0(n288_0),.q1(_w_1767));
  bfr _b_858(.a(_w_1190),.q(_w_1191));
  or_bb g214(.a(n206_0),.b(n213_0),.q(n214));
  bfr _b_790(.a(_w_1122),.q(_w_1123));
  and_bb g215(.a(n206_1),.b(n213_1),.q(n215));
  bfr _b_1239(.a(_w_1571),.q(n63));
  bfr _b_612(.a(_w_944),.q(_w_945));
  or_bb g225(.a(n219),.b(n224),.q(_w_1769));
  bfr _b_1056(.a(_w_1388),.q(_w_1389));
  and_bb g274(.a(N146_0),.b(n263_1),.q(n274));
  bfr _b_1819(.a(N55),.q(_w_2151));
  spl2 N268_s_0(.a(_w_2146),.q0(N268_0),.q1(_w_1770));
  bfr _b_1757(.a(_w_2089),.q(_w_2090));
  spl4L g179_s_2(.a(n179_5),.q0(n179_6),.q1(n179_7),.q2(n179_8),.q3(n179_9));
  bfr _b_905(.a(_w_1237),.q(n122));
  and_bb g345(.a(N210_7),.b(N91_4),.q(n345));
  bfr _b_1693(.a(_w_2025),.q(_w_2023));
  spl2 N36_s_0(.a(N36),.q0(_w_985),.q1(N36_1));
  and_bb g313(.a(N237_8),.b(n295_1),.q(n313));
  and_bb g156(.a(N447_3),.b(n144_1),.q(n156));
  bfr _b_1079(.a(_w_1411),.q(_w_1412));
  and_bb g221(.a(N183_3),.b(n179_9),.q(n221));
  bfr _b_1421(.a(_w_1753),.q(_w_1754));
  bfr _b_1164(.a(_w_1496),.q(_w_1497));
  bfr _b_718(.a(_w_1050),.q(_w_1051));
  or_bb g229(.a(n204_1),.b(n228_0),.q(n229));
  bfr _b_1779(.a(_w_2111),.q(_w_2112));
  or_bb g223(.a(n221),.b(n222),.q(_w_1800));
  bfr _b_609(.a(_w_941),.q(N219_12));
  bfr _b_1061(.a(_w_1393),.q(_w_1394));
  or_bb g321(.a(n310),.b(n320),.q(_w_1068));
  and_bi g161(.a(n160),.b(n158),.q(_w_1106));
  spl2 N261_s_0(.a(_w_2131),.q0(N261_0),.q1(_w_1803));
  bfr _b_928(.a(_w_1260),.q(_w_1261));
  or_bb g224(.a(n220),.b(n223),.q(_w_1804));
  bfr _b_1155(.a(_w_1487),.q(_w_1488));
  bfr _b_563(.a(_w_895),.q(_w_896));
  or_bb g192(.a(n189),.b(n191),.q(n192));
  and_bb g247(.a(n202_2),.b(n245_1),.q(n247));
  and_bi g168(.a(n166_0),.b(n167_0),.q(n168));
  or_bb g296(.a(N177_6),.b(n294_3),.q(_w_2006));
  or_bb g306(.a(n271_2),.b(n305),.q(_w_1823));
  bfr _b_1647(.a(_w_1979),.q(_w_1980));
  bfr _b_1439(.a(_w_1771),.q(N268_1));
  bfr _b_1363(.a(_w_1695),.q(_w_1696));
  bfr _b_1288(.a(_w_1620),.q(_w_1621));
  bfr _b_1091(.a(_w_1423),.q(_w_1424));
  and_bi g307(.a(n296_0),.b(n295_0),.q(n307));
  spl2 N143_s_0(.a(_w_2030),.q0(N143_0),.q1(_w_1825));
  bfr _b_1699(.a(_w_2031),.q(_w_2032));
  bfr _b_614(.a(_w_946),.q(_w_947));
  bfr _b_965(.a(_w_1297),.q(_w_1298));
  and_bb g238(.a(N255_1),.b(_w_2128),.q(n238));
  or_bb g212(.a(N183_6),.b(n210_3),.q(n212));
  spl3L g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1),.q2(n300_2));
  and_bi g231(.a(n229),.b(n230),.q(n231));
  bfr _b_1835(.a(_w_2167),.q(_w_2168));
  bfr _b_1024(.a(_w_1356),.q(_w_1357));
  bfr _b_781(.a(_w_1113),.q(_w_1114));
  bfr _b_1067(.a(_w_1399),.q(_w_1400));
  and_bb g232(.a(N219_4),.b(n231),.q(n232));
  spl2 g198_s_1(.a(n198_1),.q0(n198_2),.q1(n198_3));
  bfr _b_1801(.a(_w_2133),.q(_w_2134));
  and_bb g233(.a(N228_4),.b(n228_2),.q(n233));
  or_bb g304(.a(n279_2),.b(n303),.q(n304));
  bfr _b_1018(.a(_w_1350),.q(_w_1351));
  or_bb g243(.a(n233),.b(n242),.q(_w_1832));
  bfr _b_1830(.a(_w_2162),.q(_w_2161));
  spl4L g179_s_0(.a(n179),.q0(n179_0),.q1(n179_1),.q2(n179_2),.q3(n179_3));
  and_bb g177(.a(_w_2153),.b(n176),.q(n177));
  and_bb g112(.a(n101_1),.b(n110_1),.q(n112));
  or_bb g270(.a(n262),.b(n269),.q(n270));
  bfr _b_1682(.a(_w_2014),.q(n178));
  and_bi g308(.a(N219_9),.b(n298_1),.q(n308));
  bfr _b_731(.a(_w_1063),.q(_w_1064));
  or_bb g298(.a(n211_2),.b(n297),.q(n298));
  and_bb g315(.a(N177_3),.b(n179_4),.q(n315));
  and_bi g245(.a(n200_0),.b(n199_0),.q(n245));
  and_bi g120(.a(N130_3),.b(n119_0),.q(n120));
  and_bb g262(.a(N91_3),.b(n162_6),.q(n262));
  spl2 g270_s_0(.a(n270),.q0(n270_0),.q1(n270_1));
  bfr _b_865(.a(_w_1197),.q(_w_1198));
  and_bb g236(.a(N189_3),.b(n179_1),.q(n236));
  bfr _b_1481(.a(_w_1813),.q(_w_1814));
  and_bb g263(.a(N55_3),.b(n145_1),.q(n263));
  bfr _b_657(.a(_w_989),.q(_w_990));
  and_bi g341(.a(n340),.b(n338),.q(n341));
  bfr _b_1047(.a(_w_1379),.q(_w_1380));
  and_bb g267(.a(N138_2),.b(N8_1),.q(_w_1883));
  spl3L g83_s_0(.a(n83),.q0(n83_0),.q1(n83_1),.q2(n83_2));
  spl2 N91_s_1(.a(N91_2),.q0(N91_3),.q1(N91_4));
  spl2 N106_s_1(.a(N106_2),.q0(N106_3),.q1(N106_4));
  and_bb g109(.a(n104_1),.b(n107_1),.q(n109));
  bfr _b_1743(.a(_w_2075),.q(_w_2076));
  and_bb g275(.a(N138_3),.b(N51_3),.q(_w_1925));
  bfr _b_1346(.a(_w_1678),.q(_w_1679));
  bfr _b_906(.a(_w_1238),.q(_w_1239));
  or_bb g104(.a(n102),.b(n103),.q(n104));
  bfr _b_646(.a(_w_978),.q(n271_2));
  or_bb g278(.a(n273),.b(n277),.q(n278));
  or_bb g280(.a(N165_6),.b(n278_3),.q(_w_1932));
  bfr _b_1292(.a(_w_1624),.q(_w_1625));
  spl2 g270_s_1(.a(n270_1),.q0(n270_2),.q1(n270_3));
  bfr _b_520(.a(_w_852),.q(_w_853));
  and_bb g68(.a(N13_1),.b(N17_10),.q(n68));
  bfr _b_855(.a(_w_1187),.q(n144));
  or_bb g277(.a(n274),.b(n276),.q(n277));
  spl2 g194_s_0(.a(n194),.q0(n194_0),.q1(_w_1947));
  and_bb g69(.a(n67_2),.b(n68_1),.q(_w_1949));
  or_bb g286(.a(n281),.b(n285),.q(n286));
  spl2 N51_s_0(.a(_w_2150),.q0(N51_0),.q1(N51_1));
  bfr _b_1667(.a(_w_1999),.q(n295));
  bfr _b_950(.a(_w_1282),.q(_w_1283));
  bfr _b_973(.a(_w_1305),.q(_w_1306));
  or_bb g366(.a(n356),.b(n365),.q(_w_1986));
  bfr _b_829(.a(_w_1161),.q(_w_1162));
  spl3L g67_s_0(.a(n67),.q0(n67_0),.q1(n67_1),.q2(_w_2000));
  bfr _b_1719(.a(_w_2051),.q(_w_2052));
  bfr _b_1570(.a(_w_1902),.q(_w_1903));
  bfr _b_1060(.a(_w_1392),.q(_w_1393));
  bfr _b_1817(.a(_w_2149),.q(_w_2146));
  spl3L g298_s_0(.a(n298),.q0(n298_0),.q1(n298_1),.q2(n298_2));
  or_ii g80(.a(N390_2),.b(n71_1),.q(N446));
  bfr _b_540(.a(_w_872),.q(N228_7));
  spl2 N135_s_0(.a(N135),.q0(N135_0),.q1(N135_1));
  bfr _b_1642(.a(_w_1974),.q(_w_1975));
  and_bb g305(.a(n272_1),.b(n304_0),.q(n305));
  spl2 N261_s_1(.a(N261_1),.q0(N261_2),.q1(N261_3));
  bfr _b_1797(.a(N26),.q(_w_2129));
  bfr _b_1643(.a(_w_1975),.q(_w_1976));
  bfr _b_1416(.a(_w_1748),.q(_w_1749));
  spl2 g210_s_0(.a(n210),.q0(n210_0),.q1(_w_2015));
  or_bb g78(.a(N87),.b(N88),.q(n78));
  or_bb g309(.a(N228_8),.b(n308),.q(n309));
  bfr _b_1659(.a(_w_1991),.q(N880));
  and_bb g314(.a(N246_4),.b(n294_0),.q(n314));
  bfr _b_546(.a(_w_878),.q(_w_879));
  bfr _b_531(.a(_w_863),.q(n166_1));
  spl3L g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1),.q2(_w_2020));
  bfr _b_1195(.a(_w_1527),.q(_w_1528));
  and_bb g316(.a(N101_4),.b(N210_4),.q(n316));
  bfr _b_1527(.a(_w_1859),.q(_w_1860));
  bfr _b_1518(.a(_w_1850),.q(_w_1851));
  and_bb g282(.a(N149_0),.b(n263_2),.q(n282));
  bfr _b_542(.a(_w_874),.q(_w_875));
  bfr _b_543(.a(_w_875),.q(N159_4));
  and_bi g100(.a(n98_1),.b(N126_1),.q(n100));
  bfr _b_544(.a(_w_876),.q(_w_877));
  bfr _b_665(.a(_w_997),.q(_w_998));
  spl3L N17_s_1(.a(N17_1),.q0(N17_2),.q1(N17_3),.q2(N17_4));
  bfr _b_786(.a(_w_1118),.q(n265));
  bfr _b_545(.a(_w_877),.q(_w_878));
  bfr _b_833(.a(_w_1165),.q(_w_1166));
  bfr _b_549(.a(_w_881),.q(_w_882));
  bfr _b_917(.a(_w_1249),.q(_w_1250));
  and_bb g178(.a(n177),.b(n86_1),.q(_w_2014));
  bfr _b_550(.a(_w_882),.q(_w_883));
  and_bi g130(.a(N165_1),.b(N201_1),.q(n130));
  bfr _b_552(.a(_w_884),.q(_w_885));
  and_bb g180(.a(N201_3),.b(n179_0),.q(n180));
  bfr _b_899(.a(_w_1231),.q(_w_1232));
  spl2 N228_s_2(.a(N228_3),.q0(N228_4),.q1(_w_1682));
  bfr _b_555(.a(_w_887),.q(_w_888));
  bfr _b_1502(.a(_w_1834),.q(_w_1835));
  bfr _b_557(.a(_w_889),.q(N111_3));
  bfr _b_558(.a(_w_890),.q(_w_891));
  bfr _b_559(.a(_w_891),.q(_w_892));
  bfr _b_1770(.a(_w_2102),.q(_w_2087));
  spl2 N201_s_2(.a(N201_4),.q0(N201_5),.q1(N201_6));
  bfr _b_560(.a(_w_892),.q(n287_2));
  bfr _b_1365(.a(_w_1697),.q(_w_1698));
  bfr _b_685(.a(_w_1017),.q(_w_1018));
  bfr _b_1676(.a(_w_2008),.q(_w_2009));
  bfr _b_1448(.a(_w_1780),.q(_w_1781));
  bfr _b_766(.a(_w_1098),.q(_w_1099));
  bfr _b_896(.a(_w_1228),.q(_w_1229));
  bfr _b_1684(.a(_w_2016),.q(_w_2017));
  bfr _b_564(.a(_w_896),.q(_w_897));
  bfr _b_565(.a(_w_897),.q(_w_898));
  and_bb g175(.a(N246_2),.b(n165_2),.q(n175));
  bfr _b_599(.a(_w_931),.q(_w_932));
  bfr _b_567(.a(_w_899),.q(_w_900));
  bfr _b_590(.a(_w_922),.q(_w_923));
  and_bb g91(.a(N130_1),.b(N96_1),.q(n91));
  bfr _b_568(.a(_w_900),.q(_w_901));
  bfr _b_1534(.a(_w_1866),.q(_w_1867));
  bfr _b_569(.a(_w_901),.q(_w_902));
  bfr _b_1000(.a(_w_1332),.q(_w_1333));
  bfr _b_570(.a(_w_902),.q(N138_4));
  bfr _b_988(.a(_w_1320),.q(n84));
  bfr _b_571(.a(_w_903),.q(_w_904));
  bfr _b_572(.a(_w_904),.q(_w_905));
  spl3L g271_s_0(.a(n271),.q0(n271_0),.q1(n271_1),.q2(_w_976));
  bfr _b_984(.a(_w_1316),.q(_w_1317));
  bfr _b_573(.a(_w_905),.q(N165_4));
  bfr _b_1477(.a(_w_1809),.q(_w_1810));
  bfr _b_1385(.a(_w_1717),.q(_w_1718));
  bfr _b_659(.a(_w_991),.q(_w_992));
  and_bb g144(.a(_w_2063),.b(N59_2),.q(_w_1186));
  bfr _b_574(.a(_w_906),.q(_w_907));
  bfr _b_1704(.a(_w_2036),.q(_w_2037));
  bfr _b_575(.a(_w_907),.q(N8_1));
  bfr _b_1776(.a(_w_2108),.q(_w_2109));
  bfr _b_1116(.a(_w_1448),.q(_w_1449));
  bfr _b_576(.a(_w_908),.q(_w_909));
  and_bb g303(.a(n280_1),.b(n302_0),.q(n303));
  bfr _b_709(.a(_w_1041),.q(_w_1042));
  bfr _b_1661(.a(_w_1993),.q(_w_1994));
  bfr _b_578(.a(_w_910),.q(_w_911));
  bfr _b_581(.a(_w_913),.q(_w_914));
  bfr _b_640(.a(_w_972),.q(_w_973));
  bfr _b_886(.a(_w_1218),.q(_w_1219));
  bfr _b_583(.a(_w_915),.q(N121_3));
  bfr _b_651(.a(_w_983),.q(_w_984));
  bfr _b_697(.a(_w_1029),.q(_w_1030));
  bfr _b_584(.a(_w_916),.q(_w_917));
  bfr _b_1588(.a(_w_1920),.q(_w_1921));
  bfr _b_588(.a(_w_920),.q(_w_921));
  bfr _b_591(.a(_w_923),.q(_w_924));
  bfr _b_641(.a(_w_973),.q(N96_2));
  bfr _b_592(.a(_w_924),.q(N183_4));
  bfr _b_596(.a(_w_928),.q(_w_929));
  bfr _b_1755(.a(N228),.q(_w_2088));
  bfr _b_597(.a(_w_929),.q(_w_930));
  bfr _b_606(.a(_w_938),.q(_w_939));
  bfr _b_882(.a(_w_1214),.q(_w_1215));
  and_bb g255(.a(N116_2),.b(N210_2),.q(n255));
  bfr _b_598(.a(_w_930),.q(N189_4));
  bfr _b_1142(.a(_w_1474),.q(_w_1475));
  bfr _b_600(.a(_w_932),.q(_w_933));
  bfr _b_603(.a(_w_935),.q(_w_936));
  bfr _b_1135(.a(_w_1467),.q(_w_1468));
  spl2 g86_s_0(.a(n86),.q0(n86_0),.q1(n86_1));
  bfr _b_700(.a(_w_1032),.q(n347));
  bfr _b_604(.a(_w_936),.q(N189_2));
  bfr _b_610(.a(_w_942),.q(_w_943));
  bfr _b_773(.a(_w_1105),.q(n185));
  bfr _b_611(.a(_w_943),.q(N228_3));
  bfr _b_1258(.a(_w_1590),.q(_w_1591));
  bfr _b_613(.a(_w_945),.q(N219_5));
  bfr _b_617(.a(_w_949),.q(_w_950));
  bfr _b_618(.a(_w_950),.q(N237_11));
  bfr _b_1037(.a(_w_1369),.q(_w_1370));
  bfr _b_622(.a(_w_954),.q(_w_955));
  bfr _b_796(.a(_w_1128),.q(_w_1129));
  bfr _b_1425(.a(_w_1757),.q(_w_1758));
  or_bb g339(.a(n302_1),.b(n337_0),.q(n339));
  bfr _b_623(.a(_w_955),.q(N237_3));
  bfr _b_680(.a(_w_1012),.q(n350));
  bfr _b_1046(.a(_w_1378),.q(_w_1379));
  bfr _b_624(.a(_w_956),.q(_w_957));
  bfr _b_814(.a(_w_1146),.q(_w_1147));
  bfr _b_626(.a(_w_958),.q(_w_959));
  bfr _b_1509(.a(_w_1841),.q(_w_1842));
  bfr _b_632(.a(_w_964),.q(n75_1));
  bfr _b_875(.a(_w_1207),.q(_w_1208));
  bfr _b_627(.a(_w_959),.q(N55_1));
  or_bb g259(.a(n251),.b(n258),.q(_w_1640));
  and_bb g344(.a(N246_6),.b(n278_0),.q(n344));
  bfr _b_628(.a(_w_960),.q(N68_1));
  bfr _b_1569(.a(_w_1901),.q(_w_1902));
  bfr _b_747(.a(_w_1079),.q(n319));
  bfr _b_1731(.a(N156),.q(_w_2063));
  or_bb g348(.a(n344),.b(n347),.q(_w_1014));
  and_bi g153(.a(N17_2),.b(N42_4),.q(n153));
  bfr _b_876(.a(_w_1208),.q(_w_1209));
  bfr _b_629(.a(_w_961),.q(_w_962));
  bfr _b_630(.a(_w_962),.q(N91_2));
  bfr _b_1510(.a(_w_1842),.q(_w_1843));
  bfr _b_633(.a(_w_965),.q(_w_966));
  bfr _b_634(.a(_w_966),.q(_w_967));
  bfr _b_675(.a(_w_1007),.q(_w_1008));
  bfr _b_1802(.a(_w_2134),.q(_w_2135));
  bfr _b_1538(.a(_w_1870),.q(_w_1871));
  bfr _b_868(.a(_w_1200),.q(_w_1201));
  bfr _b_635(.a(_w_967),.q(N228_13));
  spl3L g202_s_0(.a(n202),.q0(n202_0),.q1(n202_1),.q2(n202_2));
  bfr _b_636(.a(_w_968),.q(N42_1));
  bfr _b_1286(.a(_w_1618),.q(_w_1619));
  bfr _b_638(.a(_w_970),.q(_w_971));
  bfr _b_620(.a(_w_952),.q(_w_953));
  bfr _b_1020(.a(_w_1352),.q(_w_1353));
  bfr _b_642(.a(_w_974),.q(_w_975));
  spl3L g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1),.q2(n304_2));
  bfr _b_644(.a(_w_976),.q(_w_977));
  bfr _b_1066(.a(_w_1398),.q(_w_1399));
  bfr _b_648(.a(_w_980),.q(_w_981));
  and_bb g79(.a(_w_2163),.b(n78_0),.q(_w_1686));
  bfr _b_768(.a(_w_1100),.q(_w_1101));
  bfr _b_682(.a(_w_1014),.q(_w_1015));
  and_bi g172(.a(n171),.b(n169),.q(n172));
  bfr _b_938(.a(_w_1270),.q(_w_1271));
  bfr _b_653(.a(_w_985),.q(N36_0));
  bfr _b_654(.a(_w_986),.q(N101_3));
  spl3L N80_s_1(.a(N80_1),.q0(N80_2),.q1(N80_3),.q2(N80_4));
  bfr _b_1044(.a(_w_1376),.q(_w_1377));
  bfr _b_662(.a(_w_994),.q(_w_995));
  bfr _b_663(.a(_w_995),.q(n272_1));
  bfr _b_1446(.a(_w_1778),.q(_w_1779));
  bfr _b_664(.a(_w_996),.q(_w_997));
  bfr _b_686(.a(_w_1018),.q(_w_1019));
  bfr _b_1685(.a(_w_2017),.q(_w_2018));
  bfr _b_979(.a(_w_1311),.q(_w_1312));
  bfr _b_1225(.a(_w_1557),.q(_w_1558));
  bfr _b_669(.a(_w_1001),.q(n296_1));
  bfr _b_1096(.a(_w_1428),.q(_w_1429));
  bfr _b_670(.a(_w_1002),.q(_w_1003));
  bfr _b_729(.a(_w_1061),.q(_w_1062));
  bfr _b_673(.a(_w_1005),.q(n364));
  bfr _b_619(.a(_w_951),.q(N237_7));
  bfr _b_839(.a(_w_1171),.q(_w_1172));
  bfr _b_501(.a(_w_833),.q(_w_834));
  bfr _b_661(.a(_w_993),.q(N101_2));
  bfr _b_676(.a(_w_1008),.q(n307_1));
  bfr _b_678(.a(_w_1010),.q(_w_1011));
  bfr _b_679(.a(_w_1011),.q(N879));
  bfr _b_1019(.a(_w_1351),.q(_w_1352));
  bfr _b_683(.a(_w_1015),.q(_w_1016));
  or_bb g198(.a(n195),.b(n197),.q(n198));
  bfr _b_688(.a(_w_1020),.q(_w_1021));
  bfr _b_689(.a(_w_1021),.q(_w_1022));
  bfr _b_691(.a(_w_1023),.q(_w_1024));
  bfr _b_694(.a(_w_1026),.q(_w_1027));
  bfr _b_698(.a(_w_1030),.q(n348));
  spl2 N8_s_0(.a(N8),.q0(N8_0),.q1(_w_906));
  bfr _b_699(.a(_w_1031),.q(_w_1032));
  bfr _b_1436(.a(_w_1768),.q(n288_1));
  bfr _b_701(.a(_w_1033),.q(n338));
  bfr _b_784(.a(_w_1116),.q(_w_1117));
  bfr _b_702(.a(_w_1034),.q(n335));
  bfr _b_703(.a(_w_1035),.q(n334));
  bfr _b_744(.a(_w_1076),.q(N874));
  bfr _b_1367(.a(_w_1699),.q(_w_1700));
  spl3L N1_s_0(.a(N1),.q0(N1_0),.q1(N1_1),.q2(_w_1111));
  bfr _b_704(.a(_w_1036),.q(_w_1037));
  bfr _b_1772(.a(_w_2104),.q(_w_2105));
  bfr _b_1326(.a(_w_1658),.q(_w_1659));
  bfr _b_556(.a(_w_888),.q(_w_889));
  bfr _b_1005(.a(_w_1337),.q(_w_1338));
  and_bb g230(.a(n204_2),.b(n228_1),.q(n230));
  bfr _b_707(.a(_w_1039),.q(_w_1040));
  bfr _b_996(.a(_w_1328),.q(_w_1329));
  bfr _b_708(.a(_w_1040),.q(_w_1041));
  bfr _b_893(.a(_w_1225),.q(n187));
  bfr _b_710(.a(_w_1042),.q(_w_1043));
  bfr _b_711(.a(_w_1043),.q(_w_1044));
  bfr _b_714(.a(_w_1046),.q(_w_1047));
  bfr _b_715(.a(_w_1047),.q(_w_1048));
  bfr _b_919(.a(_w_1251),.q(_w_1252));
  bfr _b_1653(.a(_w_1985),.q(n291));
  and_bi g148(.a(N153_1),.b(n147_0),.q(n148));
  bfr _b_639(.a(_w_971),.q(_w_972));
  bfr _b_720(.a(_w_1052),.q(_w_1053));
  bfr _b_721(.a(_w_1053),.q(_w_1054));
  spl2 g296_s_0(.a(n296),.q0(n296_0),.q1(_w_999));
  bfr _b_1049(.a(_w_1381),.q(_w_1382));
  bfr _b_615(.a(_w_947),.q(_w_948));
  bfr _b_722(.a(_w_1054),.q(_w_1055));
  bfr _b_831(.a(_w_1163),.q(_w_1164));
  bfr _b_1008(.a(_w_1340),.q(_w_1341));
  bfr _b_723(.a(_w_1055),.q(n333));
  bfr _b_724(.a(_w_1056),.q(_w_1057));
  bfr _b_1054(.a(_w_1386),.q(_w_1387));
  and_bb g159(.a(N17_0),.b(N51_0),.q(n159));
  bfr _b_1022(.a(_w_1354),.q(_w_1355));
  bfr _b_725(.a(_w_1057),.q(n332));
  bfr _b_1494(.a(_w_1826),.q(_w_1827));
  bfr _b_1238(.a(_w_1570),.q(N171_4));
  bfr _b_582(.a(_w_914),.q(_w_915));
  bfr _b_727(.a(_w_1059),.q(_w_1060));
  bfr _b_1390(.a(_w_1722),.q(N423));
  spl2 g107_s_0(.a(n107),.q0(n107_0),.q1(n107_1));
  bfr _b_728(.a(_w_1060),.q(_w_1061));
  bfr _b_734(.a(_w_1066),.q(N138_1));
  bfr _b_884(.a(_w_1216),.q(_w_1217));
  and_bi g189(.a(N146_1),.b(n147_3),.q(_w_1681));
  bfr _b_677(.a(_w_1009),.q(_w_1010));
  bfr _b_735(.a(_w_1067),.q(n323));
  and_bb g235(.a(N246_10),.b(n192_0),.q(n235));
  and_bb g149(.a(N80_0),.b(n61_0),.q(n149));
  bfr _b_738(.a(_w_1070),.q(_w_1071));
  bfr _b_739(.a(_w_1071),.q(_w_1072));
  bfr _b_740(.a(_w_1072),.q(_w_1073));
  bfr _b_1780(.a(_w_2112),.q(_w_2113));
  bfr _b_1097(.a(_w_1429),.q(_w_1430));
  bfr _b_783(.a(_w_1115),.q(_w_1116));
  bfr _b_732(.a(_w_1064),.q(_w_1065));
  bfr _b_743(.a(_w_1075),.q(_w_1076));
  and_bi g136(.a(n134_1),.b(n131_1),.q(n136));
  bfr _b_808(.a(_w_1140),.q(_w_1141));
  bfr _b_746(.a(_w_1078),.q(_w_1079));
  bfr _b_749(.a(_w_1081),.q(_w_1082));
  bfr _b_939(.a(_w_1271),.q(_w_1272));
  spl3L g204_s_0(.a(n204),.q0(n204_0),.q1(n204_1),.q2(n204_2));
  bfr _b_752(.a(_w_1084),.q(_w_1085));
  bfr _b_753(.a(_w_1085),.q(_w_1086));
  bfr _b_779(.a(_w_1111),.q(_w_1112));
  bfr _b_754(.a(_w_1086),.q(n184));
  bfr _b_1009(.a(_w_1341),.q(_w_1342));
  bfr _b_817(.a(_w_1149),.q(_w_1150));
  bfr _b_755(.a(_w_1087),.q(n186));
  bfr _b_757(.a(_w_1089),.q(_w_1090));
  bfr _b_927(.a(_w_1259),.q(_w_1260));
  bfr _b_758(.a(_w_1090),.q(_w_1091));
  and_bb g357(.a(N228_10),.b(n352_1),.q(n357));
  bfr _b_759(.a(_w_1091),.q(_w_1092));
  bfr _b_922(.a(_w_1254),.q(_w_1255));
  bfr _b_760(.a(_w_1092),.q(_w_1093));
  bfr _b_924(.a(_w_1256),.q(_w_1257));
  bfr _b_975(.a(_w_1307),.q(_w_1308));
  bfr _b_761(.a(_w_1093),.q(_w_1094));
  bfr _b_762(.a(_w_1094),.q(_w_1095));
  bfr _b_763(.a(_w_1095),.q(_w_1096));
  and_bi g142(.a(n140_1),.b(n122_1),.q(n142));
  bfr _b_764(.a(_w_1096),.q(_w_1097));
  bfr _b_1102(.a(_w_1434),.q(_w_1435));
  bfr _b_1729(.a(_w_2061),.q(_w_2062));
  and_bi g145(.a(N447_1),.b(n144_0),.q(n145));
  bfr _b_625(.a(_w_957),.q(_w_958));
  bfr _b_774(.a(_w_1106),.q(_w_1107));
  bfr _b_775(.a(_w_1107),.q(n161));
  bfr _b_852(.a(_w_1184),.q(_w_1185));
  bfr _b_776(.a(_w_1108),.q(_w_1109));
  bfr _b_1016(.a(_w_1348),.q(_w_1349));
  bfr _b_1547(.a(_w_1879),.q(_w_1880));
  bfr _b_778(.a(_w_1110),.q(N237_9));
  bfr _b_787(.a(_w_1119),.q(N219_1));
  bfr _b_788(.a(_w_1120),.q(_w_1121));
  bfr _b_791(.a(_w_1123),.q(_w_1124));
  bfr _b_771(.a(_w_1103),.q(n257));
  bfr _b_792(.a(_w_1124),.q(_w_1125));
  bfr _b_793(.a(_w_1125),.q(_w_1126));
  bfr _b_798(.a(_w_1130),.q(_w_1131));
  bfr _b_799(.a(_w_1131),.q(_w_1132));
  bfr _b_1505(.a(_w_1837),.q(_w_1838));
  bfr _b_947(.a(_w_1279),.q(N448));
  bfr _b_977(.a(_w_1309),.q(_w_1310));
  bfr _b_801(.a(_w_1133),.q(_w_1134));
  bfr _b_802(.a(_w_1134),.q(n279));
  bfr _b_1766(.a(_w_2098),.q(_w_2099));
  bfr _b_952(.a(_w_1284),.q(_w_1285));
  bfr _b_1712(.a(_w_2044),.q(_w_2045));
  bfr _b_803(.a(_w_1135),.q(_w_1136));
  bfr _b_804(.a(_w_1136),.q(_w_1137));
  bfr _b_1027(.a(_w_1359),.q(_w_1360));
  bfr _b_806(.a(_w_1138),.q(_w_1139));
  bfr _b_807(.a(_w_1139),.q(_w_1140));
  bfr _b_809(.a(_w_1141),.q(_w_1142));
  bfr _b_1308(.a(_w_1640),.q(n259));
  bfr _b_810(.a(_w_1142),.q(_w_1143));
  bfr _b_811(.a(_w_1143),.q(N116_3));
  bfr _b_826(.a(_w_1158),.q(_w_1159));
  bfr _b_812(.a(_w_1144),.q(_w_1145));
  bfr _b_813(.a(_w_1145),.q(_w_1146));
  bfr _b_1511(.a(_w_1843),.q(_w_1844));
  bfr _b_506(.a(_w_838),.q(_w_839));
  bfr _b_816(.a(_w_1148),.q(_w_1149));
  bfr _b_823(.a(_w_1155),.q(_w_1156));
  bfr _b_824(.a(_w_1156),.q(_w_1157));
  bfr _b_825(.a(_w_1157),.q(_w_1158));
  bfr _b_827(.a(_w_1159),.q(_w_1160));
  bfr _b_1828(.a(_w_2160),.q(_w_2158));
  and_bi g98(.a(n96),.b(n97),.q(n98));
  bfr _b_649(.a(_w_981),.q(_w_982));
  bfr _b_828(.a(_w_1160),.q(_w_1161));
  bfr _b_953(.a(_w_1285),.q(_w_1286));
  bfr _b_830(.a(_w_1162),.q(_w_1163));
  bfr _b_742(.a(_w_1074),.q(_w_1075));
  bfr _b_935(.a(_w_1267),.q(_w_1268));
  bfr _b_674(.a(_w_1006),.q(_w_1007));
  bfr _b_834(.a(_w_1166),.q(_w_1167));
  bfr _b_1208(.a(_w_1540),.q(_w_1541));
  or_bb g351(.a(n341),.b(n350),.q(_w_1009));
  bfr _b_835(.a(_w_1167),.q(_w_1168));
  bfr _b_836(.a(_w_1168),.q(_w_1169));
  bfr _b_1602(.a(_w_1934),.q(_w_1935));
  bfr _b_837(.a(_w_1169),.q(_w_1170));
  bfr _b_846(.a(_w_1178),.q(_w_1179));
  bfr _b_968(.a(_w_1300),.q(_w_1301));
  spl2 g68_s_0(.a(n68),.q0(n68_0),.q1(n68_1));
  bfr _b_838(.a(_w_1170),.q(_w_1171));
  bfr _b_991(.a(_w_1323),.q(_w_1324));
  bfr _b_840(.a(_w_1172),.q(_w_1173));
  bfr _b_845(.a(_w_1177),.q(_w_1178));
  and_bb g181(.a(N255_0),.b(_w_2145),.q(n181));
  bfr _b_645(.a(_w_977),.q(_w_978));
  bfr _b_667(.a(_w_999),.q(_w_1000));
  bfr _b_847(.a(_w_1179),.q(_w_1180));
  bfr _b_1840(.a(_w_2172),.q(_w_2173));
  bfr _b_850(.a(_w_1182),.q(_w_1183));
  bfr _b_851(.a(_w_1183),.q(_w_1184));
  bfr _b_1791(.a(_w_2123),.q(_w_2124));
  bfr _b_849(.a(_w_1181),.q(_w_1182));
  bfr _b_856(.a(_w_1188),.q(N146_1));
  bfr _b_1029(.a(_w_1361),.q(_w_1362));
  bfr _b_857(.a(_w_1189),.q(_w_1190));
  bfr _b_1581(.a(_w_1913),.q(_w_1914));
  and_bi g132(.a(N171_0),.b(N183_0),.q(n132));
  bfr _b_859(.a(_w_1191),.q(_w_1192));
  spl2 N219_s_1(.a(N219_1),.q0(N219_2),.q1(_w_1930));
  bfr _b_860(.a(_w_1192),.q(_w_1193));
  bfr _b_862(.a(_w_1194),.q(_w_1195));
  bfr _b_1619(.a(_w_1951),.q(_w_1952));
  bfr _b_864(.a(_w_1196),.q(_w_1197));
  bfr _b_693(.a(_w_1025),.q(_w_1026));
  bfr _b_1069(.a(_w_1401),.q(_w_1402));
  bfr _b_866(.a(_w_1198),.q(_w_1199));
  or_bb g293(.a(n290),.b(n292),.q(n293));
  bfr _b_869(.a(_w_1201),.q(_w_1202));
  spl2 N237_s_6(.a(N237_11),.q0(N237_12),.q1(_w_946));
  bfr _b_870(.a(_w_1202),.q(_w_1203));
  bfr _b_1508(.a(_w_1840),.q(_w_1841));
  bfr _b_871(.a(_w_1203),.q(_w_1204));
  bfr _b_1261(.a(_w_1593),.q(_w_1594));
  bfr _b_872(.a(_w_1204),.q(_w_1205));
  bfr _b_1478(.a(_w_1810),.q(n224));
  bfr _b_877(.a(_w_1209),.q(_w_1210));
  bfr _b_719(.a(_w_1051),.q(_w_1052));
  bfr _b_878(.a(_w_1210),.q(_w_1211));
  bfr _b_879(.a(_w_1211),.q(_w_1212));
  bfr _b_883(.a(_w_1215),.q(_w_1216));
  bfr _b_885(.a(_w_1217),.q(_w_1218));
  bfr _b_887(.a(_w_1219),.q(_w_1220));
  bfr _b_888(.a(_w_1220),.q(_w_1221));
  bfr _b_1031(.a(_w_1363),.q(_w_1364));
  bfr _b_1400(.a(_w_1732),.q(_w_1733));
  bfr _b_671(.a(_w_1003),.q(n212_1));
  bfr _b_891(.a(_w_1223),.q(n353));
  bfr _b_1383(.a(_w_1715),.q(_w_1716));
  and_bb g87(.a(_w_2155),.b(n86_0),.q(_w_1321));
  bfr _b_892(.a(_w_1224),.q(n61));
  bfr _b_925(.a(_w_1257),.q(_w_1258));
  bfr _b_1003(.a(_w_1335),.q(_w_1336));
  spl3L g322_s_0(.a(n322),.q0(n322_0),.q1(n322_1),.q2(n322_2));
  bfr _b_894(.a(_w_1226),.q(_w_1227));
  bfr _b_1469(.a(_w_1801),.q(_w_1802));
  bfr _b_534(.a(_w_866),.q(n193_2));
  bfr _b_705(.a(_w_1037),.q(_w_1038));
  bfr _b_895(.a(_w_1227),.q(_w_1228));
  bfr _b_897(.a(_w_1229),.q(_w_1230));
  bfr _b_901(.a(_w_1233),.q(_w_1234));
  bfr _b_1315(.a(_w_1647),.q(_w_1648));
  bfr _b_902(.a(_w_1234),.q(n194));
  bfr _b_1644(.a(_w_1976),.q(_w_1977));
  spl2 N42_s_1(.a(N42_1),.q0(N42_2),.q1(N42_3));
  and_bb g81(.a(N51_2),.b(n70_0),.q(N447_0));
  bfr _b_903(.a(_w_1235),.q(N228_9));
  bfr _b_601(.a(_w_933),.q(_w_934));
  bfr _b_904(.a(_w_1236),.q(_w_1237));
  spl3L g193_s_0(.a(n193),.q0(n193_0),.q1(n193_1),.q2(_w_864));
  bfr _b_907(.a(_w_1239),.q(_w_1240));
  bfr _b_908(.a(_w_1240),.q(_w_1241));
  or_bb g227(.a(n217),.b(n226),.q(_w_1811));
  bfr _b_1100(.a(_w_1432),.q(_w_1433));
  bfr _b_889(.a(_w_1221),.q(_w_1222));
  bfr _b_909(.a(_w_1241),.q(_w_1242));
  bfr _b_1105(.a(_w_1437),.q(_w_1438));
  bfr _b_911(.a(_w_1243),.q(_w_1244));
  and_bb g266(.a(n150_1),.b(n265),.q(n266));
  bfr _b_913(.a(_w_1245),.q(N171_2));
  bfr _b_684(.a(_w_1016),.q(_w_1017));
  or_bb g117(.a(N159_0),.b(N177_0),.q(n117));
  bfr _b_912(.a(_w_1244),.q(_w_1245));
  bfr _b_914(.a(_w_1246),.q(_w_1247));
  bfr _b_918(.a(_w_1250),.q(_w_1251));
  bfr _b_920(.a(_w_1252),.q(_w_1253));
  and_bb g279(.a(N165_5),.b(n278_2),.q(_w_1120));
  bfr _b_921(.a(_w_1253),.q(_w_1254));
  bfr _b_923(.a(_w_1255),.q(_w_1256));
  bfr _b_1182(.a(_w_1514),.q(_w_1515));
  bfr _b_929(.a(_w_1261),.q(_w_1262));
  bfr _b_717(.a(_w_1049),.q(_w_1050));
  bfr _b_930(.a(_w_1262),.q(_w_1263));
  bfr _b_1492(.a(_w_1824),.q(N866));
  bfr _b_1392(.a(_w_1724),.q(n226));
  or_bb g323(.a(n304_2),.b(n322_2),.q(_w_1067));
  spl3L N183_s_0(.a(N183),.q0(N183_0),.q1(N183_1),.q2(_w_1280));
  bfr _b_566(.a(_w_898),.q(N126_2));
  bfr _b_931(.a(_w_1263),.q(_w_1264));
  bfr _b_933(.a(_w_1265),.q(_w_1266));
  or_bb g94(.a(N91_1),.b(n92_1),.q(n94));
  bfr _b_848(.a(_w_1180),.q(_w_1181));
  bfr _b_1006(.a(_w_1338),.q(_w_1339));
  bfr _b_519(.a(_w_851),.q(_w_852));
  bfr _b_937(.a(_w_1269),.q(_w_1270));
  bfr _b_1668(.a(_w_2000),.q(_w_2001));
  bfr _b_941(.a(_w_1273),.q(_w_1274));
  bfr _b_1636(.a(_w_1968),.q(_w_1969));
  bfr _b_1415(.a(_w_1747),.q(_w_1748));
  bfr _b_942(.a(_w_1274),.q(_w_1275));
  bfr _b_945(.a(_w_1277),.q(_w_1278));
  bfr _b_1382(.a(_w_1714),.q(_w_1715));
  bfr _b_948(.a(_w_1280),.q(_w_1281));
  bfr _b_526(.a(_w_858),.q(_w_859));
  bfr _b_949(.a(_w_1281),.q(_w_1282));
  bfr _b_951(.a(_w_1283),.q(_w_1284));
  bfr _b_1015(.a(_w_1347),.q(_w_1348));
  bfr _b_956(.a(_w_1288),.q(_w_1289));
  bfr _b_958(.a(_w_1290),.q(_w_1291));
  bfr _b_1209(.a(_w_1541),.q(_w_1542));
  bfr _b_960(.a(_w_1292),.q(_w_1293));
  bfr _b_961(.a(_w_1293),.q(_w_1294));
  bfr _b_1353(.a(_w_1685),.q(n193));
  bfr _b_548(.a(_w_880),.q(N13_1));
  bfr _b_962(.a(_w_1294),.q(_w_1295));
  bfr _b_963(.a(_w_1295),.q(_w_1296));
  and_bb g205(.a(n194_1),.b(n204_0),.q(n205));
  bfr _b_971(.a(_w_1303),.q(_w_1304));
  bfr _b_966(.a(_w_1298),.q(_w_1299));
  bfr _b_910(.a(_w_1242),.q(_w_1243));
  bfr _b_741(.a(_w_1073),.q(_w_1074));
  bfr _b_972(.a(_w_1304),.q(_w_1305));
  bfr _b_1753(.a(_w_2085),.q(_w_2086));
  bfr _b_1284(.a(_w_1616),.q(_w_1617));
  bfr _b_1252(.a(_w_1584),.q(_w_1585));
  bfr _b_974(.a(_w_1306),.q(_w_1307));
  bfr _b_976(.a(_w_1308),.q(_w_1309));
  bfr _b_980(.a(_w_1312),.q(_w_1313));
  bfr _b_1800(.a(_w_2132),.q(_w_2133));
  bfr _b_982(.a(_w_1314),.q(_w_1315));
  bfr _b_1726(.a(_w_2058),.q(_w_2059));
  bfr _b_983(.a(_w_1315),.q(N768));
  bfr _b_1197(.a(_w_1529),.q(_w_1530));
  or_bb g362(.a(n360),.b(n361),.q(_w_1641));
  bfr _b_985(.a(_w_1317),.q(_w_1318));
  bfr _b_736(.a(_w_1068),.q(_w_1069));
  bfr _b_987(.a(_w_1319),.q(_w_1320));
  spl2 N101_s_1(.a(N101_2),.q0(_w_986),.q1(N101_4));
  bfr _b_989(.a(_w_1321),.q(n87));
  bfr _b_990(.a(_w_1322),.q(_w_1323));
  bfr _b_992(.a(_w_1324),.q(_w_1325));
  bfr _b_993(.a(_w_1325),.q(_w_1326));
  spl2 N228_s_5(.a(N228_9),.q0(N228_10),.q1(_w_868));
  bfr _b_1001(.a(_w_1333),.q(_w_1334));
  bfr _b_994(.a(_w_1326),.q(_w_1327));
  bfr _b_995(.a(_w_1327),.q(_w_1328));
  bfr _b_997(.a(_w_1329),.q(_w_1330));
  bfr _b_998(.a(_w_1330),.q(_w_1331));
  spl2 g113_s_0(.a(n113),.q0(n113_0),.q1(n113_1));
  or_bb g165(.a(n148),.b(n164),.q(n165));
  bfr _b_999(.a(_w_1331),.q(_w_1332));
  bfr _b_1002(.a(_w_1334),.q(_w_1335));
  spl3L N138_s_1(.a(N138_1),.q0(N138_2),.q1(N138_3),.q2(_w_899));
  bfr _b_1004(.a(_w_1336),.q(_w_1337));
  bfr _b_1007(.a(_w_1339),.q(_w_1340));
  bfr _b_1010(.a(_w_1342),.q(_w_1343));
  bfr _b_986(.a(_w_1318),.q(n211_2));
  bfr _b_1011(.a(_w_1343),.q(_w_1344));
  bfr _b_1013(.a(_w_1345),.q(_w_1346));
  bfr _b_1486(.a(_w_1818),.q(_w_1819));
  bfr _b_1014(.a(_w_1346),.q(_w_1347));
  bfr _b_1331(.a(_w_1663),.q(_w_1664));
  or_bb g239(.a(n237),.b(n238),.q(_w_1525));
  bfr _b_946(.a(_w_1278),.q(_w_1279));
  bfr _b_1017(.a(_w_1349),.q(_w_1350));
  bfr _b_1021(.a(_w_1353),.q(_w_1354));
  bfr _b_863(.a(_w_1195),.q(_w_1196));
  bfr _b_726(.a(_w_1058),.q(_w_1059));
  bfr _b_579(.a(_w_911),.q(_w_912));
  bfr _b_1025(.a(_w_1357),.q(_w_1358));
  or_bb g284(.a(n266_2),.b(n283),.q(n284));
  bfr _b_1032(.a(_w_1364),.q(_w_1365));
  bfr _b_1033(.a(_w_1365),.q(_w_1366));
  bfr _b_1034(.a(_w_1366),.q(_w_1367));
  bfr _b_1035(.a(_w_1367),.q(_w_1368));
  bfr _b_1036(.a(_w_1368),.q(_w_1369));
  bfr _b_1285(.a(_w_1617),.q(_w_1618));
  bfr _b_687(.a(_w_1019),.q(_w_1020));
  bfr _b_1038(.a(_w_1370),.q(_w_1371));
  spl2 N17_s_0(.a(_w_2065),.q0(N17_0),.q1(_w_1723));
  bfr _b_854(.a(_w_1186),.q(_w_1187));
  bfr _b_1041(.a(_w_1373),.q(_w_1374));
  bfr _b_1476(.a(_w_1808),.q(_w_1809));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(_w_1848));
  bfr _b_1048(.a(_w_1380),.q(_w_1381));
  bfr _b_499(.a(_w_831),.q(_w_832));
  bfr _b_608(.a(_w_940),.q(_w_941));
  bfr _b_822(.a(_w_1154),.q(_w_1155));
  bfr _b_1050(.a(_w_1382),.q(_w_1383));
  spl2 N17_s_2(.a(N17_4),.q0(N17_5),.q1(N17_6));
  and_bi g139(.a(n128_1),.b(n137_1),.q(n139));
  bfr _b_954(.a(_w_1286),.q(_w_1287));
  bfr _b_936(.a(_w_1268),.q(_w_1269));
  bfr _b_1053(.a(_w_1385),.q(_w_1386));
  bfr _b_1296(.a(_w_1628),.q(_w_1629));
  bfr _b_1058(.a(_w_1390),.q(_w_1391));
  bfr _b_1185(.a(_w_1517),.q(_w_1518));
  bfr _b_1059(.a(_w_1391),.q(_w_1392));
  bfr _b_1223(.a(_w_1555),.q(_w_1556));
  bfr _b_1062(.a(_w_1394),.q(_w_1395));
  bfr _b_1064(.a(_w_1396),.q(_w_1397));
  bfr _b_1065(.a(_w_1397),.q(_w_1398));
  bfr _b_978(.a(_w_1310),.q(_w_1311));
  bfr _b_1107(.a(_w_1439),.q(N388));
  bfr _b_1665(.a(_w_1997),.q(_w_1998));
  bfr _b_529(.a(_w_861),.q(_w_862));
  bfr _b_1068(.a(_w_1400),.q(_w_1401));
  bfr _b_1070(.a(_w_1402),.q(_w_1403));
  bfr _b_1071(.a(_w_1403),.q(_w_1404));
  bfr _b_1072(.a(_w_1404),.q(_w_1405));
  bfr _b_1184(.a(_w_1516),.q(_w_1517));
  bfr _b_561(.a(_w_893),.q(N149_1));
  bfr _b_1074(.a(_w_1406),.q(N421));
  bfr _b_1803(.a(_w_2135),.q(_w_2136));
  bfr _b_1075(.a(_w_1407),.q(_w_1408));
  bfr _b_1076(.a(_w_1408),.q(_w_1409));
  bfr _b_1438(.a(_w_1770),.q(_w_1771));
  bfr _b_1078(.a(_w_1410),.q(_w_1411));
  bfr _b_881(.a(_w_1213),.q(_w_1214));
  bfr _b_1080(.a(_w_1412),.q(_w_1413));
  bfr _b_1081(.a(_w_1413),.q(_w_1414));
  bfr _b_621(.a(_w_953),.q(N237_5));
  bfr _b_1082(.a(_w_1414),.q(_w_1415));
  bfr _b_1084(.a(_w_1416),.q(_w_1417));
  bfr _b_1088(.a(_w_1420),.q(_w_1421));
  bfr _b_1718(.a(_w_2050),.q(_w_2051));
  spl3L g352_s_0(.a(n352),.q0(n352_0),.q1(n352_1),.q2(n352_2));
  bfr _b_805(.a(_w_1137),.q(_w_1138));
  bfr _b_1089(.a(_w_1421),.q(_w_1422));
  bfr _b_1090(.a(_w_1422),.q(_w_1423));
  spl2 N75_s_0(.a(N75),.q0(N75_0),.q1(N75_1));
  bfr _b_1093(.a(_w_1425),.q(_w_1426));
  bfr _b_1094(.a(_w_1426),.q(_w_1427));
  bfr _b_900(.a(_w_1232),.q(N159_2));
  bfr _b_819(.a(_w_1151),.q(_w_1152));
  bfr _b_1095(.a(_w_1427),.q(_w_1428));
  bfr _b_1099(.a(_w_1431),.q(_w_1432));
  bfr _b_1101(.a(_w_1433),.q(_w_1434));
  bfr _b_1104(.a(_w_1436),.q(_w_1437));
  bfr _b_1612(.a(_w_1944),.q(_w_1945));
  bfr _b_1106(.a(_w_1438),.q(_w_1439));
  bfr _b_1558(.a(_w_1890),.q(_w_1891));
  bfr _b_1108(.a(_w_1440),.q(_w_1441));
endmodule
