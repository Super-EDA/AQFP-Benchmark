module c1908 (G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G4,G5,G6,G7,G8,G9,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908);
  input G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G4,G5,G6,G7,G8,G9;
  output G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908;
  wire _w_1854,_w_1851,_w_1850,_w_1849,_w_1848,_w_1846,_w_1841,_w_1840,_w_1839,_w_1838,_w_1836,_w_1829,_w_1828,_w_1827,_w_1826,_w_1825,_w_1824,_w_1823,_w_1820,_w_1819,_w_1818,_w_1816,_w_1811,_w_1810,_w_1808,_w_1805,_w_1835,_w_1803,_w_1802,_w_1799,_w_1797,_w_1794,_w_1793,_w_1792,_w_1791,_w_1790,_w_1789,_w_1787,_w_1853,_w_1784,_w_1783,_w_1782,_w_1781,_w_1780,_w_1779,_w_1778,_w_1777,_w_1776,_w_1775,_w_1774,_w_1772,_w_1771,_w_1770,_w_1768,_w_1766,_w_1763,_w_1760,_w_1759,_w_1757,_w_1755,_w_1752,_w_1747,_w_1744,_w_1743,_w_1738,_w_1731,_w_1726,_w_1724,_w_1720,_w_1719,_w_1718,_w_1716,_w_1714,_w_1812,_w_1712,_w_1711,_w_1710,_w_1707,_w_1706,_w_1704,_w_1703,_w_1700,_w_1698,_w_1695,_w_1694,_w_1687,_w_1685,_w_1680,_w_1676,_w_1674,_w_1673,_w_1672,_w_1666,_w_1665,_w_1660,_w_1814,_w_1658,_w_1657,_w_1655,_w_1654,_w_1653,_w_1652,_w_1649,_w_1644,_w_1642,_w_1641,_w_1639,_w_1832,_w_1638,_w_1637,_w_1634,_w_1633,_w_1630,_w_1626,_w_1625,_w_1623,_w_1622,_w_1614,_w_1612,_w_1611,_w_1609,_w_1606,_w_1605,_w_1603,_w_1601,_w_1597,_w_1595,_w_1592,_w_1590,_w_1589,_w_1588,_w_1833,_w_1584,_w_1582,_w_1581,_w_1580,_w_1579,_w_1578,_w_1837,_w_1576,_w_1575,_w_1574,_w_1573,_w_1572,_w_1571,_w_1570,_w_1569,_w_1567,_w_1565,_w_1645,_w_1563,_w_1561,_w_1559,_w_1558,_w_1557,_w_1552,_w_1551,_w_1550,_w_1549,_w_1548,_w_1545,_w_1543,_w_1542,_w_1541,_w_1555,_w_1537,_w_1535,_w_1534,_w_1544,_w_1533,_w_1532,_w_1530,_w_1693,_w_1560,_w_1527,_w_1524,_w_1831,_w_1522,_w_1520,_w_1519,_w_1518,_w_1513,_w_1511,_w_1510,_w_1507,_w_1505,_w_1502,_w_1501,_w_1499,_w_1497,_w_1495,_w_1494,_w_1761,_w_1493,_w_1492,_w_1491,_w_1490,_w_1489,_w_1488,_w_1806,_w_1486,_w_1484,_w_1482,_w_1481,_w_1809,_w_1479,_w_1478,_w_1476,_w_1474,_w_1472,_w_1471,_w_1470,_w_1469,_w_1467,_w_1628,_w_1465,_w_1463,_w_1460,_w_1457,_w_1456,_w_1452,_w_1451,_w_1447,_w_1444,_w_1855,_w_1443,_w_1442,_w_1441,_w_1440,_w_1439,_w_1648,_w_1438,_w_1434,_w_1433,_w_1427,_w_1425,_w_1424,_w_1423,_w_1667,_w_1422,_w_1496,_w_1420,_w_1656,_w_1419,_w_1475,_w_1417,_w_1415,_w_1414,_w_1413,_w_1410,_w_1406,_w_1405,_w_1402,_w_1400,_w_1399,_w_1616,_w_1392,_w_1515,_w_1391,_w_1390,_w_1388,_w_1387,_w_1383,_w_1547,_w_1381,_w_1379,_w_1678,_w_1376,_w_1375,_w_1371,_w_1705,_w_1454,_w_1370,_w_1369,_w_1713,_w_1368,_w_1367,_w_1365,_w_1364,_w_1362,_w_1360,_w_1358,_w_1357,_w_1356,_w_1354,_w_1677,_w_1353,_w_1350,_w_1348,_w_1346,_w_1343,_w_1342,_w_1430,_w_1339,_w_1807,_w_1337,_w_1335,_w_1334,_w_1598,_w_1344,_w_1333,_w_1332,_w_1331,_w_1330,_w_1699,_w_1329,_w_1327,_w_1323,_w_1322,_w_1321,_w_1320,_w_1319,_w_1318,_w_1315,_w_1312,_w_1310,_w_1307,_w_1306,_w_1303,_w_1301,_w_1300,_w_1297,_w_1296,_w_1295,_w_1689,_w_1294,_w_1293,_w_1291,_w_1290,_w_1288,_w_1546,_w_1287,_w_1521,_w_1286,_w_1285,_w_1349,_w_1284,_w_1283,_w_1282,_w_1280,_w_1279,_w_1277,_w_1276,_w_1275,_w_1709,_w_1271,_w_1485,_w_1270,_w_1264,_w_1263,_w_1748,_w_1262,_w_1261,_w_1259,_w_1688,_w_1257,_w_1255,_w_1254,_w_1253,_w_1459,_w_1251,_w_1250,_w_1340,_w_1249,_w_1248,_w_1242,_w_1237,_w_1596,_w_1233,_w_1232,_w_1230,_w_1228,_w_1224,_w_1222,_w_1428,_w_1221,_w_1409,_w_1243,_w_1220,_w_1480,_w_1217,_w_1735,_w_1215,_w_1214,_w_1213,_w_1211,_w_1210,_w_1206,_w_1204,_w_1203,_w_1201,_w_1200,_w_1199,_w_1197,_w_1196,_w_1585,_w_1194,_w_1191,_w_1190,_w_1817,_w_1187,_w_1432,_w_1184,_w_1219,_w_1183,_w_1182,_w_1180,_w_1179,_w_1176,_w_1174,_w_1173,_w_1171,_w_1664,_w_1166,_w_1164,_w_1396,_w_1163,_w_1161,_w_1159,_w_1483,_w_1158,_w_1157,_w_1156,_w_1246,_w_1155,_w_1152,_w_1151,_w_1150,_w_1617,_w_1146,_w_1145,_w_1140,_w_1139,_w_1138,_w_1137,_w_1134,_w_1131,_w_1130,_w_1129,_w_1127,_w_1126,_w_1122,_w_1121,_w_1120,_w_1118,_w_1117,_w_1216,_w_1115,_w_1114,_w_1435,_w_1113,_w_1112,_w_1111,_w_1110,G22_0,_w_795,_w_934,_w_1785,n135,G11_7,_w_906,n182_1,n57_1,_w_956,_w_1056,n42,n205_0,n172_1,n199_0,_w_1341,n273,n105_2,G19_0,_w_1377,_w_853,G21_0,n110_1,n113_1,_w_1822,n235,n235_8,G24_3,n163,_w_825,_w_862,G5_1,G33_9,G33_8,G33_6,_w_1737,G15_5,_w_860,G33_1,G16_6,n78_0,G16_4,G16_3,n203_7,G16_1,n41_4,_w_1696,n206_6,_w_1773,_w_1729,n109_0,n199_1,n142_1,n203_0,n222_10,n41_3,_w_1722,n222_8,n222_4,n222_3,_w_1345,_w_802,n222_2,_w_1503,n203_9,_w_1756,n222_1,_w_928,n222_0,n248,G10_6,G2_5,G2_4,_w_1593,G2_2,n309,G1_2,_w_1728,n137,_w_922,G28_0,n316,G19_1,n60_1,n162,n50_3,_w_1272,n50_2,_w_1205,_w_1198,n47_1,n128,n56_2,n72_0,_w_1715,_w_1070,n235_3,_w_1607,n56_1,_w_1477,_w_953,_w_1325,_w_847,n35_3,_w_1256,n275_0,n34_0,_w_1830,G15_7,n145_1,_w_1053,G15_6,_w_1177,G5_3,G15_4,G15_2,G15_1,_w_880,_w_1075,n92_1,_w_1734,_w_1352,_w_1202,G33_14,n89,_w_1235,n92_0,n161_1,n141,n87_7,n50_1,n103,n234,_w_1758,G33_2,n87_5,_w_1226,n258,n87_0,_w_867,_w_1643,G29_0,_w_938,n88_1,G16_7,_w_913,G15_3,_w_1175,G8_2,_w_871,n146,_w_1845,n95_1,_w_887,G30_1,G4_3,_w_1241,n254_6,_w_1701,n105_3,G26_2,n182,_w_1355,n254_4,G25_1,G31_20,n185_1,_w_1458,n254_3,n61,_w_884,G10_4,G2_3,n312_1,n317,n320,_w_1506,n318,G1_7,_w_1144,_w_1154,n310,n239,_w_1188,_w_1092,n46,n308,n108_1,n57_0,_w_833,n306,_w_891,n304,n199,n300,n113_0,_w_1487,_w_1236,n297,_w_1553,_w_1010,G15_0,G9_7,_w_1635,n296,G28_1,n265,n34,_w_1108,_w_1229,G1_6,n284,n72_1,n283,n268,n282,G31_14,n281,_w_1723,n302,n233,_w_976,G24_2,n53_0,n152_0,_w_1148,n276,G16_0,n142_0,n116_0,n272,_w_1668,n206_4,_w_963,_w_994,_w_1398,G27_2,n262,_w_1834,n50_0,n259,_w_978,_w_1227,_w_998,G10_7,n106,_w_1192,n113,G1_0,n252,n250,_w_1621,n254_5,_w_1708,_w_1269,n315,n114,_w_1308,G2_0,_w_1671,n300_0,_w_1554,n246,_w_1462,n245,G16_5,G7_5,_w_1446,n195_1,n206_12,n243,_w_1133,n60_0,n261,_w_1351,G14_6,_w_807,_w_1681,G1_4,G8_8,G24_1,_w_1473,n304_1,n74_1,_w_1064,n153,n186,_w_1366,n198_0,_w_902,n291,n86,G8_10,G9_3,n87,_w_1384,n85,n161,n254_9,n81,_w_1577,n80,_w_1762,_w_820,_w_1162,n281_1,n293,_w_1741,n184,n156,_w_1167,n188_1,_w_1195,n79,G31_19,n73_1,n96,_w_1260,n305,_w_1382,n54,_w_897,n195,n198,G33_7,n174,_w_1101,_w_952,_w_1448,n41,n65,n64,_w_1753,_w_1119,G10_1,n87_1,G16_2,_w_1087,n145,_w_921,n313,_w_1105,n173,_w_1632,_w_1181,_w_828,_w_1842,G8_0,n182_0,_w_1586,n56,G5_6,_w_1717,n87_4,_w_1085,n125,_w_1032,_w_1153,G31_6,n227,n53,n148_1,G11_2,_w_1436,n52,n72,n55,G5_0,n47_0,n50,n221_2,_w_1691,n40,n53_1,n49,n221_0,_w_1461,_w_842,_w_1000,_w_1764,n47,n41_2,n74,G11_5,n60,_w_1239,n71,n68,_w_925,_w_1536,G8_3,n289,_w_1646,_w_1149,_w_1421,_w_1038,G13_2,_w_1683,_w_1526,G9_6,G9_0,n206_1,n200,_w_1404,_w_972,n109_1,_w_1629,_w_949,n109,n59,n78,n67,_w_810,_w_1373,_w_918,_w_1613,n58,_w_1292,n128_1,G5_5,_w_967,_w_1843,G33_10,_w_1608,_w_1063,G10_3,G4_7,n101,n90,_w_1662,_w_1273,n95_0,_w_1750,_w_1800,_w_837,n89_1,n75,_w_1566,n131,n38_1,n292,G4_10,n172,_w_1684,_w_816,n105_4,n159,n179_1,n205,n222_7,n217,n111,n235_2,n316_1,_w_1095,n87_6,n82,_w_1096,_w_1821,_w_1453,n77,G1_5,n176,_w_1767,_w_1509,_w_1169,G33_0,G11_1,G10_5,n57,n132,n196,G11_6,_w_1568,_w_1650,G33_3,_w_1796,_w_1274,_w_995,n277,n76,_w_1314,n48,G2_1,n203_6,G7_3,G4_5,n169,n128_0,_w_1528,G13_7,n91,_w_1587,n35_1,_w_1801,G26_0,_w_1393,_w_869,_w_1209,_w_872,G25_2,_w_1651,n177_1,G10_2,n301,n66_0,_w_1225,_w_969,G5_2,_w_1844,n281_0,G12_0,n311,_w_950,_w_1788,_w_1143,n87_2,_w_1769,n197,n94,n117,n124,_w_1240,_w_948,n271,n172_0,n151,n303,n89_0,_w_966,_w_1599,G31_18,n275_1,n178,n154,_w_1401,n254_0,_w_1464,n145_0,n105,G8_9,_w_1372,_w_1223,n44,n129,n83,n203_4,_w_1278,_w_1172,_w_1071,_w_1426,n177,_w_1304,n211,G22_1,n192,n88_0,_w_818,n312_0,_w_1313,n171,_w_1449,n287,_w_1065,n112,n73_0,n69,_w_1407,_w_939,_w_1186,n254_2,_w_1073,_w_1231,n39,n311_1,G33_13,_w_1640,_w_1512,n84_1,n144,_w_1316,n164,_w_936,n104,n93,_w_1266,n56_0,n255,n267_0,n223,n222_9,n110,n63_0,_w_1001,_w_1378,G33_11,n187,n311_0,G8_4,n242,_w_1094,n206,n116,n206_2,_w_1302,G30_0,n206_0,_w_1636,_w_1252,G10_0,n51,G31_12,n222_11,G26_1,_w_806,n120,n122,_w_1247,n125_1,_w_874,_w_1006,n105_1,n123,_w_1374,n98_1,_w_937,n127,_w_1234,G33_4,n256,_w_1123,_w_912,_w_1631,_w_1142,_w_1078,_w_1077,_w_1099,n130,n248_0,n175,_w_1619,_w_1281,G23_3,_w_1125,_w_979,n81_1,_w_926,n224,_w_852,_w_942,n133,n118,n235_1,n136,n216,_w_1514,n267,n254_8,G31_8,_w_1395,_w_857,G3_1,n168,_w_831,n314,n97,n66,_w_1265,n204,n138,n100,_w_1027,_w_1135,n41_1,n139,n288,n158,_w_993,G2_6,n84,n207,_w_1765,G33_5,G11_3,n151_0,n249,G12_1,n321,n147,n222_6,n108_2,n148,_w_1659,n254_7,n142,G1_3,_w_798,n115,_w_885,G29_1,_w_973,_w_1591,_w_1508,G1_1,n202,_w_896,n226,n234_1,_w_1397,G11_4,n152,G27_1,n180,n155,n157,n136_1,_w_1385,n193,_w_1061,n143,_w_1326,_w_1189,_w_1042,n185,_w_1268,G3_3,n214,n160,n203_5,_w_927,n222_5,_w_803,n194,n81_0,G4_9,n165,n166,_w_1178,n181,n183,G3_6,n206_8,_w_1504,n235_5,n300_1,_w_1538,n77_2,_w_1847,_w_1258,n43,n205_1,G18_1,_w_1682,_w_1084,n189,_w_907,n70,_w_935,_w_899,n125_0,n190,n229,n191,n201,_w_982,n236,_w_1539,n162_1,_w_845,n99,_w_1389,n195_0,_w_1005,n203,_w_1289,n41_0,n66_1,_w_1615,_w_1107,n208,n88,G8_7,G3_7,n213,G3_5,n220,_w_1128,_w_841,n295,_w_886,_w_1523,n230,n77_0,n232,_w_1359,n149,G8_6,n237,n73_2,G3_0,G3_2,n102,G3_4,_w_1305,n119_0,_w_916,n35,n119_1,_w_1702,n77_1,_w_1018,n197_1,G32_0,_w_1104,G11_0,G32_1,n178_0,_w_1361,_w_989,n178_1,_w_910,_w_1082,_w_1742,_w_1098,_w_1008,n219,n204_0,G17_0,_w_1583,G6_0,_w_1795,n34_1,n316_0,G17_1,G6_1,G6_2,_w_1562,G4_6,G6_3,_w_1749,G6_4,n170,G6_5,_w_1324,_w_915,G6_6,_w_1062,n108,G6_7,_w_1338,n140,G7_0,_w_1733,G7_1,G7_4,_w_856,_w_1445,G8_5,G7_6,G7_7,n270,G18_0,G9_1,_w_1620,_w_1045,G9_2,_w_1721,G9_4,_w_1564,_w_1380,G13_6,_w_1141,G9_5,n37,n44_0,_w_1147,n44_1,_w_1813,_w_1540,_w_1309,n177_0,n200_1,_w_1498,_w_1103,_w_1431,G31_9,_w_848,n177_2,n177_3,n299_1,n198_1,G31_0,_w_888,G31_1,G31_2,G31_3,_w_1600,_w_1466,_w_808,G31_5,_w_965,G23_2,G31_7,_w_1311,G14_2,_w_1663,_w_1109,_w_908,G31_11,G33_12,G31_13,_w_1745,_w_813,G31_15,_w_954,G31_16,G31_17,n304_0,G20_0,G5_4,G5_7,n122_0,n35_0,n35_2,n74_0,n74_2,_w_1049,n98_0,n171_0,n221,_w_829,n188,n178_2,n108_0,n108_3,n110_0,_w_1679,_w_1067,n98,n206_3,_w_929,_w_1675,n206_5,G12_2,_w_1525,n210,n206_7,n206_9,n69_1,G7_2,_w_900,n206_11,n206_13,_w_1106,_w_1208,n116_1,n122_1,G4_0,G4_1,_w_1739,_w_1002,G4_2,G4_4,G4_8,n126_0,n126_1,_w_1604,n127_0,_w_1556,n128_2,_w_1394,n203_1,n133_0,n139_1,n201_1,n133_1,G14_3,G14_4,_w_1647,_w_801,_w_809,_w_981,G14_5,_w_1238,G21_1,G13_0,_w_1068,G13_1,G13_4,G13_5,n136_0,n267_1,n38_0,_w_991,G2_7,n267_2,_w_821,_w_1468,_w_1267,n267_3,n267_4,n36,G14_0,n267_5,n78_1,n267_6,n267_7,_w_1363,n168_0,n168_1,_w_827,n204_1,_w_964,n139_0,n158_1,n161_0,_w_1013,n84_0,_w_1136,n254_1,n63_1,_w_1450,n253,n63_2,n235_0,n63_3,_w_988,_w_1754,_w_1732,_w_1437,_w_1412,n148_0,_w_1015,n151_1,n152_1,G12_4,G12_5,_w_1011,G12_6,n158_0,G12_7,_w_1730,_w_1193,n185_0,n179,_w_1036,_w_1244,n162_0,_w_1624,n165_0,_w_1670,n127_1,n165_1,n92,n179_0,n188_0,n200_0,n191_0,_w_1037,n191_1,_w_1048,n192_0,_w_1661,_w_1429,_w_1298,n206_10,n192_1,n192_2,n45,n248_1,_w_958,n134,n105_0,n201_0,_w_1594,_w_1245,n87_3,n99_0,n203_2,n203_3,_w_844,_w_1627,_w_1610,n203_8,n312,n66_2,n219_0,n219_1,n221_1,_w_1531,_w_960,n234_0,n254,G20_1,n235_4,n235_6,n235_7,_w_1336,n171_1,_w_1020,n235_9,_w_1815,_w_1403,_w_1207,_w_974,_w_796,_w_797,_w_799,_w_804,n62,_w_811,_w_1132,_w_812,_w_962,_w_814,_w_815,_w_817,_w_1686,_w_822,n121,_w_1097,n119,_w_932,_w_1328,n240,_w_834,_w_1168,_w_835,_w_850,_w_1725,_w_836,_w_838,_w_1076,_w_839,_w_840,_w_1602,_w_843,_w_1418,n197_0,_w_846,n299_0,_w_849,_w_944,n278,_w_851,_w_1529,_w_854,_w_855,_w_858,_w_1618,_w_859,_w_861,_w_863,_w_864,G27_0,_w_1019,G31_4,_w_865,_w_868,G23_1,_w_870,_w_873,_w_1697,_w_875,_w_876,_w_1852,n178_3,_w_931,_w_1170,_w_1044,_w_866,_w_877,_w_1669,_w_878,_w_879,_w_881,_w_882,_w_883,_w_1299,_w_889,_w_890,_w_832,n299,_w_892,_w_893,_w_1727,_w_894,n99_1,_w_895,_w_898,n150,_w_901,_w_990,_w_903,n73,_w_904,_w_1804,_w_905,_w_909,_w_823,_w_911,n38,_w_914,_w_819,_w_917,_w_919,_w_1386,_w_826,_w_920,_w_1009,_w_923,_w_1124,_w_924,_w_930,_w_824,_w_933,n126,_w_940,_w_941,_w_943,_w_951,_w_945,_w_1455,_w_946,_w_947,_w_800,G14_7,_w_955,_w_957,_w_1212,_w_959,n107,_w_961,_w_1317,_w_968,_w_1411,G8_1,_w_970,_w_1690,_w_971,_w_1093,_w_975,_w_1517,_w_1408,n63,_w_977,_w_980,_w_983,_w_1786,_w_984,_w_985,_w_1160,_w_1024,n279,_w_986,_w_987,_w_992,_w_996,_w_997,_w_999,_w_1003,_w_1090,_w_1004,_w_1692,_w_1500,_w_1007,_w_1012,G14_1,_w_1025,_w_805,_w_1054,n66_3,G31_10,_w_1014,_w_1751,_w_1165,_w_1016,_w_1798,_w_1516,_w_1017,_w_1021,_w_1022,_w_1416,n285,_w_1023,_w_1026,n195_2,_w_1028,_w_1029,_w_1030,_w_1736,_w_1347,_w_1031,n264,_w_1040,n269,_w_1033,_w_1746,_w_794,n222,_w_1034,_w_1035,G13_3,_w_1039,_w_1041,_w_1043,G23_0,_w_1046,G24_0,_w_1047,_w_1116,G28_2,_w_1050,_w_1051,_w_1052,_w_1055,_w_1185,_w_1057,G25_0,n275,_w_1058,_w_1059,n167,G12_3,_w_1060,_w_1066,_w_1069,_w_1072,n69_0,_w_1074,_w_1740,_w_1079,_w_1080,_w_1081,_w_1218,_w_830,_w_1083,n95,_w_1086,_w_1088,_w_1089,_w_1091,_w_1100,_w_1102;

  bfr _b_1539(.a(_w_1853),.q(_w_1854));
  bfr _b_1537(.a(G7),.q(_w_1851));
  bfr _b_1536(.a(G6),.q(_w_1850));
  bfr _b_1535(.a(_w_1849),.q(_w_1847));
  bfr _b_1533(.a(G5),.q(_w_1848));
  bfr _b_1541(.a(G9),.q(_w_1855));
  bfr _b_1528(.a(_w_1842),.q(_w_1843));
  bfr _b_1526(.a(_w_1840),.q(_w_1841));
  bfr _b_1523(.a(_w_1837),.q(_w_1838));
  bfr _b_1522(.a(_w_1836),.q(_w_1837));
  bfr _b_1521(.a(_w_1835),.q(_w_1836));
  bfr _b_1520(.a(_w_1834),.q(_w_1835));
  bfr _b_1519(.a(_w_1833),.q(_w_1834));
  bfr _b_1516(.a(G30),.q(_w_1830));
  bfr _b_1515(.a(_w_1829),.q(_w_1814));
  bfr _b_1513(.a(_w_1827),.q(_w_1828));
  bfr _b_1512(.a(_w_1826),.q(_w_1827));
  bfr _b_1507(.a(_w_1821),.q(_w_1822));
  bfr _b_1506(.a(_w_1820),.q(_w_1821));
  bfr _b_1504(.a(_w_1818),.q(_w_1819));
  bfr _b_1503(.a(_w_1817),.q(_w_1818));
  bfr _b_1501(.a(_w_1815),.q(_w_1816));
  bfr _b_1500(.a(G29),.q(_w_1815));
  bfr _b_1499(.a(_w_1813),.q(_w_1800));
  bfr _b_1497(.a(_w_1811),.q(_w_1812));
  bfr _b_1496(.a(_w_1810),.q(_w_1811));
  bfr _b_1495(.a(_w_1809),.q(_w_1810));
  bfr _b_1493(.a(_w_1807),.q(_w_1808));
  bfr _b_1491(.a(_w_1805),.q(_w_1806));
  bfr _b_1490(.a(_w_1804),.q(_w_1805));
  bfr _b_1489(.a(_w_1803),.q(_w_1804));
  bfr _b_1485(.a(_w_1799),.q(_w_1785));
  bfr _b_1480(.a(_w_1794),.q(_w_1795));
  bfr _b_1479(.a(_w_1793),.q(_w_1794));
  bfr _b_1475(.a(_w_1789),.q(_w_1790));
  bfr _b_1474(.a(_w_1788),.q(_w_1789));
  bfr _b_1473(.a(_w_1787),.q(_w_1788));
  bfr _b_1472(.a(_w_1786),.q(_w_1787));
  bfr _b_1470(.a(_w_1784),.q(_w_1770));
  bfr _b_1468(.a(_w_1782),.q(_w_1783));
  bfr _b_1466(.a(_w_1780),.q(_w_1781));
  bfr _b_1465(.a(_w_1779),.q(_w_1780));
  bfr _b_1463(.a(_w_1777),.q(_w_1778));
  bfr _b_1462(.a(_w_1776),.q(_w_1777));
  bfr _b_1459(.a(_w_1773),.q(_w_1774));
  bfr _b_1458(.a(_w_1772),.q(_w_1773));
  bfr _b_1456(.a(G26),.q(_w_1771));
  bfr _b_1455(.a(_w_1769),.q(_w_1754));
  bfr _b_1454(.a(_w_1768),.q(_w_1769));
  bfr _b_1453(.a(_w_1767),.q(_w_1768));
  bfr _b_1450(.a(_w_1764),.q(_w_1765));
  bfr _b_1449(.a(_w_1763),.q(_w_1764));
  bfr _b_1444(.a(_w_1758),.q(_w_1759));
  bfr _b_1461(.a(_w_1775),.q(_w_1776));
  bfr _b_1441(.a(_w_1755),.q(_w_1756));
  bfr _b_1440(.a(G25),.q(_w_1755));
  bfr _b_1433(.a(_w_1747),.q(_w_1746));
  bfr _b_1432(.a(G18),.q(_w_1747));
  bfr _b_1429(.a(_w_1743),.q(_w_1741));
  bfr _b_1427(.a(G16),.q(_w_1742));
  bfr _b_1426(.a(_w_1740),.q(_w_1739));
  bfr _b_1424(.a(_w_1738),.q(_w_1736));
  bfr _b_1423(.a(_w_1737),.q(_w_1738));
  bfr _b_1422(.a(G1),.q(_w_1737));
  bfr _b_1420(.a(_w_1734),.q(_w_1735));
  bfr _b_1419(.a(_w_1733),.q(_w_1734));
  bfr _b_1418(.a(_w_1732),.q(n69));
  bfr _b_1417(.a(_w_1731),.q(_w_1732));
  bfr _b_1416(.a(_w_1730),.q(_w_1731));
  bfr _b_1412(.a(_w_1726),.q(G31_4));
  bfr _b_1410(.a(_w_1724),.q(_w_1725));
  bfr _b_1409(.a(_w_1723),.q(_w_1724));
  bfr _b_1408(.a(_w_1722),.q(_w_1723));
  bfr _b_1407(.a(_w_1721),.q(_w_1722));
  bfr _b_1406(.a(_w_1720),.q(_w_1721));
  bfr _b_1405(.a(_w_1719),.q(_w_1720));
  bfr _b_1404(.a(_w_1718),.q(_w_1719));
  bfr _b_1403(.a(_w_1717),.q(_w_1718));
  bfr _b_1402(.a(_w_1716),.q(G31_2));
  bfr _b_1399(.a(_w_1713),.q(_w_1714));
  bfr _b_1398(.a(_w_1712),.q(_w_1713));
  bfr _b_1396(.a(_w_1710),.q(_w_1711));
  bfr _b_1391(.a(_w_1705),.q(_w_1706));
  bfr _b_1388(.a(_w_1702),.q(G1897));
  bfr _b_1387(.a(_w_1701),.q(_w_1702));
  bfr _b_1384(.a(_w_1698),.q(G1893));
  bfr _b_1381(.a(_w_1695),.q(_w_1696));
  bfr _b_1380(.a(_w_1694),.q(n232));
  bfr _b_1379(.a(_w_1693),.q(G1890));
  bfr _b_1378(.a(_w_1692),.q(_w_1693));
  bfr _b_1377(.a(_w_1691),.q(_w_1692));
  bfr _b_1413(.a(_w_1727),.q(_w_1728));
  bfr _b_1375(.a(_w_1689),.q(_w_1690));
  bfr _b_1374(.a(_w_1688),.q(_w_1689));
  bfr _b_1373(.a(_w_1687),.q(_w_1688));
  bfr _b_1371(.a(_w_1685),.q(_w_1686));
  bfr _b_1369(.a(_w_1683),.q(_w_1684));
  bfr _b_1366(.a(_w_1680),.q(n221));
  bfr _b_1364(.a(_w_1678),.q(_w_1679));
  bfr _b_1360(.a(_w_1674),.q(_w_1675));
  bfr _b_1359(.a(_w_1673),.q(_w_1674));
  bfr _b_1356(.a(_w_1670),.q(_w_1671));
  bfr _b_1354(.a(_w_1668),.q(_w_1669));
  bfr _b_1352(.a(_w_1666),.q(_w_1667));
  bfr _b_1351(.a(_w_1665),.q(_w_1666));
  bfr _b_1350(.a(_w_1664),.q(_w_1665));
  bfr _b_1349(.a(_w_1663),.q(_w_1664));
  bfr _b_1348(.a(_w_1662),.q(_w_1663));
  bfr _b_1347(.a(_w_1661),.q(_w_1662));
  bfr _b_1460(.a(_w_1774),.q(_w_1775));
  bfr _b_1345(.a(_w_1659),.q(_w_1660));
  bfr _b_1342(.a(_w_1656),.q(_w_1657));
  bfr _b_1341(.a(_w_1655),.q(_w_1656));
  bfr _b_1338(.a(_w_1652),.q(_w_1653));
  bfr _b_1337(.a(_w_1651),.q(G1888));
  bfr _b_1336(.a(_w_1650),.q(_w_1651));
  bfr _b_1335(.a(_w_1649),.q(_w_1650));
  bfr _b_1334(.a(_w_1648),.q(G1886));
  bfr _b_1330(.a(_w_1644),.q(_w_1645));
  bfr _b_1329(.a(_w_1643),.q(_w_1644));
  bfr _b_1325(.a(_w_1639),.q(n273));
  bfr _b_1332(.a(_w_1646),.q(_w_1647));
  bfr _b_1322(.a(_w_1636),.q(_w_1637));
  bfr _b_1321(.a(_w_1635),.q(_w_1636));
  bfr _b_1320(.a(_w_1634),.q(_w_1635));
  bfr _b_1525(.a(_w_1839),.q(_w_1840));
  bfr _b_1319(.a(_w_1633),.q(n191));
  bfr _b_1317(.a(_w_1631),.q(G1892));
  bfr _b_1314(.a(_w_1628),.q(_w_1629));
  bfr _b_1312(.a(_w_1626),.q(_w_1627));
  bfr _b_1397(.a(_w_1711),.q(_w_1712));
  bfr _b_1311(.a(_w_1625),.q(G2_2));
  bfr _b_1307(.a(_w_1621),.q(_w_1622));
  bfr _b_1306(.a(_w_1620),.q(_w_1621));
  bfr _b_1305(.a(_w_1619),.q(G1896));
  bfr _b_1304(.a(_w_1618),.q(_w_1619));
  bfr _b_1303(.a(_w_1617),.q(_w_1618));
  bfr _b_1302(.a(_w_1616),.q(_w_1617));
  bfr _b_1301(.a(_w_1615),.q(G9_2));
  bfr _b_1300(.a(_w_1614),.q(G26_2));
  bfr _b_1298(.a(_w_1612),.q(_w_1613));
  bfr _b_1297(.a(_w_1611),.q(_w_1612));
  bfr _b_1295(.a(_w_1609),.q(_w_1610));
  bfr _b_1294(.a(_w_1608),.q(_w_1609));
  bfr _b_1290(.a(_w_1604),.q(_w_1605));
  bfr _b_1289(.a(_w_1603),.q(_w_1604));
  bfr _b_1514(.a(_w_1828),.q(_w_1829));
  bfr _b_1287(.a(_w_1601),.q(_w_1602));
  bfr _b_1283(.a(_w_1597),.q(G1903));
  bfr _b_1282(.a(_w_1596),.q(n72_1));
  bfr _b_1279(.a(_w_1593),.q(_w_1594));
  bfr _b_1276(.a(_w_1590),.q(_w_1591));
  bfr _b_1274(.a(_w_1588),.q(_w_1589));
  bfr _b_1278(.a(_w_1592),.q(_w_1593));
  bfr _b_1272(.a(_w_1586),.q(_w_1587));
  bfr _b_1268(.a(_w_1582),.q(_w_1583));
  bfr _b_1277(.a(_w_1591),.q(_w_1592));
  bfr _b_1267(.a(_w_1581),.q(_w_1582));
  bfr _b_1264(.a(_w_1578),.q(_w_1579));
  bfr _b_1299(.a(_w_1613),.q(_w_1614));
  bfr _b_1262(.a(_w_1576),.q(_w_1577));
  bfr _b_1259(.a(_w_1573),.q(_w_1574));
  bfr _b_1253(.a(_w_1567),.q(G1895));
  bfr _b_1250(.a(_w_1564),.q(_w_1565));
  bfr _b_1249(.a(_w_1563),.q(_w_1564));
  bfr _b_1248(.a(_w_1562),.q(n308));
  bfr _b_1247(.a(_w_1561),.q(_w_1562));
  bfr _b_1372(.a(_w_1686),.q(G1894));
  bfr _b_1246(.a(_w_1560),.q(_w_1561));
  bfr _b_1243(.a(_w_1557),.q(_w_1558));
  bfr _b_1242(.a(_w_1556),.q(_w_1557));
  bfr _b_1241(.a(_w_1555),.q(n74));
  bfr _b_1240(.a(_w_1554),.q(_w_1555));
  bfr _b_1324(.a(_w_1638),.q(_w_1639));
  bfr _b_1235(.a(_w_1549),.q(_w_1550));
  bfr _b_1234(.a(_w_1548),.q(_w_1549));
  bfr _b_1233(.a(_w_1547),.q(_w_1548));
  bfr _b_1361(.a(_w_1675),.q(_w_1676));
  bfr _b_1232(.a(_w_1546),.q(_w_1547));
  bfr _b_1230(.a(_w_1544),.q(n192_2));
  bfr _b_1229(.a(_w_1543),.q(_w_1544));
  bfr _b_1228(.a(_w_1542),.q(_w_1543));
  bfr _b_1227(.a(_w_1541),.q(_w_1542));
  bfr _b_1370(.a(_w_1684),.q(_w_1685));
  bfr _b_1323(.a(_w_1637),.q(_w_1638));
  bfr _b_1226(.a(_w_1540),.q(_w_1541));
  bfr _b_1224(.a(_w_1538),.q(_w_1539));
  bfr _b_1221(.a(_w_1535),.q(_w_1536));
  bfr _b_1270(.a(_w_1584),.q(_w_1585));
  bfr _b_1263(.a(_w_1577),.q(_w_1578));
  bfr _b_1220(.a(_w_1534),.q(_w_1535));
  bfr _b_1219(.a(_w_1533),.q(_w_1534));
  bfr _b_1217(.a(_w_1531),.q(_w_1532));
  bfr _b_1443(.a(_w_1757),.q(_w_1758));
  bfr _b_1216(.a(_w_1530),.q(n73_2));
  bfr _b_1362(.a(_w_1676),.q(_w_1677));
  bfr _b_1215(.a(_w_1529),.q(_w_1530));
  bfr _b_1214(.a(_w_1528),.q(_w_1529));
  bfr _b_1213(.a(_w_1527),.q(_w_1528));
  bfr _b_1211(.a(_w_1525),.q(_w_1526));
  bfr _b_1207(.a(_w_1521),.q(_w_1522));
  bfr _b_1206(.a(_w_1520),.q(_w_1521));
  bfr _b_1205(.a(_w_1519),.q(_w_1520));
  bfr _b_1204(.a(_w_1518),.q(_w_1519));
  bfr _b_1201(.a(_w_1515),.q(_w_1516));
  bfr _b_1200(.a(_w_1514),.q(_w_1515));
  bfr _b_1199(.a(_w_1513),.q(_w_1514));
  bfr _b_1198(.a(_w_1512),.q(_w_1513));
  bfr _b_1196(.a(_w_1510),.q(_w_1511));
  bfr _b_1194(.a(_w_1508),.q(_w_1509));
  bfr _b_1193(.a(_w_1507),.q(_w_1508));
  bfr _b_1192(.a(_w_1506),.q(_w_1507));
  bfr _b_1191(.a(_w_1505),.q(_w_1506));
  bfr _b_1190(.a(_w_1504),.q(_w_1505));
  bfr _b_1189(.a(_w_1503),.q(_w_1504));
  bfr _b_1187(.a(_w_1501),.q(_w_1502));
  bfr _b_1186(.a(_w_1500),.q(_w_1501));
  bfr _b_1180(.a(_w_1494),.q(n162));
  bfr _b_1179(.a(_w_1493),.q(_w_1494));
  bfr _b_1178(.a(_w_1492),.q(n125_1));
  bfr _b_1177(.a(_w_1491),.q(_w_1492));
  bfr _b_1176(.a(_w_1490),.q(_w_1491));
  bfr _b_1174(.a(_w_1488),.q(_w_1489));
  bfr _b_1173(.a(_w_1487),.q(_w_1488));
  bfr _b_1171(.a(_w_1485),.q(_w_1486));
  bfr _b_1169(.a(_w_1483),.q(_w_1484));
  bfr _b_1168(.a(_w_1482),.q(_w_1483));
  bfr _b_1167(.a(_w_1481),.q(_w_1482));
  bfr _b_1166(.a(_w_1480),.q(_w_1481));
  bfr _b_1163(.a(_w_1477),.q(_w_1478));
  bfr _b_1162(.a(_w_1476),.q(_w_1477));
  bfr _b_1161(.a(_w_1475),.q(n178));
  bfr _b_1159(.a(_w_1473),.q(_w_1474));
  bfr _b_1158(.a(_w_1472),.q(_w_1473));
  bfr _b_1157(.a(_w_1471),.q(_w_1472));
  bfr _b_1156(.a(_w_1470),.q(_w_1471));
  bfr _b_1154(.a(_w_1468),.q(_w_1469));
  bfr _b_1153(.a(_w_1467),.q(_w_1468));
  bfr _b_1152(.a(_w_1466),.q(_w_1467));
  bfr _b_1148(.a(_w_1462),.q(G33_12));
  bfr _b_1147(.a(_w_1461),.q(_w_1462));
  bfr _b_1146(.a(_w_1460),.q(_w_1461));
  bfr _b_1144(.a(_w_1458),.q(_w_1459));
  bfr _b_1141(.a(_w_1455),.q(_w_1456));
  bfr _b_1140(.a(_w_1454),.q(_w_1455));
  bfr _b_1138(.a(_w_1452),.q(_w_1453));
  bfr _b_1137(.a(_w_1451),.q(_w_1452));
  bfr _b_1136(.a(_w_1450),.q(_w_1451));
  bfr _b_1134(.a(_w_1448),.q(_w_1449));
  bfr _b_1133(.a(_w_1447),.q(_w_1448));
  bfr _b_1132(.a(_w_1446),.q(_w_1447));
  bfr _b_1293(.a(_w_1607),.q(_w_1608));
  bfr _b_1131(.a(_w_1445),.q(_w_1446));
  bfr _b_1129(.a(_w_1443),.q(_w_1444));
  bfr _b_1128(.a(_w_1442),.q(_w_1443));
  bfr _b_1127(.a(_w_1441),.q(_w_1442));
  bfr _b_1126(.a(_w_1440),.q(_w_1441));
  bfr _b_1124(.a(_w_1438),.q(_w_1439));
  bfr _b_1160(.a(_w_1474),.q(_w_1475));
  bfr _b_1122(.a(_w_1436),.q(_w_1437));
  bfr _b_1120(.a(_w_1434),.q(_w_1435));
  bfr _b_1119(.a(_w_1433),.q(_w_1434));
  bfr _b_1118(.a(_w_1432),.q(_w_1433));
  bfr _b_1114(.a(_w_1428),.q(_w_1429));
  bfr _b_1113(.a(_w_1427),.q(_w_1428));
  bfr _b_1111(.a(_w_1425),.q(_w_1426));
  bfr _b_1110(.a(_w_1424),.q(_w_1425));
  bfr _b_1109(.a(_w_1423),.q(_w_1424));
  bfr _b_538(.a(_w_852),.q(_w_853));
  bfr _b_537(.a(_w_851),.q(_w_852));
  bfr _b_536(.a(_w_850),.q(_w_851));
  and_bb g97(.a(n87_4),.b(n95_1),.q(n97));
  bfr _b_656(.a(_w_970),.q(_w_971));
  bfr _b_528(.a(_w_842),.q(_w_843));
  and_bi g276(.a(n275_0),.b(G31_19),.q(n276));
  bfr _b_524(.a(_w_838),.q(_w_839));
  bfr _b_523(.a(_w_837),.q(_w_838));
  bfr _b_522(.a(_w_836),.q(_w_837));
  bfr _b_517(.a(_w_831),.q(G13_2));
  bfr _b_1394(.a(_w_1708),.q(_w_1709));
  spl3L G9_s_1(.a(G9_2),.q0(G9_3),.q1(G9_4),.q2(_w_918));
  bfr _b_516(.a(_w_830),.q(_w_831));
  spl2 g197_s_0(.a(n197),.q0(n197_0),.q1(n197_1));
  spl2 g125_s_0(.a(n125),.q0(n125_0),.q1(_w_1476));
  bfr _b_511(.a(_w_825),.q(_w_826));
  bfr _b_509(.a(_w_823),.q(_w_824));
  bfr _b_785(.a(_w_1099),.q(_w_1100));
  bfr _b_815(.a(_w_1129),.q(_w_1130));
  bfr _b_1055(.a(_w_1369),.q(_w_1370));
  bfr _b_504(.a(_w_818),.q(_w_819));
  spl2 G13_s_2(.a(G13_5),.q0(G13_6),.q1(G13_7));
  and_bb g253(.a(n252),.b(n77_2),.q(n253));
  bfr _b_510(.a(_w_824),.q(_w_825));
  bfr _b_497(.a(_w_811),.q(G12_0));
  bfr _b_494(.a(_w_808),.q(_w_809));
  bfr _b_490(.a(_w_804),.q(_w_805));
  bfr _b_862(.a(_w_1176),.q(_w_1177));
  bfr _b_514(.a(_w_828),.q(n151_1));
  bfr _b_488(.a(_w_802),.q(_w_803));
  spl3L G15_s_1(.a(G15_2),.q0(G15_3),.q1(G15_4),.q2(_w_1360));
  and_bi g52(.a(n44_1),.b(n50_1),.q(n52));
  bfr _b_485(.a(_w_799),.q(_w_800));
  bfr _b_513(.a(_w_827),.q(_w_828));
  and_bi g271(.a(n77_1),.b(n270),.q(n271));
  bfr _b_480(.a(_w_794),.q(_w_795));
  bfr _b_767(.a(_w_1081),.q(_w_1082));
  bfr _b_1389(.a(_w_1703),.q(_w_1704));
  bfr _b_1183(.a(_w_1497),.q(G1887));
  spl4L g235_s_2(.a(n235_1),.q0(n235_6),.q1(n235_7),.q2(n235_8),.q3(n235_9));
  bfr _b_518(.a(_w_832),.q(_w_833));
  and_bb g138(.a(n133_1),.b(n136_1),.q(n138));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(n235_1));
  spl4L g203_s_3(.a(n203_5),.q0(n203_6),.q1(n203_7),.q2(n203_8),.q3(n203_9));
  spl2 g201_s_0(.a(n201),.q0(n201_0),.q1(n201_1));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(_w_794));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  and_bi g188(.a(n186),.b(n187),.q(n188));
  and_bi g295(.a(n128_2),.b(G31_17),.q(n295));
  and_bb g288(.a(n267_4),.b(n287),.q(n288));
  spl2 G12_s_0(.a(_w_1739),.q0(_w_811),.q1(G12_1));
  bfr _b_845(.a(_w_1159),.q(_w_1160));
  spl2 g151_s_0(.a(n151),.q0(n151_0),.q1(_w_812));
  or_bb g88(.a(G24_0),.b(G33_0),.q(n88));
  bfr _b_483(.a(_w_797),.q(_w_798));
  spl4L g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1),.q2(n63_2),.q3(n63_3));
  spl3L G14_s_1(.a(G14_2),.q0(G14_3),.q1(G14_4),.q2(_w_832));
  bfr _b_995(.a(_w_1309),.q(_w_1310));
  and_bi g83(.a(n81_1),.b(G12_2),.q(n83));
  bfr _b_1467(.a(_w_1781),.q(_w_1782));
  bfr _b_643(.a(_w_957),.q(_w_958));
  or_bb g274(.a(n268),.b(n273),.q(_w_1652));
  spl2 g122_s_0(.a(n122),.q0(n122_0),.q1(n122_1));
  bfr _b_1275(.a(_w_1589),.q(_w_1590));
  spl2 g116_s_0(.a(n116),.q0(n116_0),.q1(n116_1));
  or_bi g209(.a(n208),.b(n207),.q(_w_1598));
  spl4L g206_s_3(.a(n206_5),.q0(n206_10),.q1(n206_11),.q2(n206_12),.q3(n206_13));
  bfr _b_776(.a(_w_1090),.q(_w_1091));
  bfr _b_1016(.a(_w_1330),.q(_w_1331));
  spl2 g110_s_0(.a(n110),.q0(n110_0),.q1(n110_1));
  bfr _b_648(.a(_w_962),.q(_w_963));
  bfr _b_1245(.a(_w_1559),.q(_w_1560));
  spl2 g35_s_0(.a(n35),.q0(n35_0),.q1(_w_903));
  bfr _b_993(.a(_w_1307),.q(_w_1308));
  spl2 G5_s_2(.a(G5_5),.q0(G5_6),.q1(G5_7));
  or_bi g244(.a(n243),.b(n242),.q(_w_1695));
  spl2 G5_s_0(.a(_w_1847),.q0(_w_904),.q1(G5_1));
  spl2 G20_s_0(.a(_w_1750),.q0(G20_0),.q1(_w_905));
  spl2 G32_s_0(.a(_w_1832),.q0(G32_0),.q1(_w_985));
  spl2 g34_s_0(.a(n34),.q0(n34_0),.q1(n34_1));
  bfr _b_1261(.a(_w_1575),.q(_w_1576));
  bfr _b_872(.a(_w_1186),.q(_w_1187));
  spl3L g74_s_0(.a(n74),.q0(n74_0),.q1(n74_1),.q2(_w_892));
  bfr _b_484(.a(_w_798),.q(_w_799));
  bfr _b_1079(.a(_w_1393),.q(_w_1394));
  spl4L G31_s_6(.a(G31_14),.q0(G31_15),.q1(G31_16),.q2(G31_17),.q3(_w_906));
  and_bb g194(.a(G25_1),.b(n192_1),.q(n194));
  spl2 G31_s_5(.a(G31_12),.q0(G31_13),.q1(_w_907));
  and_bi g76(.a(n74_1),.b(n73_1),.q(n76));
  bfr _b_1271(.a(_w_1585),.q(_w_1586));
  and_bi g107(.a(G16_4),.b(n105_1),.q(n107));
  bfr _b_666(.a(_w_980),.q(_w_981));
  bfr _b_832(.a(_w_1146),.q(_w_1147));
  spl2 g127_s_0(.a(n127),.q0(n127_0),.q1(n127_1));
  spl4L G31_s_2(.a(G31_4),.q0(G31_5),.q1(G31_6),.q2(G31_7),.q3(G31_8));
  spl2 g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1));
  spl4L g267_s_0(.a(n267),.q0(n267_0),.q1(n267_1),.q2(n267_2),.q3(n267_3));
  spl2 g177_s_0(.a(n177),.q0(n177_0),.q1(n177_1));
  bfr _b_811(.a(_w_1125),.q(_w_1126));
  bfr _b_826(.a(_w_1140),.q(_w_1141));
  bfr _b_486(.a(_w_800),.q(_w_801));
  spl2 g44_s_0(.a(n44),.q0(n44_0),.q1(n44_1));
  bfr _b_1328(.a(_w_1642),.q(n205));
  spl3L G7_s_1(.a(G7_2),.q0(G7_3),.q1(G7_4),.q2(_w_940));
  bfr _b_860(.a(_w_1174),.q(_w_1175));
  spl2 G6_s_2(.a(G6_5),.q0(G6_6),.q1(G6_7));
  spl3L G6_s_1(.a(G6_2),.q0(G6_3),.q1(G6_4),.q2(_w_962));
  bfr _b_1105(.a(_w_1419),.q(G16_5));
  spl2 g178_s_0(.a(n178),.q0(n178_0),.q1(n178_1));
  bfr _b_545(.a(_w_859),.q(_w_860));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(n119_1));
  bfr _b_750(.a(_w_1064),.q(_w_1065));
  spl3L G3_s_1(.a(G3_2),.q0(G3_3),.q1(G3_4),.q2(_w_998));
  bfr _b_958(.a(_w_1272),.q(_w_1273));
  spl2 G22_s_0(.a(_w_1753),.q0(G22_0),.q1(G22_1));
  and_bi g85(.a(n84_0),.b(n66_2),.q(n85));
  or_bb g261(.a(G13_6),.b(n254_6),.q(n261));
  spl2 G11_s_2(.a(G11_5),.q0(G11_6),.q1(G11_7));
  bfr _b_1210(.a(_w_1524),.q(_w_1525));
  bfr _b_898(.a(_w_1212),.q(_w_1213));
  bfr _b_592(.a(_w_906),.q(G31_18));
  spl3L G25_s_0(.a(_w_1754),.q0(G25_0),.q1(G25_1),.q2(_w_1063));
  bfr _b_1486(.a(G28),.q(_w_1801));
  bfr _b_1014(.a(_w_1328),.q(_w_1329));
  spl3L G3_s_0(.a(G3),.q0(G3_0),.q1(G3_1),.q2(_w_1075));
  bfr _b_1125(.a(_w_1439),.q(_w_1440));
  spl2 g105_s_1(.a(n105_2),.q0(n105_3),.q1(n105_4));
  spl2 g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1));
  spl2 G4_s_3(.a(G4_8),.q0(G4_9),.q1(G4_10));
  bfr _b_751(.a(_w_1065),.q(_w_1066));
  and_bi g146(.a(G2_3),.b(n145_0),.q(n146));
  bfr _b_1231(.a(_w_1545),.q(_w_1546));
  bfr _b_647(.a(_w_961),.q(G7_5));
  spl3L g105_s_0(.a(n105),.q0(n105_0),.q1(n105_1),.q2(_w_1077));
  spl2 G19_s_0(.a(_w_1748),.q0(G19_0),.q1(_w_1083));
  spl2 G21_s_0(.a(_w_1752),.q0(_w_1084),.q1(G21_1));
  bfr _b_502(.a(_w_816),.q(_w_817));
  bfr _b_1540(.a(_w_1854),.q(_w_1852));
  bfr _b_681(.a(_w_995),.q(_w_996));
  spl3L g77_s_0(.a(n77),.q0(n77_0),.q1(n77_1),.q2(_w_1099));
  or_bb g84(.a(n82),.b(n83),.q(n84));
  bfr _b_668(.a(_w_982),.q(_w_983));
  bfr _b_1260(.a(_w_1574),.q(_w_1575));
  bfr _b_498(.a(_w_812),.q(_w_813));
  spl2 G24_s_1(.a(G24_1),.q0(_w_1102),.q1(G24_3));
  or_bb g174(.a(G28_1),.b(n172_1),.q(n174));
  spl2 g53_s_0(.a(n53),.q0(n53_0),.q1(n53_1));
  bfr _b_1273(.a(_w_1587),.q(_w_1588));
  bfr _b_861(.a(_w_1175),.q(_w_1176));
  spl2 G24_s_0(.a(G24),.q0(G24_0),.q1(G24_1));
  bfr _b_1357(.a(_w_1671),.q(_w_1672));
  spl3L G33_s_3(.a(G33_7),.q0(G33_8),.q1(G33_9),.q2(_w_1103));
  spl2 G33_s_2(.a(G33_5),.q0(G33_6),.q1(G33_7));
  bfr _b_1316(.a(_w_1630),.q(_w_1631));
  and_bi g195(.a(n193),.b(n194),.q(n195));
  bfr _b_1451(.a(_w_1765),.q(_w_1766));
  bfr _b_1393(.a(_w_1707),.q(_w_1708));
  bfr _b_1343(.a(_w_1657),.q(_w_1658));
  bfr _b_795(.a(_w_1109),.q(_w_1110));
  spl3L G33_s_0(.a(G33),.q0(G33_0),.q1(G33_1),.q2(G33_2));
  spl2 G16_s_2(.a(G16_5),.q0(G16_6),.q1(G16_7));
  and_bb g305(.a(n299_0),.b(n304_0),.q(n305));
  spl3L G16_s_0(.a(_w_1741),.q0(G16_0),.q1(G16_1),.q2(G16_2));
  bfr _b_1431(.a(_w_1745),.q(_w_1744));
  spl2 g222_s_2(.a(n222_4),.q0(n222_6),.q1(n222_7));
  bfr _b_739(.a(_w_1053),.q(_w_1054));
  or_bb g176(.a(n155),.b(n175),.q(n176));
  bfr _b_1471(.a(G27),.q(_w_1786));
  spl3L G28_s_0(.a(_w_1800),.q0(G28_0),.q1(G28_1),.q2(_w_1123));
  bfr _b_982(.a(_w_1296),.q(_w_1297));
  spl2 g222_s_1(.a(n222_3),.q0(n222_4),.q1(n222_5));
  bfr _b_918(.a(_w_1232),.q(_w_1233));
  bfr _b_559(.a(_w_873),.q(_w_874));
  spl2 G10_s_2(.a(G10_5),.q0(G10_6),.q1(G10_7));
  bfr _b_951(.a(_w_1265),.q(_w_1266));
  spl3L G10_s_0(.a(G10),.q0(G10_0),.q1(G10_1),.q2(_w_1157));
  spl2 G14_s_2(.a(G14_5),.q0(G14_6),.q1(G14_7));
  bfr _b_1534(.a(_w_1848),.q(_w_1849));
  bfr _b_569(.a(_w_883),.q(_w_884));
  spl2 G12_s_2(.a(G12_5),.q0(G12_6),.q1(G12_7));
  spl3L G4_s_2(.a(G4_5),.q0(G4_6),.q1(G4_7),.q2(_w_1183));
  bfr _b_864(.a(_w_1178),.q(_w_1179));
  and_bb g268(.a(G32_1),.b(n267_0),.q(n268));
  spl3L G1_s_1(.a(G1_2),.q0(G1_3),.q1(G1_4),.q2(_w_1206));
  bfr _b_807(.a(_w_1121),.q(_w_1122));
  bfr _b_1254(.a(_w_1568),.q(_w_1569));
  spl4L g267_s_1(.a(n267_3),.q0(n267_4),.q1(n267_5),.q2(n267_6),.q3(n267_7));
  spl4L g50_s_0(.a(n50),.q0(n50_0),.q1(n50_1),.q2(n50_2),.q3(n50_3));
  bfr _b_721(.a(_w_1035),.q(_w_1036));
  bfr _b_1049(.a(_w_1363),.q(_w_1364));
  bfr _b_535(.a(_w_849),.q(_w_850));
  and_bb g43(.a(G4_4),.b(G8_1),.q(n43));
  or_bb g182(.a(n180),.b(n181),.q(n182));
  spl2 g47_s_0(.a(n47),.q0(n47_0),.q1(n47_1));
  and_bi g191(.a(n189),.b(n190),.q(_w_1632));
  bfr _b_1222(.a(_w_1536),.q(_w_1537));
  spl2 g275_s_0(.a(n275),.q0(n275_0),.q1(n275_1));
  spl2 g198_s_0(.a(n198),.q0(n198_0),.q1(n198_1));
  spl3L g195_s_0(.a(n195),.q0(n195_0),.q1(n195_1),.q2(n195_2));
  bfr _b_1340(.a(_w_1654),.q(G1900));
  and_bb g173(.a(G28_0),.b(n172_0),.q(n173));
  spl3L G15_s_0(.a(G15),.q0(G15_0),.q1(G15_1),.q2(G15_2));
  bfr _b_1355(.a(_w_1669),.q(_w_1670));
  spl2 g203_s_2(.a(n203_3),.q0(_w_1235),.q1(n203_5));
  spl2 g161_s_0(.a(n161),.q0(n161_0),.q1(n161_1));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  bfr _b_1075(.a(_w_1389),.q(_w_1390));
  spl3L g87_s_1(.a(n87_2),.q0(n87_3),.q1(n87_4),.q2(n87_5));
  spl2 g89_s_0(.a(n89),.q0(n89_0),.q1(n89_1));
  bfr _b_1064(.a(_w_1378),.q(_w_1379));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  bfr _b_571(.a(_w_885),.q(_w_886));
  spl3L G8_s_1(.a(G8_2),.q0(G8_3),.q1(G8_4),.q2(_w_1236));
  bfr _b_730(.a(_w_1044),.q(_w_1045));
  bfr _b_1256(.a(_w_1570),.q(_w_1571));
  bfr _b_765(.a(_w_1079),.q(_w_1080));
  spl2 g95_s_0(.a(n95),.q0(n95_0),.q1(n95_1));
  or_bb g34(.a(G24_2),.b(G31_3),.q(n34));
  spl2 g38_s_0(.a(n38),.q0(n38_0),.q1(n38_1));
  bfr _b_1291(.a(_w_1605),.q(_w_1606));
  spl4L g254_s_2(.a(n254_1),.q0(n254_6),.q1(n254_7),.q2(n254_8),.q3(n254_9));
  or_bb g213(.a(G3_6),.b(n206_10),.q(n213));
  spl2 g145_s_0(.a(n145),.q0(n145_0),.q1(n145_1));
  spl4L g254_s_1(.a(n254_0),.q0(n254_2),.q1(n254_3),.q2(n254_4),.q3(n254_5));
  bfr _b_794(.a(_w_1108),.q(_w_1109));
  bfr _b_1028(.a(_w_1342),.q(_w_1343));
  spl3L G4_s_0(.a(G4),.q0(G4_0),.q1(G4_1),.q2(_w_1237));
  bfr _b_990(.a(_w_1304),.q(_w_1305));
  and_bi g322(.a(n321),.b(n320),.q(_w_1239));
  and_bb g320(.a(G26_2),.b(n267_7),.q(n320));
  bfr _b_1143(.a(_w_1457),.q(G1899));
  and_ii g319(.a(n317),.b(n318),.q(_w_1241));
  bfr _b_505(.a(_w_819),.q(_w_820));
  and_bb g314(.a(n222_2),.b(n312_1),.q(n314));
  bfr _b_546(.a(_w_860),.q(_w_861));
  or_bb g156(.a(G3_3),.b(G6_3),.q(n156));
  or_bb g313(.a(n222_1),.b(n312_0),.q(n313));
  and_bb g312(.a(G22_0),.b(G30_0),.q(_w_1242));
  bfr _b_1445(.a(_w_1759),.q(_w_1760));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(n88_1));
  and_bi g289(.a(n151_1),.b(n288),.q(n289));
  bfr _b_874(.a(_w_1188),.q(_w_1189));
  bfr _b_1281(.a(_w_1595),.q(_w_1596));
  and_bb g311(.a(n308),.b(n310),.q(_w_1265));
  or_bb g127(.a(G23_2),.b(G31_0),.q(n127));
  and_bi g310(.a(n219_1),.b(n309),.q(n310));
  bfr _b_1123(.a(_w_1437),.q(_w_1438));
  and_bb g196(.a(n178_2),.b(n195_0),.q(n196));
  and_bi g78(.a(n35_2),.b(n77_0),.q(n78));
  and_bb g309(.a(n105_3),.b(n87_6),.q(_w_1274));
  or_bi g307(.a(n305),.b(n306),.q(_w_1280));
  bfr _b_1395(.a(_w_1709),.q(_w_1710));
  bfr _b_1151(.a(_w_1465),.q(_w_1466));
  bfr _b_1139(.a(_w_1453),.q(G5_5));
  or_bb g219(.a(G30_1),.b(G33_9),.q(n219));
  bfr _b_1530(.a(_w_1844),.q(_w_1845));
  bfr _b_1401(.a(_w_1715),.q(_w_1716));
  bfr _b_692(.a(_w_1006),.q(_w_1007));
  bfr _b_1063(.a(_w_1377),.q(_w_1378));
  spl2 g219_s_0(.a(n219),.q0(n219_0),.q1(n219_1));
  bfr _b_543(.a(_w_857),.q(_w_858));
  spl2 g200_s_0(.a(n200),.q0(n200_0),.q1(_w_1281));
  spl2 g168_s_0(.a(n168),.q0(n168_0),.q1(n168_1));
  and_bb g300(.a(G21_0),.b(G29_0),.q(_w_1282));
  or_bb g92(.a(n90),.b(n91),.q(n92));
  and_bb g299(.a(n199_1),.b(n56_2),.q(_w_1290));
  spl2 g171_s_0(.a(n171),.q0(n171_0),.q1(_w_1300));
  spl2 G23_s_0(.a(G23),.q0(G23_0),.q1(G23_1));
  and_bi g315(.a(n313),.b(n314),.q(n315));
  and_bb g298(.a(n203_9),.b(n297),.q(_w_1318));
  or_bb g297(.a(n125_1),.b(n296),.q(n297));
  bfr _b_1484(.a(_w_1798),.q(_w_1799));
  and_bi g294(.a(n203_8),.b(n293),.q(_w_1319));
  and_bb g292(.a(n267_5),.b(n291),.q(n292));
  and_bi g158(.a(n156),.b(n157),.q(n158));
  bfr _b_580(.a(_w_894),.q(_w_895));
  bfr _b_797(.a(_w_1111),.q(_w_1112));
  bfr _b_489(.a(_w_803),.q(_w_804));
  bfr _b_634(.a(_w_948),.q(_w_949));
  bfr _b_675(.a(_w_989),.q(_w_990));
  bfr _b_1339(.a(_w_1653),.q(_w_1654));
  and_bi g58(.a(n57_0),.b(G9_3),.q(n58));
  bfr _b_908(.a(_w_1222),.q(_w_1223));
  and_bb g190(.a(n188_1),.b(n87_1),.q(n190));
  bfr _b_1386(.a(_w_1700),.q(_w_1701));
  bfr _b_1244(.a(_w_1558),.q(_w_1559));
  bfr _b_873(.a(_w_1187),.q(_w_1188));
  or_bb g105(.a(n103),.b(n104),.q(n105));
  and_bi g38(.a(n36),.b(n37),.q(n38));
  bfr _b_1195(.a(_w_1509),.q(_w_1510));
  spl3L G2_s_1(.a(G2_2),.q0(G2_3),.q1(G2_4),.q2(_w_1163));
  or_bb g316(.a(G33_14),.b(n315),.q(n316));
  and_bi g155(.a(n154),.b(n153),.q(n155));
  spl2 g206_s_1(.a(n206_3),.q0(n206_4),.q1(n206_5));
  bfr _b_992(.a(_w_1306),.q(_w_1307));
  bfr _b_512(.a(_w_826),.q(_w_827));
  bfr _b_503(.a(_w_817),.q(_w_818));
  spl2 g99_s_0(.a(n99),.q0(n99_0),.q1(n99_1));
  spl2 g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1));
  bfr _b_703(.a(_w_1017),.q(_w_1018));
  bfr _b_744(.a(_w_1058),.q(_w_1059));
  and_bi g147(.a(n145_1),.b(G2_4),.q(n147));
  and_bb g240(.a(G6_7),.b(n235_5),.q(n240));
  and_bb g39(.a(G5_0),.b(n38_0),.q(n39));
  bfr _b_1145(.a(_w_1459),.q(_w_1460));
  or_bb g151(.a(n149),.b(n150),.q(n151));
  and_bi g318(.a(n316_1),.b(n311_1),.q(n318));
  bfr _b_880(.a(_w_1194),.q(_w_1195));
  bfr _b_1130(.a(_w_1444),.q(_w_1445));
  bfr _b_890(.a(_w_1204),.q(_w_1205));
  and_bb g140(.a(n108_2),.b(n139_0),.q(n140));
  or_bb g137(.a(n133_0),.b(n136_0),.q(n137));
  spl2 G29_s_0(.a(_w_1814),.q0(G29_0),.q1(G29_1));
  spl2 g133_s_0(.a(n133),.q0(n133_0),.q1(n133_1));
  or_bb g154(.a(G27_1),.b(n152_1),.q(n154));
  spl3L G27_s_0(.a(_w_1785),.q0(G27_0),.q1(G27_1),.q2(_w_1321));
  and_bi g200(.a(G24_3),.b(G23_3),.q(_w_1334));
  spl2 g203_s_0(.a(n203),.q0(n203_0),.q1(_w_1347));
  bfr _b_588(.a(_w_902),.q(n74_2));
  bfr _b_1083(.a(_w_1397),.q(_w_1398));
  spl2 g35_s_1(.a(n35_1),.q0(n35_2),.q1(_w_1358));
  and_bi g90(.a(n89_0),.b(G1_3),.q(n90));
  spl2 g203_s_1(.a(n203_1),.q0(n203_2),.q1(n203_3));
  and_bi g95(.a(n93),.b(n94),.q(n95));
  or_bb g160(.a(G8_7),.b(n158_1),.q(n160));
  bfr _b_491(.a(_w_805),.q(_w_806));
  and_bi g152(.a(n151_0),.b(G31_7),.q(n152));
  bfr _b_552(.a(_w_866),.q(_w_867));
  or_bb g130(.a(n126_1),.b(n128_1),.q(n130));
  bfr _b_967(.a(_w_1281),.q(n200_1));
  bfr _b_540(.a(_w_854),.q(_w_855));
  and_bi g61(.a(G10_0),.b(G15_0),.q(n61));
  or_bb g242(.a(G7_6),.b(n235_6),.q(n242));
  bfr _b_957(.a(_w_1271),.q(_w_1272));
  bfr _b_495(.a(_w_809),.q(_w_810));
  and_bi g248(.a(n234_0),.b(n221_1),.q(n248));
  and_bb g129(.a(n126_0),.b(n128_0),.q(n129));
  or_bb g53(.a(n51),.b(n52),.q(n53));
  bfr _b_1117(.a(_w_1431),.q(n35));
  and_bb g187(.a(n185_1),.b(n50_3),.q(n187));
  and_bb g128(.a(G19_1),.b(n127_0),.q(_w_1387));
  or_bb g193(.a(G25_0),.b(n192_0),.q(n193));
  bfr _b_926(.a(_w_1240),.q(G1908));
  or_bb g126(.a(G31_6),.b(n125_0),.q(n126));
  spl3L G16_s_1(.a(G16_2),.q0(G16_3),.q1(G16_4),.q2(_w_1397));
  bfr _b_1531(.a(_w_1845),.q(_w_1846));
  and_bi g125(.a(n124),.b(n123),.q(n125));
  bfr _b_554(.a(_w_868),.q(_w_869));
  bfr _b_696(.a(_w_1010),.q(_w_1011));
  and_bb g123(.a(n116_0),.b(n122_0),.q(n123));
  or_bb g119(.a(n117),.b(n118),.q(n119));
  bfr _b_844(.a(_w_1158),.q(_w_1159));
  bfr _b_1318(.a(_w_1632),.q(_w_1633));
  and_bb g256(.a(G11_7),.b(n254_3),.q(n256));
  and_bi g118(.a(G7_4),.b(G4_7),.q(n118));
  bfr _b_1265(.a(_w_1579),.q(_w_1580));
  bfr _b_1212(.a(_w_1526),.q(_w_1527));
  bfr _b_585(.a(_w_899),.q(_w_900));
  spl2 G30_s_0(.a(_w_1830),.q0(G30_0),.q1(_w_1108));
  spl2 g312_s_0(.a(n312),.q0(n312_0),.q1(n312_1));
  and_bi g250(.a(n248_1),.b(G9_7),.q(n250));
  bfr _b_853(.a(_w_1167),.q(_w_1168));
  spl2 g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1));
  spl2 G23_s_1(.a(G23_1),.q0(G23_2),.q1(G23_3));
  bfr _b_842(.a(_w_1156),.q(G10_5));
  bfr _b_515(.a(_w_829),.q(_w_830));
  and_bi g234(.a(n233),.b(n78_1),.q(n234));
  and_bi g111(.a(n110_0),.b(G13_3),.q(n111));
  and_bi g110(.a(G20_0),.b(n109_0),.q(n110));
  bfr _b_605(.a(_w_919),.q(_w_920));
  and_bi g222(.a(n198_1),.b(n221_0),.q(n222));
  or_bb g220(.a(n201_1),.b(n219_0),.q(n220));
  and_bi g150(.a(n142_1),.b(n148_1),.q(n150));
  or_bb g63(.a(n61),.b(n62),.q(n63));
  or_bb g164(.a(G12_4),.b(n63_3),.q(n164));
  bfr _b_768(.a(_w_1082),.q(n105_2));
  and_bi g79(.a(G13_0),.b(G11_0),.q(n79));
  or_bb g113(.a(n111),.b(n112),.q(n113));
  or_bb g201(.a(G31_13),.b(n200_0),.q(n201));
  spl2 g57_s_0(.a(n57),.q0(n57_0),.q1(n57_1));
  and_bi g56(.a(n54),.b(n55),.q(n56));
  bfr _b_1498(.a(_w_1812),.q(_w_1813));
  and_bi g249(.a(G9_6),.b(n248_0),.q(n249));
  bfr _b_1482(.a(_w_1796),.q(_w_1797));
  bfr _b_1203(.a(_w_1517),.q(G8_8));
  bfr _b_607(.a(_w_921),.q(_w_922));
  bfr _b_1085(.a(_w_1399),.q(_w_1400));
  bfr _b_1042(.a(_w_1356),.q(_w_1357));
  bfr _b_1043(.a(_w_1357),.q(n203_1));
  and_bb g135(.a(G11_4),.b(G15_4),.q(n135));
  or_bb g96(.a(n87_3),.b(n95_0),.q(n96));
  bfr _b_1414(.a(_w_1728),.q(G17_1));
  or_bb g73(.a(G31_11),.b(n72_0),.q(n73));
  and_bi g114(.a(n113_0),.b(n108_0),.q(n114));
  bfr _b_551(.a(_w_865),.q(_w_866));
  and_bi g62(.a(G15_1),.b(G10_1),.q(n62));
  bfr _b_1077(.a(_w_1391),.q(_w_1392));
  spl2 G3_s_2(.a(G3_5),.q0(G3_6),.q1(G3_7));
  bfr _b_1476(.a(_w_1790),.q(_w_1791));
  bfr _b_1048(.a(_w_1362),.q(_w_1363));
  bfr _b_530(.a(_w_844),.q(_w_845));
  spl2 g87_s_2(.a(n87_5),.q0(n87_6),.q1(n87_7));
  spl3L G9_s_0(.a(_w_1855),.q0(G9_0),.q1(G9_1),.q2(_w_1615));
  and_bi g254(.a(n253),.b(n221_2),.q(n254));
  bfr _b_482(.a(_w_796),.q(_w_797));
  spl2 G33_s_4(.a(G33_10),.q0(G33_11),.q1(_w_1458));
  or_bb g108(.a(n106),.b(n107),.q(n108));
  and_bi g197(.a(n177_0),.b(n196),.q(n197));
  bfr _b_1237(.a(_w_1551),.q(_w_1552));
  or_bb g203(.a(G32_0),.b(G33_6),.q(n203));
  bfr _b_713(.a(_w_1027),.q(_w_1028));
  bfr _b_820(.a(_w_1134),.q(_w_1135));
  or_bb g141(.a(n108_3),.b(n139_1),.q(n141));
  and_bi g59(.a(G9_4),.b(n57_1),.q(n59));
  bfr _b_508(.a(_w_822),.q(_w_823));
  bfr _b_1310(.a(_w_1624),.q(_w_1625));
  or_bb g93(.a(n41_0),.b(n92_0),.q(n93));
  bfr _b_562(.a(_w_876),.q(_w_877));
  spl2 G8_s_3(.a(G8_8),.q0(G8_9),.q1(G8_10));
  bfr _b_519(.a(_w_833),.q(_w_834));
  bfr _b_937(.a(_w_1251),.q(_w_1252));
  or_bb g45(.a(G2_0),.b(G3_0),.q(n45));
  bfr _b_1266(.a(_w_1580),.q(G33_5));
  bfr _b_1172(.a(_w_1486),.q(_w_1487));
  or_bb g49(.a(G1_1),.b(n47_1),.q(n49));
  and_bb g302(.a(n206_2),.b(n300_1),.q(n302));
  bfr _b_1529(.a(_w_1843),.q(_w_1844));
  spl2 g92_s_0(.a(n92),.q0(n92_0),.q1(n92_1));
  bfr _b_733(.a(_w_1047),.q(_w_1048));
  bfr _b_1434(.a(G19),.q(_w_1749));
  spl2 g98_s_0(.a(n98),.q0(n98_0),.q1(_w_1022));
  or_bb g186(.a(n185_0),.b(n50_2),.q(n186));
  spl2 g162_s_0(.a(n162),.q0(n162_0),.q1(n162_1));
  or_bb g226(.a(G15_6),.b(n222_8),.q(n226));
  and_bi g143(.a(G5_3),.b(G8_3),.q(n143));
  bfr _b_1181(.a(_w_1495),.q(_w_1496));
  bfr _b_1103(.a(_w_1417),.q(_w_1418));
  and_bb g265(.a(G14_7),.b(n254_9),.q(n265));
  or_bb g207(.a(G1_6),.b(n206_6),.q(n207));
  bfr _b_769(.a(_w_1083),.q(G19_1));
  bfr _b_1202(.a(_w_1516),.q(_w_1517));
  bfr _b_672(.a(_w_986),.q(_w_987));
  or_bb g124(.a(n116_1),.b(n122_1),.q(n124));
  or_bb g245(.a(G8_9),.b(n235_8),.q(n245));
  bfr _b_1524(.a(_w_1838),.q(_w_1839));
  spl4L g222_s_3(.a(n222_5),.q0(n222_8),.q1(n222_9),.q2(n222_10),.q3(n222_11));
  and_bi g47(.a(n45),.b(n46),.q(n47));
  and_bi g162(.a(G19_0),.b(n109_1),.q(_w_1493));
  spl4L g206_s_0(.a(n206),.q0(n206_0),.q1(n206_1),.q2(n206_2),.q3(n206_3));
  bfr _b_1488(.a(_w_1802),.q(_w_1803));
  bfr _b_1333(.a(_w_1647),.q(_w_1648));
  bfr _b_712(.a(_w_1026),.q(_w_1027));
  bfr _b_589(.a(_w_903),.q(n35_1));
  bfr _b_932(.a(_w_1246),.q(_w_1247));
  and_bi g75(.a(n73_0),.b(n74_0),.q(n75));
  spl2 G1_s_2(.a(G1_5),.q0(G1_6),.q1(G1_7));
  bfr _b_1165(.a(_w_1479),.q(_w_1480));
  or_bi g218(.a(n217),.b(n216),.q(_w_1495));
  and_bi g57(.a(G21_1),.b(G33_3),.q(n57));
  bfr _b_1457(.a(_w_1771),.q(_w_1772));
  or_bb g122(.a(n120),.b(n121),.q(n122));
  and_bi g86(.a(n66_3),.b(n84_1),.q(n86));
  and_bi g321(.a(n203_2),.b(n98_1),.q(n321));
  and_bi g161(.a(n160),.b(n159),.q(n161));
  and_bi g291(.a(G28_2),.b(G31_16),.q(n291));
  bfr _b_1313(.a(_w_1627),.q(G18_1));
  or_bi g241(.a(n240),.b(n239),.q(_w_1628));
  bfr _b_631(.a(_w_945),.q(_w_946));
  or_bb g40(.a(G5_2),.b(n38_1),.q(n40));
  and_bb g281(.a(G25_2),.b(n267_2),.q(n281));
  bfr _b_1428(.a(_w_1742),.q(_w_1743));
  bfr _b_1376(.a(_w_1690),.q(G1891));
  bfr _b_1039(.a(_w_1353),.q(_w_1354));
  or_bb g77(.a(n75),.b(n76),.q(n77));
  bfr _b_1149(.a(_w_1463),.q(_w_1464));
  bfr _b_1086(.a(_w_1400),.q(_w_1401));
  bfr _b_1170(.a(_w_1484),.q(_w_1485));
  or_bb g42(.a(G4_3),.b(G8_0),.q(n42));
  and_bi g41(.a(n40),.b(n39),.q(n41));
  bfr _b_527(.a(_w_841),.q(_w_842));
  bfr _b_1437(.a(_w_1751),.q(_w_1750));
  spl2 g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1));
  spl3L G4_s_1(.a(G4_2),.q0(G4_3),.q1(G4_4),.q2(G4_5));
  and_bi g171(.a(n169),.b(n170),.q(n171));
  bfr _b_1255(.a(_w_1569),.q(_w_1570));
  spl3L G8_s_2(.a(G8_5),.q0(G8_6),.q1(G8_7),.q2(_w_1498));
  bfr _b_615(.a(_w_929),.q(_w_930));
  bfr _b_722(.a(_w_1036),.q(_w_1037));
  bfr _b_831(.a(_w_1145),.q(_w_1146));
  bfr _b_500(.a(_w_814),.q(_w_815));
  and_bb g237(.a(G5_7),.b(n235_3),.q(n237));
  spl2 g126_s_0(.a(n126),.q0(n126_0),.q1(n126_1));
  or_bb g258(.a(G12_6),.b(n254_4),.q(n258));
  spl2 g81_s_0(.a(n81),.q0(n81_0),.q1(n81_1));
  bfr _b_1435(.a(_w_1749),.q(_w_1748));
  and_bi g133(.a(G18_0),.b(n88_1),.q(n133));
  bfr _b_1057(.a(_w_1371),.q(_w_1372));
  and_bb g246(.a(G8_10),.b(n235_9),.q(n246));
  bfr _b_1121(.a(_w_1435),.q(_w_1436));
  bfr _b_695(.a(_w_1009),.q(_w_1010));
  and_bb g37(.a(G6_1),.b(G7_1),.q(n37));
  spl2 g248_s_0(.a(n248),.q0(n248_0),.q1(n248_1));
  bfr _b_507(.a(_w_821),.q(_w_822));
  bfr _b_1115(.a(_w_1429),.q(_w_1430));
  spl3L g73_s_0(.a(n73),.q0(n73_0),.q1(n73_1),.q2(_w_1518));
  and_bi g102(.a(n100),.b(n101),.q(n102));
  bfr _b_1327(.a(_w_1641),.q(_w_1642));
  bfr _b_1280(.a(_w_1594),.q(_w_1595));
  spl2 G2_s_2(.a(G2_5),.q0(G2_6),.q1(G2_7));
  and_bb g46(.a(G2_1),.b(G3_1),.q(n46));
  spl2 g113_s_0(.a(n113),.q0(n113_0),.q1(n113_1));
  bfr _b_999(.a(_w_1313),.q(_w_1314));
  and_bi g165(.a(n164),.b(n163),.q(n165));
  spl3L g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1),.q2(_w_1531));
  bfr _b_1150(.a(_w_1464),.q(_w_1465));
  spl2 G31_s_4(.a(G31_10),.q0(G31_11),.q1(G31_12));
  and_bi g64(.a(n63_0),.b(G16_0),.q(n64));
  or_bb g66(.a(n64),.b(n65),.q(n66));
  and_bb g35(.a(G18_1),.b(n34_1),.q(_w_1420));
  or_bb g210(.a(G2_6),.b(n206_8),.q(n210));
  and_bb g74(.a(G17_1),.b(n34_0),.q(_w_1545));
  or_bb g269(.a(n178_0),.b(n35_0),.q(n269));
  and_bi g287(.a(G27_2),.b(G31_15),.q(n287));
  bfr _b_496(.a(_w_810),.q(n191_1));
  or_bb g99(.a(G31_5),.b(n98_0),.q(n99));
  bfr _b_595(.a(_w_909),.q(_w_910));
  bfr _b_1052(.a(_w_1366),.q(_w_1367));
  spl3L G11_s_1(.a(G11_2),.q0(G11_3),.q1(G11_4),.q2(_w_1038));
  and_bb g208(.a(G1_7),.b(n206_7),.q(n208));
  bfr _b_758(.a(_w_1072),.q(_w_1073));
  and_bi g103(.a(G9_0),.b(G14_3),.q(n103));
  or_bb g72(.a(n70),.b(n71),.q(n72));
  bfr _b_533(.a(_w_847),.q(_w_848));
  bfr _b_493(.a(_w_807),.q(_w_808));
  spl2 g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1));
  bfr _b_1452(.a(_w_1766),.q(_w_1767));
  bfr _b_1051(.a(_w_1365),.q(_w_1366));
  or_bb g283(.a(n191_1),.b(n282),.q(n283));
  or_bb g36(.a(G6_0),.b(G7_0),.q(n36));
  spl2 G31_s_0(.a(_w_1831),.q0(G31_0),.q1(G31_1));
  bfr _b_899(.a(_w_1213),.q(_w_1214));
  and_bi g180(.a(G4_0),.b(G14_0),.q(n180));
  spl3L g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1),.q2(_w_857));
  spl2 g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1));
  spl3L g41_s_0(.a(n41),.q0(n41_0),.q1(n41_1),.q2(_w_1386));
  and_bi g184(.a(n182_1),.b(n179_1),.q(n184));
  bfr _b_1040(.a(_w_1354),.q(_w_1355));
  or_bb g308(.a(n105_4),.b(n87_7),.q(_w_1556));
  bfr _b_731(.a(_w_1045),.q(_w_1046));
  and_ii g251(.a(n249),.b(n250),.q(_w_1563));
  and_bi g112(.a(G13_4),.b(n110_1),.q(n112));
  or_bb g270(.a(n195_1),.b(n269),.q(n270));
  and_bi g50(.a(n49),.b(n48),.q(n50));
  spl4L g108_s_0(.a(n108),.q0(n108_0),.q1(n108_1),.q2(n108_2),.q3(n108_3));
  and_bb g296(.a(n267_6),.b(n295),.q(n296));
  or_bb g168(.a(n166),.b(n167),.q(n168));
  and_bi g80(.a(G11_1),.b(G13_1),.q(n80));
  spl2 G31_s_3(.a(G31_8),.q0(G31_9),.q1(G31_10));
  spl3L G33_s_1(.a(G33_2),.q0(G33_3),.q1(G33_4),.q2(_w_1568));
  or_bb g134(.a(G11_3),.b(G15_3),.q(n134));
  spl2 g72_s_0(.a(n72),.q0(n72_0),.q1(_w_1581));
  and_bi g89(.a(G17_0),.b(n88_0),.q(n89));
  bfr _b_652(.a(_w_966),.q(_w_967));
  and_bi g65(.a(G16_1),.b(n63_1),.q(n65));
  and_bb g163(.a(G12_3),.b(n63_2),.q(n163));
  and_bi g166(.a(n162_0),.b(n165_0),.q(n166));
  bfr _b_959(.a(_w_1273),.q(n311));
  and_bi g167(.a(n165_1),.b(n162_1),.q(n167));
  bfr _b_1045(.a(_w_1359),.q(n35_3));
  spl3L G26_s_0(.a(_w_1770),.q0(G26_0),.q1(G26_1),.q2(_w_1601));
  bfr _b_821(.a(_w_1135),.q(_w_1136));
  or_bb g306(.a(n299_1),.b(n304_1),.q(n306));
  bfr _b_1439(.a(G22),.q(_w_1753));
  bfr _b_1363(.a(_w_1677),.q(G12_5));
  bfr _b_1288(.a(_w_1602),.q(_w_1603));
  bfr _b_1091(.a(_w_1405),.q(_w_1406));
  or_bb g169(.a(n161_0),.b(n168_0),.q(n169));
  bfr _b_525(.a(_w_839),.q(_w_840));
  bfr _b_547(.a(_w_861),.q(_w_862));
  spl2 G33_s_5(.a(G33_12),.q0(G33_13),.q1(G33_14));
  and_bb g170(.a(n161_1),.b(n168_1),.q(n170));
  spl3L G14_s_0(.a(G14),.q0(G14_0),.q1(G14_1),.q2(G14_2));
  bfr _b_1269(.a(_w_1583),.q(_w_1584));
  bfr _b_1087(.a(_w_1401),.q(_w_1402));
  bfr _b_1218(.a(_w_1532),.q(_w_1533));
  and_bi g290(.a(n203_7),.b(n289),.q(_w_1597));
  and_bi g285(.a(n203_6),.b(n284),.q(n285));
  spl4L g206_s_2(.a(n206_4),.q0(n206_6),.q1(n206_7),.q2(n206_8),.q3(n206_9));
  spl2 G7_s_2(.a(G7_5),.q0(G7_6),.q1(G7_7));
  spl2 G15_s_2(.a(G15_5),.q0(G15_6),.q1(G15_7));
  bfr _b_1081(.a(_w_1395),.q(_w_1396));
  spl3L G8_s_0(.a(_w_1852),.q0(G8_0),.q1(G8_1),.q2(G8_2));
  bfr _b_1197(.a(_w_1511),.q(_w_1512));
  bfr _b_985(.a(_w_1299),.q(n299));
  bfr _b_1257(.a(_w_1571),.q(_w_1572));
  and_bb g252(.a(n197_1),.b(n35_3),.q(n252));
  bfr _b_521(.a(_w_835),.q(_w_836));
  bfr _b_841(.a(_w_1155),.q(_w_1156));
  and_bi g179(.a(G22_1),.b(G33_4),.q(n179));
  bfr _b_1344(.a(_w_1658),.q(_w_1659));
  and_bi g317(.a(n311_0),.b(n316_0),.q(n317));
  bfr _b_650(.a(_w_964),.q(_w_965));
  or_bi g257(.a(n256),.b(n255),.q(_w_1616));
  bfr _b_915(.a(_w_1229),.q(_w_1230));
  and_bi g131(.a(n130),.b(n129),.q(n131));
  or_bb g216(.a(G4_9),.b(n206_12),.q(n216));
  or_bi g228(.a(n227),.b(n226),.q(_w_1733));
  bfr _b_777(.a(_w_1091),.q(_w_1092));
  spl3L G2_s_0(.a(G2),.q0(G2_0),.q1(G2_1),.q2(_w_1620));
  spl2 G31_s_7(.a(G31_18),.q0(G31_19),.q1(G31_20));
  or_bb g185(.a(n183),.b(n184),.q(n185));
  bfr _b_1442(.a(_w_1756),.q(_w_1757));
  spl2 G18_s_0(.a(_w_1746),.q0(G18_0),.q1(_w_1626));
  or_bb g273(.a(G33_11),.b(n272),.q(_w_1634));
  bfr _b_1092(.a(_w_1406),.q(_w_1407));
  and_bb g157(.a(G3_4),.b(G6_4),.q(n157));
  bfr _b_772(.a(_w_1086),.q(_w_1087));
  or_bb g199(.a(G29_1),.b(G33_8),.q(n199));
  or_bb g202(.a(n199_0),.b(n201_0),.q(n202));
  bfr _b_1175(.a(_w_1489),.q(_w_1490));
  bfr _b_660(.a(_w_974),.q(_w_975));
  and_bi g198(.a(n197_0),.b(n78_0),.q(n198));
  bfr _b_688(.a(_w_1002),.q(_w_1003));
  or_bb g204(.a(n200_1),.b(n203_0),.q(n204));
  bfr _b_531(.a(_w_845),.q(_w_846));
  bfr _b_928(.a(_w_1242),.q(_w_1243));
  bfr _b_1532(.a(_w_1846),.q(_w_1832));
  bfr _b_1464(.a(_w_1778),.q(_w_1779));
  bfr _b_1309(.a(_w_1623),.q(_w_1624));
  spl3L g221_s_0(.a(n221),.q0(n221_0),.q1(n221_1),.q2(n221_2));
  and_bi g82(.a(G12_0),.b(n81_0),.q(n82));
  or_bb g301(.a(n206_1),.b(n300_0),.q(n301));
  bfr _b_943(.a(_w_1257),.q(_w_1258));
  and_bi g71(.a(n69_1),.b(n56_1),.q(n71));
  bfr _b_1112(.a(_w_1426),.q(_w_1427));
  and_bi g206(.a(n198_0),.b(n205_0),.q(n206));
  bfr _b_594(.a(_w_908),.q(_w_909));
  and_bi g106(.a(n105_0),.b(G16_3),.q(n106));
  and_bi g115(.a(n108_1),.b(n113_1),.q(n115));
  spl3L G13_s_1(.a(G13_2),.q0(G13_3),.q1(G13_4),.q2(_w_870));
  and_bb g211(.a(G2_7),.b(n206_9),.q(n211));
  bfr _b_1358(.a(_w_1672),.q(_w_1673));
  bfr _b_706(.a(_w_1020),.q(_w_1021));
  and_bi g70(.a(n56_0),.b(n69_0),.q(n70));
  bfr _b_1236(.a(_w_1550),.q(_w_1551));
  and_bi g67(.a(n66_0),.b(n60_0),.q(n67));
  and_bb g214(.a(G3_7),.b(n206_11),.q(n214));
  bfr _b_1239(.a(_w_1553),.q(_w_1554));
  bfr _b_612(.a(_w_926),.q(_w_927));
  spl4L g222_s_0(.a(n222),.q0(n222_0),.q1(n222_1),.q2(n222_2),.q3(n222_3));
  or_bi g225(.a(n224),.b(n223),.q(_w_1649));
  bfr _b_1056(.a(_w_1370),.q(_w_1371));
  spl4L G12_s_1(.a(G12_1),.q0(G12_2),.q1(G12_3),.q2(G12_4),.q3(_w_1655));
  and_bb g217(.a(G4_10),.b(n206_13),.q(n217));
  spl3L G13_s_0(.a(G13),.q0(G13_0),.q1(G13_1),.q2(_w_829));
  spl3L g87_s_0(.a(n87),.q0(n87_0),.q1(n87_1),.q2(n87_2));
  or_bb g116(.a(n114),.b(n115),.q(n116));
  bfr _b_553(.a(_w_867),.q(_w_868));
  or_bi g215(.a(n214),.b(n213),.q(_w_1646));
  bfr _b_790(.a(_w_1104),.q(_w_1105));
  and_bb g221(.a(n204_1),.b(n220),.q(_w_1678));
  bfr _b_1421(.a(_w_1735),.q(G1889));
  bfr _b_1164(.a(_w_1478),.q(_w_1479));
  bfr _b_718(.a(_w_1032),.q(_w_1033));
  or_bb g229(.a(G16_6),.b(n222_10),.q(n229));
  spl2 g41_s_1(.a(n41_2),.q0(n41_3),.q1(n41_4));
  or_bb g223(.a(G10_6),.b(n222_6),.q(n223));
  bfr _b_829(.a(_w_1143),.q(_w_1144));
  bfr _b_609(.a(_w_923),.q(_w_924));
  bfr _b_1061(.a(_w_1375),.q(_w_1376));
  and_bi g277(.a(n72_1),.b(n276),.q(n277));
  and_bb g224(.a(G10_7),.b(n222_7),.q(n224));
  bfr _b_1100(.a(_w_1414),.q(_w_1415));
  and_bb g227(.a(G15_7),.b(n222_9),.q(n227));
  spl2 g84_s_0(.a(n84),.q0(n84_0),.q1(n84_1));
  bfr _b_944(.a(_w_1258),.q(_w_1259));
  bfr _b_970(.a(_w_1284),.q(_w_1285));
  or_bi g247(.a(n246),.b(n245),.q(_w_1683));
  and_bi g121(.a(n119_1),.b(G10_4),.q(n121));
  spl3L G11_s_0(.a(G11),.q0(G11_0),.q1(G11_1),.q2(G11_2));
  or_bi g238(.a(n237),.b(n236),.q(_w_1687));
  or_bi g212(.a(n211),.b(n210),.q(_w_1643));
  spl2 g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1));
  or_bi g231(.a(n230),.b(n229),.q(_w_1691));
  bfr _b_487(.a(_w_801),.q(_w_802));
  bfr _b_1067(.a(_w_1381),.q(_w_1382));
  and_bi g232(.a(n178_3),.b(n195_2),.q(_w_1694));
  and_bb g233(.a(n177_2),.b(n232),.q(n233));
  or_bb g304(.a(G33_13),.b(n303),.q(n304));
  bfr _b_1018(.a(_w_1332),.q(_w_1333));
  and_bi g149(.a(n148_0),.b(n142_0),.q(n149));
  bfr _b_738(.a(_w_1052),.q(_w_1053));
  and_bi g235(.a(n234_1),.b(n205_1),.q(n235));
  bfr _b_1069(.a(_w_1383),.q(_w_1384));
  spl3L G6_s_0(.a(_w_1850),.q0(G6_0),.q1(G6_1),.q2(_w_1320));
  bfr _b_693(.a(_w_1007),.q(_w_1008));
  and_bb g243(.a(G7_7),.b(n235_7),.q(n243));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(n179_1));
  and_bi g177(.a(n132),.b(n176),.q(n177));
  and_bi g183(.a(n179_0),.b(n182_0),.q(n183));
  and_bb g101(.a(G26_1),.b(n99_1),.q(n101));
  or_bi g260(.a(n259),.b(n258),.q(_w_1699));
  and_bi g120(.a(G10_3),.b(n119_0),.q(n120));
  and_bb g262(.a(G13_7),.b(n254_7),.q(n262));
  or_bb g236(.a(G5_6),.b(n235_2),.q(n236));
  bfr _b_1481(.a(_w_1795),.q(_w_1796));
  or_bi g263(.a(n262),.b(n261),.q(_w_1703));
  bfr _b_657(.a(_w_971),.q(_w_972));
  bfr _b_1047(.a(_w_1361),.q(_w_1362));
  bfr _b_1188(.a(_w_1502),.q(_w_1503));
  bfr _b_481(.a(_w_795),.q(_w_796));
  bfr _b_565(.a(_w_879),.q(_w_880));
  bfr _b_1517(.a(G31),.q(_w_1831));
  or_bb g264(.a(G14_6),.b(n254_8),.q(n264));
  spl3L G31_s_1(.a(G31_1),.q0(_w_1707),.q1(G31_3),.q2(_w_1717));
  bfr _b_971(.a(_w_1285),.q(_w_1286));
  and_bb g205(.a(n202),.b(n204_0),.q(_w_1640));
  bfr _b_966(.a(_w_1280),.q(G1906));
  or_bb g60(.a(n58),.b(n59),.q(n60));
  or_bb g267(.a(n206_0),.b(n222_0),.q(n267));
  or_bb g109(.a(G23_0),.b(G33_1),.q(n109));
  bfr _b_532(.a(_w_846),.q(_w_847));
  and_bb g272(.a(n177_3),.b(n271),.q(n272));
  bfr _b_616(.a(_w_930),.q(_w_931));
  bfr _b_492(.a(_w_806),.q(_w_807));
  and_bb g275(.a(n267_1),.b(n74_2),.q(n275));
  and_bi g104(.a(G14_4),.b(G9_1),.q(n104));
  bfr _b_646(.a(_w_960),.q(_w_961));
  spl2 g148_s_0(.a(n148),.q0(n148_0),.q1(n148_1));
  and_bi g278(.a(n275_1),.b(n73_2),.q(n278));
  spl2 g205_s_0(.a(n205),.q0(n205_0),.q1(n205_1));
  bfr _b_1093(.a(_w_1407),.q(_w_1408));
  and_bi g280(.a(n279),.b(n277),.q(G1901));
  bfr _b_1292(.a(_w_1606),.q(_w_1607));
  bfr _b_520(.a(_w_834),.q(_w_835));
  and_bi g68(.a(n60_1),.b(n66_1),.q(n68));
  bfr _b_855(.a(_w_1169),.q(_w_1170));
  spl2 G17_s_0(.a(_w_1744),.q0(G17_0),.q1(_w_1727));
  or_bb g69(.a(n67),.b(n68),.q(_w_1730));
  and_bb g286(.a(n283),.b(n285),.q(G1902));
  and_bb g55(.a(n41_4),.b(n53_1),.q(n55));
  bfr _b_541(.a(_w_855),.q(_w_856));
  bfr _b_1527(.a(_w_1841),.q(_w_1842));
  bfr _b_1518(.a(G32),.q(_w_1833));
  and_bi g282(.a(n281_0),.b(G31_20),.q(n282));
  bfr _b_542(.a(_w_856),.q(G14_5));
  or_bb g100(.a(G26_0),.b(n99_0),.q(n100));
  bfr _b_544(.a(_w_858),.q(_w_859));
  bfr _b_665(.a(_w_979),.q(_w_980));
  bfr _b_786(.a(_w_1100),.q(_w_1101));
  bfr _b_833(.a(_w_1147),.q(_w_1148));
  bfr _b_549(.a(_w_863),.q(_w_864));
  bfr _b_917(.a(_w_1231),.q(_w_1232));
  and_bb g178(.a(G20_1),.b(n127_1),.q(_w_1463));
  bfr _b_550(.a(_w_864),.q(_w_865));
  bfr _b_555(.a(_w_869),.q(n128_2));
  bfr _b_1502(.a(_w_1816),.q(_w_1817));
  bfr _b_557(.a(_w_871),.q(_w_872));
  spl2 g158_s_0(.a(n158),.q0(n158_0),.q1(n158_1));
  bfr _b_558(.a(_w_872),.q(_w_873));
  bfr _b_560(.a(_w_874),.q(_w_875));
  bfr _b_1365(.a(_w_1679),.q(_w_1680));
  bfr _b_685(.a(_w_999),.q(_w_1000));
  bfr _b_1448(.a(_w_1762),.q(_w_1763));
  spl4L g66_s_0(.a(n66),.q0(n66_0),.q1(n66_1),.q2(n66_2),.q3(n66_3));
  bfr _b_766(.a(_w_1080),.q(_w_1081));
  bfr _b_896(.a(_w_1210),.q(_w_1211));
  bfr _b_1155(.a(_w_1469),.q(_w_1470));
  and_bi g192(.a(n191_0),.b(G31_9),.q(n192));
  bfr _b_563(.a(_w_877),.q(_w_878));
  bfr _b_564(.a(_w_878),.q(_w_879));
  and_bi g175(.a(n174),.b(n173),.q(_w_1729));
  bfr _b_599(.a(_w_913),.q(_w_914));
  bfr _b_1082(.a(_w_1396),.q(n128));
  bfr _b_621(.a(_w_935),.q(_w_936));
  bfr _b_567(.a(_w_881),.q(_w_882));
  bfr _b_590(.a(_w_904),.q(G5_0));
  and_bi g91(.a(G1_4),.b(n89_1),.q(n91));
  bfr _b_568(.a(_w_882),.q(_w_883));
  bfr _b_1000(.a(_w_1314),.q(_w_1315));
  bfr _b_570(.a(_w_884),.q(_w_885));
  bfr _b_988(.a(_w_1302),.q(_w_1303));
  bfr _b_572(.a(_w_886),.q(_w_887));
  bfr _b_984(.a(_w_1298),.q(_w_1299));
  bfr _b_573(.a(_w_887),.q(_w_888));
  bfr _b_1477(.a(_w_1791),.q(_w_1792));
  bfr _b_1385(.a(_w_1699),.q(_w_1700));
  bfr _b_659(.a(_w_973),.q(_w_974));
  and_bi g144(.a(G8_4),.b(G5_4),.q(n144));
  bfr _b_574(.a(_w_888),.q(_w_889));
  bfr _b_575(.a(_w_889),.q(_w_890));
  bfr _b_1116(.a(_w_1430),.q(_w_1431));
  bfr _b_576(.a(_w_890),.q(_w_891));
  and_bi g303(.a(n301),.b(n302),.q(n303));
  bfr _b_709(.a(_w_1023),.q(_w_1024));
  spl2 g254_s_0(.a(n254),.q0(n254_0),.q1(n254_1));
  spl2 g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1));
  bfr _b_577(.a(_w_891),.q(G13_5));
  bfr _b_578(.a(_w_892),.q(_w_893));
  spl2 g311_s_0(.a(n311),.q0(n311_0),.q1(n311_1));
  bfr _b_581(.a(_w_895),.q(_w_896));
  bfr _b_640(.a(_w_954),.q(_w_955));
  bfr _b_886(.a(_w_1200),.q(_w_1201));
  bfr _b_583(.a(_w_897),.q(_w_898));
  bfr _b_651(.a(_w_965),.q(_w_966));
  bfr _b_697(.a(_w_1011),.q(_w_1012));
  bfr _b_584(.a(_w_898),.q(_w_899));
  bfr _b_586(.a(_w_900),.q(_w_901));
  spl3L G10_s_1(.a(G10_2),.q0(G10_3),.q1(G10_4),.q2(_w_1137));
  bfr _b_782(.a(_w_1096),.q(_w_1097));
  bfr _b_1251(.a(_w_1565),.q(_w_1566));
  bfr _b_587(.a(_w_901),.q(_w_902));
  bfr _b_1098(.a(_w_1412),.q(_w_1413));
  bfr _b_591(.a(_w_905),.q(G20_1));
  bfr _b_641(.a(_w_955),.q(_w_956));
  bfr _b_596(.a(_w_910),.q(_w_911));
  bfr _b_597(.a(_w_911),.q(_w_912));
  bfr _b_606(.a(_w_920),.q(_w_921));
  bfr _b_882(.a(_w_1196),.q(_w_1197));
  or_bb g255(.a(G11_6),.b(n254_2),.q(n255));
  bfr _b_598(.a(_w_912),.q(_w_913));
  bfr _b_1142(.a(_w_1456),.q(_w_1457));
  bfr _b_600(.a(_w_914),.q(_w_915));
  bfr _b_904(.a(_w_1218),.q(_w_1219));
  bfr _b_601(.a(_w_915),.q(_w_916));
  bfr _b_602(.a(_w_916),.q(_w_917));
  bfr _b_603(.a(_w_917),.q(G31_14));
  bfr _b_1135(.a(_w_1449),.q(_w_1450));
  bfr _b_700(.a(_w_1014),.q(_w_1015));
  bfr _b_604(.a(_w_918),.q(_w_919));
  bfr _b_610(.a(_w_924),.q(_w_925));
  bfr _b_773(.a(_w_1087),.q(_w_1088));
  bfr _b_611(.a(_w_925),.q(_w_926));
  bfr _b_1258(.a(_w_1572),.q(_w_1573));
  bfr _b_613(.a(_w_927),.q(_w_928));
  bfr _b_614(.a(_w_928),.q(_w_929));
  or_bb g54(.a(n41_3),.b(n53_0),.q(n54));
  bfr _b_965(.a(_w_1279),.q(n309));
  bfr _b_617(.a(_w_931),.q(_w_932));
  bfr _b_618(.a(_w_932),.q(_w_933));
  bfr _b_1037(.a(_w_1351),.q(_w_1352));
  bfr _b_622(.a(_w_936),.q(_w_937));
  bfr _b_796(.a(_w_1110),.q(_w_1111));
  bfr _b_1425(.a(G12),.q(_w_1740));
  bfr _b_623(.a(_w_937),.q(_w_938));
  bfr _b_680(.a(_w_994),.q(_w_995));
  bfr _b_1046(.a(_w_1360),.q(_w_1361));
  bfr _b_624(.a(_w_938),.q(_w_939));
  bfr _b_814(.a(_w_1128),.q(_w_1129));
  bfr _b_626(.a(_w_940),.q(_w_941));
  bfr _b_1509(.a(_w_1823),.q(_w_1824));
  bfr _b_632(.a(_w_946),.q(_w_947));
  bfr _b_875(.a(_w_1189),.q(_w_1190));
  spl2 G9_s_2(.a(G9_5),.q0(G9_6),.q1(G9_7));
  bfr _b_627(.a(_w_941),.q(_w_942));
  and_bb g259(.a(G12_7),.b(n254_5),.q(n259));
  bfr _b_628(.a(_w_942),.q(_w_943));
  bfr _b_747(.a(_w_1061),.q(_w_1062));
  and_bb g153(.a(G27_0),.b(n152_0),.q(n153));
  bfr _b_876(.a(_w_1190),.q(_w_1191));
  bfr _b_629(.a(_w_943),.q(_w_944));
  bfr _b_630(.a(_w_944),.q(_w_945));
  bfr _b_1510(.a(_w_1824),.q(_w_1825));
  bfr _b_633(.a(_w_947),.q(_w_948));
  bfr _b_1538(.a(G8),.q(_w_1853));
  bfr _b_868(.a(_w_1182),.q(G2_5));
  bfr _b_635(.a(_w_949),.q(_w_950));
  bfr _b_636(.a(_w_950),.q(_w_951));
  bfr _b_1286(.a(_w_1600),.q(G1884));
  bfr _b_638(.a(_w_952),.q(_w_953));
  bfr _b_620(.a(_w_934),.q(_w_935));
  bfr _b_1020(.a(_w_1334),.q(_w_1335));
  bfr _b_642(.a(_w_956),.q(_w_957));
  spl2 g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1));
  bfr _b_644(.a(_w_958),.q(_w_959));
  bfr _b_1066(.a(_w_1380),.q(_w_1381));
  bfr _b_828(.a(_w_1142),.q(_w_1143));
  spl2 g234_s_0(.a(n234),.q0(n234_0),.q1(n234_1));
  and_bi g98(.a(n96),.b(n97),.q(n98));
  bfr _b_649(.a(_w_963),.q(_w_964));
  bfr _b_653(.a(_w_967),.q(_w_968));
  bfr _b_654(.a(_w_968),.q(_w_969));
  bfr _b_655(.a(_w_969),.q(_w_970));
  bfr _b_818(.a(_w_1132),.q(_w_1133));
  bfr _b_637(.a(_w_951),.q(_w_952));
  bfr _b_981(.a(_w_1295),.q(_w_1296));
  bfr _b_1368(.a(_w_1682),.q(G7_2));
  bfr _b_658(.a(_w_972),.q(_w_973));
  bfr _b_1044(.a(_w_1358),.q(_w_1359));
  bfr _b_662(.a(_w_976),.q(_w_977));
  bfr _b_663(.a(_w_977),.q(_w_978));
  bfr _b_1446(.a(_w_1760),.q(_w_1761));
  bfr _b_664(.a(_w_978),.q(_w_979));
  bfr _b_686(.a(_w_1000),.q(_w_1001));
  bfr _b_979(.a(_w_1293),.q(_w_1294));
  bfr _b_1225(.a(_w_1539),.q(_w_1540));
  bfr _b_669(.a(_w_983),.q(_w_984));
  bfr _b_1096(.a(_w_1410),.q(_w_1411));
  bfr _b_670(.a(_w_984),.q(G6_5));
  bfr _b_1400(.a(_w_1714),.q(_w_1715));
  bfr _b_891(.a(_w_1205),.q(G4_8));
  bfr _b_671(.a(_w_985),.q(_w_986));
  bfr _b_729(.a(_w_1043),.q(_w_1044));
  bfr _b_673(.a(_w_987),.q(_w_988));
  bfr _b_619(.a(_w_933),.q(_w_934));
  bfr _b_839(.a(_w_1153),.q(_w_1154));
  bfr _b_501(.a(_w_815),.q(_w_816));
  bfr _b_661(.a(_w_975),.q(_w_976));
  bfr _b_676(.a(_w_990),.q(_w_991));
  bfr _b_678(.a(_w_992),.q(_w_993));
  bfr _b_679(.a(_w_993),.q(_w_994));
  bfr _b_1019(.a(_w_1333),.q(G27_2));
  bfr _b_938(.a(_w_1252),.q(_w_1253));
  and_bi g172(.a(n171_0),.b(G31_2),.q(n172));
  and_bb g48(.a(G1_0),.b(n47_0),.q(n48));
  bfr _b_682(.a(_w_996),.q(_w_997));
  bfr _b_683(.a(_w_997),.q(G32_1));
  bfr _b_689(.a(_w_1003),.q(_w_1004));
  bfr _b_690(.a(_w_1004),.q(_w_1005));
  bfr _b_691(.a(_w_1005),.q(_w_1006));
  bfr _b_694(.a(_w_1008),.q(_w_1009));
  bfr _b_698(.a(_w_1012),.q(_w_1013));
  bfr _b_699(.a(_w_1013),.q(_w_1014));
  bfr _b_1436(.a(G20),.q(_w_1751));
  bfr _b_701(.a(_w_1015),.q(_w_1016));
  bfr _b_784(.a(_w_1098),.q(G21_0));
  bfr _b_702(.a(_w_1016),.q(_w_1017));
  bfr _b_1367(.a(_w_1681),.q(_w_1682));
  bfr _b_704(.a(_w_1018),.q(_w_1019));
  bfr _b_1326(.a(_w_1640),.q(_w_1641));
  bfr _b_556(.a(_w_870),.q(_w_871));
  bfr _b_1005(.a(_w_1319),.q(G1904));
  and_bb g230(.a(G16_7),.b(n222_11),.q(n230));
  bfr _b_707(.a(_w_1021),.q(G3_5));
  bfr _b_996(.a(_w_1310),.q(_w_1311));
  bfr _b_708(.a(_w_1022),.q(_w_1023));
  bfr _b_893(.a(_w_1207),.q(_w_1208));
  bfr _b_710(.a(_w_1024),.q(_w_1025));
  bfr _b_711(.a(_w_1025),.q(_w_1026));
  bfr _b_714(.a(_w_1028),.q(_w_1029));
  bfr _b_715(.a(_w_1029),.q(_w_1030));
  bfr _b_919(.a(_w_1233),.q(_w_1234));
  bfr _b_716(.a(_w_1030),.q(_w_1031));
  bfr _b_930(.a(_w_1244),.q(_w_1245));
  bfr _b_717(.a(_w_1031),.q(_w_1032));
  or_bb g148(.a(n146),.b(n147),.q(n148));
  bfr _b_639(.a(_w_953),.q(_w_954));
  bfr _b_720(.a(_w_1034),.q(_w_1035));
  bfr _b_1008(.a(_w_1322),.q(_w_1323));
  bfr _b_723(.a(_w_1037),.q(n98_1));
  bfr _b_724(.a(_w_1038),.q(_w_1039));
  bfr _b_1054(.a(_w_1368),.q(_w_1369));
  and_bb g159(.a(G8_6),.b(n158_0),.q(n159));
  bfr _b_1022(.a(_w_1336),.q(_w_1337));
  bfr _b_725(.a(_w_1039),.q(_w_1040));
  bfr _b_1494(.a(_w_1808),.q(_w_1809));
  bfr _b_1238(.a(_w_1552),.q(_w_1553));
  bfr _b_582(.a(_w_896),.q(_w_897));
  bfr _b_727(.a(_w_1041),.q(_w_1042));
  bfr _b_1390(.a(_w_1704),.q(_w_1705));
  bfr _b_728(.a(_w_1042),.q(_w_1043));
  bfr _b_734(.a(_w_1048),.q(_w_1049));
  bfr _b_884(.a(_w_1198),.q(_w_1199));
  or_bb g189(.a(n188_0),.b(n87_0),.q(n189));
  bfr _b_677(.a(_w_991),.q(_w_992));
  bfr _b_735(.a(_w_1049),.q(_w_1050));
  bfr _b_1483(.a(_w_1797),.q(_w_1798));
  bfr _b_737(.a(_w_1051),.q(_w_1052));
  bfr _b_740(.a(_w_1054),.q(_w_1055));
  bfr _b_1097(.a(_w_1411),.q(_w_1412));
  bfr _b_732(.a(_w_1046),.q(_w_1047));
  bfr _b_783(.a(_w_1097),.q(_w_1098));
  bfr _b_743(.a(_w_1057),.q(_w_1058));
  and_bi g136(.a(n134),.b(n135),.q(n136));
  bfr _b_808(.a(_w_1122),.q(G30_1));
  bfr _b_745(.a(_w_1059),.q(_w_1060));
  bfr _b_746(.a(_w_1060),.q(_w_1061));
  bfr _b_748(.a(_w_1062),.q(G11_5));
  bfr _b_749(.a(_w_1063),.q(_w_1064));
  bfr _b_939(.a(_w_1253),.q(_w_1254));
  spl2 g204_s_0(.a(n204),.q0(n204_0),.q1(n204_1));
  bfr _b_752(.a(_w_1066),.q(_w_1067));
  bfr _b_753(.a(_w_1067),.q(_w_1068));
  bfr _b_779(.a(_w_1093),.q(_w_1094));
  bfr _b_754(.a(_w_1068),.q(_w_1069));
  bfr _b_1009(.a(_w_1323),.q(_w_1324));
  bfr _b_817(.a(_w_1131),.q(_w_1132));
  bfr _b_755(.a(_w_1069),.q(_w_1070));
  bfr _b_756(.a(_w_1070),.q(_w_1071));
  bfr _b_757(.a(_w_1071),.q(_w_1072));
  bfr _b_927(.a(_w_1241),.q(G1907));
  bfr _b_759(.a(_w_1073),.q(_w_1074));
  bfr _b_922(.a(_w_1236),.q(G8_5));
  bfr _b_760(.a(_w_1074),.q(G25_2));
  bfr _b_924(.a(_w_1238),.q(G4_2));
  bfr _b_762(.a(_w_1076),.q(G3_2));
  bfr _b_763(.a(_w_1077),.q(_w_1078));
  and_bi g142(.a(n141),.b(n140),.q(n142));
  bfr _b_764(.a(_w_1078),.q(_w_1079));
  bfr _b_770(.a(_w_1084),.q(_w_1085));
  bfr _b_940(.a(_w_1254),.q(_w_1255));
  bfr _b_781(.a(_w_1095),.q(_w_1096));
  bfr _b_1024(.a(_w_1338),.q(_w_1339));
  bfr _b_1102(.a(_w_1416),.q(_w_1417));
  or_bb g145(.a(n143),.b(n144),.q(n145));
  bfr _b_625(.a(_w_939),.q(G9_5));
  bfr _b_774(.a(_w_1088),.q(_w_1089));
  bfr _b_775(.a(_w_1089),.q(_w_1090));
  bfr _b_852(.a(_w_1166),.q(_w_1167));
  bfr _b_778(.a(_w_1092),.q(_w_1093));
  bfr _b_1430(.a(G17),.q(_w_1745));
  bfr _b_539(.a(_w_853),.q(_w_854));
  bfr _b_780(.a(_w_1094),.q(_w_1095));
  bfr _b_787(.a(_w_1101),.q(n77_2));
  bfr _b_788(.a(_w_1102),.q(G24_2));
  bfr _b_789(.a(_w_1103),.q(_w_1104));
  bfr _b_791(.a(_w_1105),.q(_w_1106));
  bfr _b_771(.a(_w_1085),.q(_w_1086));
  bfr _b_792(.a(_w_1106),.q(_w_1107));
  bfr _b_793(.a(_w_1107),.q(G33_10));
  bfr _b_798(.a(_w_1112),.q(_w_1113));
  bfr _b_799(.a(_w_1113),.q(_w_1114));
  bfr _b_1505(.a(_w_1819),.q(_w_1820));
  spl2 g139_s_0(.a(n139),.q0(n139_0),.q1(n139_1));
  bfr _b_947(.a(_w_1261),.q(_w_1262));
  bfr _b_977(.a(_w_1291),.q(_w_1292));
  bfr _b_801(.a(_w_1115),.q(_w_1116));
  bfr _b_802(.a(_w_1116),.q(_w_1117));
  bfr _b_952(.a(_w_1266),.q(_w_1267));
  bfr _b_803(.a(_w_1117),.q(_w_1118));
  bfr _b_804(.a(_w_1118),.q(_w_1119));
  bfr _b_1089(.a(_w_1403),.q(_w_1404));
  bfr _b_805(.a(_w_1119),.q(_w_1120));
  bfr _b_1027(.a(_w_1341),.q(_w_1342));
  bfr _b_806(.a(_w_1120),.q(_w_1121));
  bfr _b_809(.a(_w_1123),.q(_w_1124));
  bfr _b_1308(.a(_w_1622),.q(_w_1623));
  bfr _b_810(.a(_w_1124),.q(_w_1125));
  bfr _b_812(.a(_w_1126),.q(_w_1127));
  bfr _b_813(.a(_w_1127),.q(_w_1128));
  bfr _b_1511(.a(_w_1825),.q(_w_1826));
  bfr _b_506(.a(_w_820),.q(_w_821));
  bfr _b_816(.a(_w_1130),.q(_w_1131));
  bfr _b_900(.a(_w_1214),.q(_w_1215));
  bfr _b_1095(.a(_w_1409),.q(_w_1410));
  bfr _b_819(.a(_w_1133),.q(_w_1134));
  bfr _b_823(.a(_w_1137),.q(_w_1138));
  bfr _b_824(.a(_w_1138),.q(_w_1139));
  bfr _b_825(.a(_w_1139),.q(_w_1140));
  bfr _b_827(.a(_w_1141),.q(_w_1142));
  bfr _b_953(.a(_w_1267),.q(_w_1268));
  bfr _b_830(.a(_w_1144),.q(_w_1145));
  bfr _b_742(.a(_w_1056),.q(_w_1057));
  bfr _b_935(.a(_w_1249),.q(_w_1250));
  bfr _b_674(.a(_w_988),.q(_w_989));
  bfr _b_834(.a(_w_1148),.q(_w_1149));
  bfr _b_1208(.a(_w_1522),.q(_w_1523));
  spl3L g56_s_0(.a(n56),.q0(n56_0),.q1(n56_1),.q2(_w_1229));
  bfr _b_835(.a(_w_1149),.q(_w_1150));
  bfr _b_836(.a(_w_1150),.q(_w_1151));
  bfr _b_837(.a(_w_1151),.q(_w_1152));
  bfr _b_846(.a(_w_1160),.q(_w_1161));
  bfr _b_968(.a(_w_1282),.q(_w_1283));
  bfr _b_838(.a(_w_1152),.q(_w_1153));
  bfr _b_991(.a(_w_1305),.q(_w_1306));
  bfr _b_840(.a(_w_1154),.q(_w_1155));
  bfr _b_1411(.a(_w_1725),.q(_w_1726));
  bfr _b_843(.a(_w_1157),.q(_w_1158));
  and_bi g181(.a(G14_1),.b(G4_1),.q(n181));
  bfr _b_645(.a(_w_959),.q(_w_960));
  bfr _b_667(.a(_w_981),.q(_w_982));
  bfr _b_847(.a(_w_1161),.q(_w_1162));
  bfr _b_850(.a(_w_1164),.q(_w_1165));
  spl3L G1_s_0(.a(_w_1736),.q0(G1_0),.q1(G1_1),.q2(G1_2));
  bfr _b_851(.a(_w_1165),.q(_w_1166));
  bfr _b_849(.a(_w_1163),.q(_w_1164));
  bfr _b_856(.a(_w_1170),.q(_w_1171));
  spl2 g178_s_1(.a(n178_1),.q0(n178_2),.q1(n178_3));
  bfr _b_1029(.a(_w_1343),.q(_w_1344));
  bfr _b_857(.a(_w_1171),.q(_w_1172));
  bfr _b_858(.a(_w_1172),.q(_w_1173));
  and_bb g132(.a(n102),.b(n131),.q(n132));
  bfr _b_859(.a(_w_1173),.q(_w_1174));
  bfr _b_865(.a(_w_1179),.q(_w_1180));
  bfr _b_866(.a(_w_1180),.q(_w_1181));
  and_bi g293(.a(n171_1),.b(n292),.q(n293));
  and_bi g51(.a(n50_0),.b(n44_0),.q(n51));
  bfr _b_869(.a(_w_1183),.q(_w_1184));
  bfr _b_870(.a(_w_1184),.q(_w_1185));
  bfr _b_1508(.a(_w_1822),.q(_w_1823));
  bfr _b_871(.a(_w_1185),.q(_w_1186));
  bfr _b_1478(.a(_w_1792),.q(_w_1793));
  bfr _b_877(.a(_w_1191),.q(_w_1192));
  bfr _b_719(.a(_w_1033),.q(_w_1034));
  bfr _b_878(.a(_w_1192),.q(_w_1193));
  bfr _b_879(.a(_w_1193),.q(_w_1194));
  bfr _b_883(.a(_w_1197),.q(_w_1198));
  spl3L G7_s_0(.a(_w_1851),.q0(G7_0),.q1(G7_1),.q2(_w_1681));
  bfr _b_885(.a(_w_1199),.q(_w_1200));
  bfr _b_887(.a(_w_1201),.q(_w_1202));
  bfr _b_888(.a(_w_1202),.q(_w_1203));
  bfr _b_1031(.a(_w_1345),.q(_w_1346));
  bfr _b_909(.a(_w_1223),.q(_w_1224));
  bfr _b_889(.a(_w_1203),.q(_w_1204));
  bfr _b_1383(.a(_w_1697),.q(_w_1698));
  spl4L G5_s_1(.a(G5_1),.q0(G5_2),.q1(G5_3),.q2(G5_4),.q3(_w_1432));
  or_bb g87(.a(n85),.b(n86),.q(n87));
  bfr _b_892(.a(_w_1206),.q(_w_1207));
  bfr _b_925(.a(_w_1239),.q(_w_1240));
  bfr _b_1003(.a(_w_1317),.q(n171_1));
  bfr _b_894(.a(_w_1208),.q(_w_1209));
  bfr _b_1469(.a(_w_1783),.q(_w_1784));
  bfr _b_534(.a(_w_848),.q(_w_849));
  bfr _b_705(.a(_w_1019),.q(_w_1020));
  bfr _b_895(.a(_w_1209),.q(_w_1210));
  bfr _b_897(.a(_w_1211),.q(_w_1212));
  bfr _b_901(.a(_w_1215),.q(_w_1216));
  bfr _b_1315(.a(_w_1629),.q(_w_1630));
  spl4L g235_s_1(.a(n235_0),.q0(n235_2),.q1(n235_3),.q2(n235_4),.q3(n235_5));
  bfr _b_902(.a(_w_1216),.q(_w_1217));
  or_bb g81(.a(n79),.b(n80),.q(n81));
  bfr _b_903(.a(_w_1217),.q(_w_1218));
  bfr _b_905(.a(_w_1219),.q(_w_1220));
  bfr _b_1346(.a(_w_1660),.q(_w_1661));
  bfr _b_906(.a(_w_1220),.q(_w_1221));
  spl2 g60_s_0(.a(n60),.q0(n60_0),.q1(n60_1));
  bfr _b_907(.a(_w_1221),.q(_w_1222));
  bfr _b_911(.a(_w_1225),.q(_w_1226));
  or_bi g266(.a(n265),.b(n264),.q(_w_1454));
  bfr _b_913(.a(_w_1227),.q(_w_1228));
  and_bi g117(.a(G4_6),.b(G7_3),.q(n117));
  bfr _b_684(.a(_w_998),.q(_w_999));
  bfr _b_912(.a(_w_1226),.q(_w_1227));
  bfr _b_914(.a(_w_1228),.q(G1_5));
  bfr _b_916(.a(_w_1230),.q(_w_1231));
  bfr _b_920(.a(_w_1234),.q(n56_2));
  and_bi g279(.a(n203_4),.b(n278),.q(n279));
  bfr _b_921(.a(_w_1235),.q(n203_4));
  bfr _b_923(.a(_w_1237),.q(_w_1238));
  bfr _b_1182(.a(_w_1496),.q(_w_1497));
  bfr _b_929(.a(_w_1243),.q(_w_1244));
  bfr _b_1492(.a(_w_1806),.q(_w_1807));
  bfr _b_1392(.a(_w_1706),.q(G1898));
  bfr _b_566(.a(_w_880),.q(_w_881));
  bfr _b_931(.a(_w_1245),.q(_w_1246));
  bfr _b_933(.a(_w_1247),.q(_w_1248));
  bfr _b_848(.a(_w_1162),.q(G10_2));
  and_bb g94(.a(n41_1),.b(n92_1),.q(n94));
  bfr _b_1006(.a(_w_1320),.q(G6_2));
  bfr _b_934(.a(_w_1248),.q(_w_1249));
  bfr _b_941(.a(_w_1255),.q(_w_1256));
  bfr _b_1415(.a(_w_1729),.q(n175));
  bfr _b_942(.a(_w_1256),.q(_w_1257));
  bfr _b_945(.a(_w_1259),.q(_w_1260));
  bfr _b_1382(.a(_w_1696),.q(_w_1697));
  bfr _b_948(.a(_w_1262),.q(_w_1263));
  bfr _b_526(.a(_w_840),.q(_w_841));
  bfr _b_949(.a(_w_1263),.q(_w_1264));
  spl2 g177_s_1(.a(n177_1),.q0(n177_2),.q1(n177_3));
  bfr _b_950(.a(_w_1264),.q(n312));
  bfr _b_973(.a(_w_1287),.q(_w_1288));
  spl2 g136_s_0(.a(n136),.q0(n136_0),.q1(n136_1));
  bfr _b_593(.a(_w_907),.q(_w_908));
  bfr _b_955(.a(_w_1269),.q(_w_1270));
  bfr _b_761(.a(_w_1075),.q(_w_1076));
  bfr _b_975(.a(_w_1289),.q(n300));
  bfr _b_1015(.a(_w_1329),.q(_w_1330));
  bfr _b_956(.a(_w_1270),.q(_w_1271));
  bfr _b_1209(.a(_w_1523),.q(_w_1524));
  bfr _b_960(.a(_w_1274),.q(_w_1275));
  bfr _b_961(.a(_w_1275),.q(_w_1276));
  bfr _b_1353(.a(_w_1667),.q(_w_1668));
  spl2 g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1));
  bfr _b_548(.a(_w_862),.q(_w_863));
  bfr _b_962(.a(_w_1276),.q(_w_1277));
  bfr _b_963(.a(_w_1277),.q(_w_1278));
  bfr _b_964(.a(_w_1278),.q(_w_1279));
  bfr _b_969(.a(_w_1283),.q(_w_1284));
  spl2 g281_s_0(.a(n281),.q0(n281_0),.q1(n281_1));
  bfr _b_910(.a(_w_1224),.q(_w_1225));
  bfr _b_741(.a(_w_1055),.q(_w_1056));
  bfr _b_972(.a(_w_1286),.q(_w_1287));
  bfr _b_1284(.a(_w_1598),.q(_w_1599));
  bfr _b_1252(.a(_w_1566),.q(_w_1567));
  bfr _b_974(.a(_w_1288),.q(_w_1289));
  bfr _b_976(.a(_w_1290),.q(_w_1291));
  bfr _b_980(.a(_w_1294),.q(_w_1295));
  bfr _b_983(.a(_w_1297),.q(_w_1298));
  bfr _b_736(.a(_w_1050),.q(_w_1051));
  bfr _b_987(.a(_w_1301),.q(_w_1302));
  bfr _b_989(.a(_w_1303),.q(_w_1304));
  bfr _b_997(.a(_w_1311),.q(_w_1312));
  and_bi g44(.a(n42),.b(n43),.q(n44));
  bfr _b_998(.a(_w_1312),.q(_w_1313));
  bfr _b_994(.a(_w_1308),.q(_w_1309));
  bfr _b_1001(.a(_w_1315),.q(_w_1316));
  bfr _b_1002(.a(_w_1316),.q(_w_1317));
  bfr _b_1004(.a(_w_1318),.q(G1905));
  bfr _b_1007(.a(_w_1321),.q(_w_1322));
  bfr _b_1010(.a(_w_1324),.q(_w_1325));
  bfr _b_986(.a(_w_1300),.q(_w_1301));
  bfr _b_1011(.a(_w_1325),.q(_w_1326));
  bfr _b_1487(.a(_w_1801),.q(_w_1802));
  bfr _b_1012(.a(_w_1326),.q(_w_1327));
  bfr _b_1013(.a(_w_1327),.q(_w_1328));
  bfr _b_1331(.a(_w_1645),.q(G1885));
  bfr _b_946(.a(_w_1260),.q(_w_1261));
  or_bb g239(.a(G6_6),.b(n235_4),.q(n239));
  bfr _b_1017(.a(_w_1331),.q(_w_1332));
  bfr _b_1021(.a(_w_1335),.q(_w_1336));
  bfr _b_867(.a(_w_1181),.q(_w_1182));
  bfr _b_1023(.a(_w_1337),.q(_w_1338));
  bfr _b_726(.a(_w_1040),.q(_w_1041));
  bfr _b_863(.a(_w_1177),.q(_w_1178));
  bfr _b_579(.a(_w_893),.q(_w_894));
  bfr _b_1025(.a(_w_1339),.q(_w_1340));
  bfr _b_800(.a(_w_1114),.q(_w_1115));
  bfr _b_1026(.a(_w_1340),.q(_w_1341));
  bfr _b_1030(.a(_w_1344),.q(_w_1345));
  and_bb g284(.a(n192_2),.b(n281_1),.q(n284));
  bfr _b_1032(.a(_w_1346),.q(n200));
  bfr _b_1033(.a(_w_1347),.q(_w_1348));
  bfr _b_1034(.a(_w_1348),.q(_w_1349));
  bfr _b_1035(.a(_w_1349),.q(_w_1350));
  bfr _b_1036(.a(_w_1350),.q(_w_1351));
  bfr _b_1285(.a(_w_1599),.q(_w_1600));
  bfr _b_687(.a(_w_1001),.q(_w_1002));
  bfr _b_1038(.a(_w_1352),.q(_w_1353));
  bfr _b_854(.a(_w_1168),.q(_w_1169));
  bfr _b_1041(.a(_w_1355),.q(_w_1356));
  bfr _b_499(.a(_w_813),.q(_w_814));
  bfr _b_822(.a(_w_1136),.q(G28_2));
  bfr _b_608(.a(_w_922),.q(_w_923));
  bfr _b_1050(.a(_w_1364),.q(_w_1365));
  and_bi g139(.a(n137),.b(n138),.q(n139));
  bfr _b_954(.a(_w_1268),.q(_w_1269));
  bfr _b_936(.a(_w_1250),.q(_w_1251));
  bfr _b_1053(.a(_w_1367),.q(_w_1368));
  bfr _b_1296(.a(_w_1610),.q(_w_1611));
  bfr _b_1058(.a(_w_1372),.q(_w_1373));
  bfr _b_1185(.a(_w_1499),.q(_w_1500));
  bfr _b_1059(.a(_w_1373),.q(_w_1374));
  bfr _b_1060(.a(_w_1374),.q(_w_1375));
  bfr _b_1223(.a(_w_1537),.q(_w_1538));
  bfr _b_1062(.a(_w_1376),.q(_w_1377));
  bfr _b_1065(.a(_w_1379),.q(_w_1380));
  bfr _b_978(.a(_w_1292),.q(_w_1293));
  bfr _b_1107(.a(_w_1421),.q(_w_1422));
  bfr _b_529(.a(_w_843),.q(_w_844));
  bfr _b_1068(.a(_w_1382),.q(_w_1383));
  bfr _b_1070(.a(_w_1384),.q(_w_1385));
  bfr _b_1071(.a(_w_1385),.q(G15_5));
  bfr _b_1072(.a(_w_1386),.q(n41_2));
  bfr _b_1447(.a(_w_1761),.q(_w_1762));
  bfr _b_1073(.a(_w_1387),.q(_w_1388));
  bfr _b_1184(.a(_w_1498),.q(_w_1499));
  bfr _b_561(.a(_w_875),.q(_w_876));
  bfr _b_1074(.a(_w_1388),.q(_w_1389));
  bfr _b_1076(.a(_w_1390),.q(_w_1391));
  bfr _b_1438(.a(G21),.q(_w_1752));
  bfr _b_1078(.a(_w_1392),.q(_w_1393));
  bfr _b_881(.a(_w_1195),.q(_w_1196));
  bfr _b_1080(.a(_w_1394),.q(_w_1395));
  bfr _b_1084(.a(_w_1398),.q(_w_1399));
  bfr _b_1088(.a(_w_1402),.q(_w_1403));
  bfr _b_1090(.a(_w_1404),.q(_w_1405));
  bfr _b_1094(.a(_w_1408),.q(_w_1409));
  bfr _b_1099(.a(_w_1413),.q(_w_1414));
  bfr _b_1101(.a(_w_1415),.q(_w_1416));
  bfr _b_1104(.a(_w_1418),.q(_w_1419));
  spl2 g316_s_0(.a(n316),.q0(n316_0),.q1(n316_1));
  bfr _b_1106(.a(_w_1420),.q(_w_1421));
  bfr _b_1108(.a(_w_1422),.q(_w_1423));
endmodule
