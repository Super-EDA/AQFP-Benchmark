module comparator (
    bn0,
    bn1,
    bn2,
    bn3,
    bn4,
    bn5,
    bn6,
    bn7,
    bn8,
    bn9,
    bn10,
    bn11,
    bn12,
    bn13,
    bn14,
    bn15,
    bn16,
    bn17,
    bn18,
    bn19,
    bn20,
    bn21,
    bn22,
    bn23,
    bn24,
    bn25,
    bn26,
    bn27,
    bn28,
    bn29,
    bn30,
    bn31,
    rn0,
    rn1,
    rn2,
    rn3,
    rn4,
    rn5,
    rn6,
    rn7,
    rn8,
    rn9,
    rn10,
    rn11,
    rn12,
    rn13,
    rn14,
    rn15,
    rn16,
    rn17,
    rn18,
    rn19,
    rn20,
    rn21,
    rn22,
    rn23,
    rn24,
    rn25,
    rn26,
    rn27,
    rn28,
    rn29,
    rn30,
    rn31,
    s
);
  wire nn_0_;
  wire nn_1_;
  wire nn_2_;
  wire nn_3_;
  wire nn_4_;
  wire nn_5_;
  wire nn_6_;
  wire nn_7_;
  wire nn_8_;
  wire nn_9_;
  wire nn_10_;
  wire nn_11_;
  wire nn_12_;
  wire nn_13_;
  wire nn_14_;
  wire nn_15_;
  wire nn_16_;
  wire nn_17_;
  wire nn_18_;
  wire nn_19_;
  wire nn_20_;
  wire nn_21_;
  wire nn_22_;
  wire nn_23_;
  wire nn_24_;
  wire nn_25_;
  wire nn_26_;
  wire nn_27_;
  wire nn_28_;
  wire nn_29_;
  wire nn_30_;
  wire nn_31_;
  wire nn_32_;
  wire nn_33_;
  wire nn_34_;
  wire nn_35_;
  wire nn_36_;
  wire nn_37_;
  wire nn_38_;
  wire nn_39_;
  wire nn_40_;
  wire nn_41_;
  wire nn_42_;
  wire nn_43_;
  wire nn_44_;
  wire nn_45_;
  wire nn_46_;
  wire nn_47_;
  wire nn_48_;
  wire nn_49_;
  wire nn_50_;
  wire nn_51_;
  wire nn_52_;
  wire nn_53_;
  wire nn_54_;
  wire nn_55_;
  wire nn_56_;
  wire nn_57_;
  wire nn_58_;
  wire nn_59_;
  wire nn_60_;
  wire nn_61_;
  wire nn_62_;
  wire nn_63_;
  wire nn_64_;
  wire nn_65_;
  wire nn_66_;
  wire nn_67_;
  wire nn_68_;
  wire nn_69_;
  wire nn_70_;
  wire nn_71_;
  wire nn_72_;
  wire nn_73_;
  wire nn_74_;
  wire nn_75_;
  wire nn_76_;
  wire nn_77_;
  wire nn_78_;
  wire nn_79_;
  wire nn_80_;
  wire nn_81_;
  wire nn_82_;
  wire nn_83_;
  wire nn_84_;
  wire nn_85_;
  wire nn_86_;
  wire nn_87_;
  wire nn_88_;
  wire nn_89_;
  wire nn_90_;
  wire nn_91_;
  wire nn_92_;
  wire nn_93_;
  wire nn_94_;
  wire nn_95_;
  wire nn_96_;
  wire nn_97_;
  wire nn_98_;
  wire nn_99_;
  wire nn_100_;
  wire nn_101_;
  wire nn_102_;
  wire nn_103_;
  wire nn_104_;
  wire nn_105_;
  wire nn_106_;
  wire nn_107_;
  wire nn_108_;
  wire nn_109_;
  wire nn_110_;
  wire nn_111_;
  wire nn_112_;
  wire nn_113_;
  wire nn_114_;
  wire nn_115_;
  wire nn_116_;
  wire nn_117_;
  wire nn_118_;
  wire nn_119_;
  wire nn_120_;
  wire nn_121_;
  wire nn_122_;
  wire nn_123_;
  wire nn_124_;
  wire nn_125_;
  wire nn_126_;
  wire nn_127_;
  wire nn_128_;
  wire nn_129_;
  wire nn_130_;
  wire nn_131_;
  wire nn_132_;
  wire nn_133_;
  wire nn_134_;
  wire nn_135_;
  wire nn_136_;
  wire nn_137_;
  wire nn_138_;
  wire nn_139_;
  wire nn_140_;
  wire nn_141_;
  wire nn_142_;
  wire nn_143_;
  wire nn_144_;
  wire nn_145_;
  wire nn_146_;
  wire nn_147_;
  wire nn_148_;
  wire nn_149_;
  wire nn_150_;
  wire nn_151_;
  wire nn_152_;
  wire nn_153_;
  wire nn_154_;
  wire nn_155_;
  wire nn_156_;
  wire nn_157_;
  wire nn_158_;
  wire nn_159_;
  wire nn_160_;
  wire nn_161_;
  wire nn_162_;
  wire nn_163_;
  wire nn_164_;
  wire nn_165_;
  wire nn_166_;
  wire nn_167_;
  wire nn_168_;
  wire nn_169_;
  wire nn_170_;
  wire nn_171_;
  wire nn_172_;
  wire nn_173_;
  wire nn_174_;
  wire nn_175_;
  wire nn_176_;
  wire nn_177_;
  wire nn_178_;
  wire nn_179_;
  wire nn_180_;
  wire nn_181_;
  wire nn_182_;
  wire nn_183_;
  wire nn_184_;
  wire nn_185_;
  wire nn_186_;
  wire nn_187_;
  wire nn_188_;
  wire nn_189_;
  wire nn_190_;
  wire nn_191_;
  wire nn_192_;
  wire nn_193_;
  wire nn_194_;
  wire nn_195_;
  wire nn_196_;
  wire nn_197_;
  wire nn_198_;
  wire nn_199_;
  wire nn_200_;
  wire nn_201_;
  wire nn_202_;
  wire nn_203_;
  wire nn_204_;
  wire nn_205_;
  wire nn_206_;
  wire nn_207_;
  wire nn_208_;
  wire nn_209_;
  wire nn_210_;
  wire nn_211_;
  wire nn_212_;
  wire nn_213_;
  wire nn_214_;
  wire nn_215_;
  wire nn_216_;
  wire nn_217_;
  wire nn_218_;
  wire nn_219_;
  wire nn_220_;
  wire nn_221_;
  wire nn_222_;
  wire nn_223_;
  wire nn_224_;
  wire nn_225_;
  wire nn_226_;
  wire nn_227_;
  wire nn_228_;
  wire nn_229_;
  wire nn_230_;
  wire nn_231_;
  wire nn_232_;
  wire nn_233_;
  wire nn_234_;
  wire nn_235_;
  wire nn_236_;
  wire nn_237_;
  wire nn_238_;
  wire nn_239_;
  wire nn_240_;
  wire nn_241_;
  wire nn_242_;
  wire nn_243_;
  wire nn_244_;
  wire nn_245_;
  wire nn_246_;
  wire nn_247_;
  wire nn_248_;
  wire nn_249_;
  wire nn_250_;
  wire nn_251_;
  wire nn_252_;
  wire nn_253_;
  wire nn_254_;
  wire nn_255_;
  wire nn_256_;
  wire nn_257_;
  wire nn_258_;
  wire nn_259_;
  wire nn_260_;
  wire nn_261_;
  wire nn_262_;
  wire nn_263_;
  wire nn_264_;
  wire nn_265_;
  wire nn_266_;
  wire nn_267_;
  wire nn_268_;
  wire nn_269_;
  wire nn_270_;
  wire nn_271_;
  wire nn_272_;
  wire nn_273_;
  wire nn_274_;
  wire nn_275_;
  wire nn_276_;
  wire nn_277_;
  wire nn_278_;
  wire nn_279_;
  wire nn_280_;
  wire nn_281_;
  wire nn_282_;
  wire nn_283_;
  wire nn_284_;
  wire nn_285_;
  wire nn_286_;
  wire nn_287_;
  wire nn_288_;
  wire nn_289_;
  wire nn_290_;
  wire nn_291_;
  wire nn_292_;
  wire nn_293_;
  wire nn_294_;
  wire nn_295_;
  wire nn_296_;
  wire nn_297_;
  wire nn_298_;
  wire nn_299_;
  wire nn_300_;
  wire nn_301_;
  wire nn_302_;
  wire nn_303_;
  wire nn_304_;
  wire nn_305_;
  wire nn_306_;
  wire nn_307_;
  wire nn_308_;
  wire nn_309_;
  wire nn_310_;
  wire nn_311_;
  wire nn_312_;
  wire nn_313_;
  wire nn_314_;
  wire nn_315_;
  wire nn_316_;
  wire nn_317_;
  wire nn_318_;
  wire nn_319_;
  wire nn_320_;
  wire nn_321_;
  wire nn_322_;
  wire nn_323_;
  wire nn_324_;
  wire nn_325_;
  wire nn_326_;
  wire nn_327_;
  wire nn_328_;
  wire nn_329_;
  wire nn_330_;
  wire nn_331_;
  wire nn_332_;
  wire nn_333_;
  wire nn_334_;
  wire nn_335_;
  wire nn_336_;
  wire nn_337_;
  wire nn_338_;
  wire nn_339_;
  wire nn_340_;
  wire nn_341_;
  wire nn_342_;
  wire nn_343_;
  wire nn_344_;
  wire nn_345_;
  wire nn_346_;
  wire nn_347_;
  wire nn_348_;
  wire nn_349_;
  wire nn_350_;
  wire nn_351_;
  wire nn_352_;
  wire nn_353_;
  wire nn_354_;
  wire nn_355_;
  wire nn_356_;
  wire nn_357_;
  wire nn_358_;
  wire nn_359_;
  wire nn_360_;
  wire nn_361_;
  wire nn_362_;
  wire nn_363_;
  wire nn_364_;
  wire nn_365_;
  wire nn_366_;
  wire nn_367_;
  wire nn_368_;
  wire nn_369_;
  wire nn_370_;
  wire nn_371_;
  wire nn_372_;
  wire nn_373_;
  wire nn_374_;
  wire nn_375_;
  wire nn_376_;
  wire nn_377_;
  wire nn_378_;
  wire nn_379_;
  wire nn_380_;
  wire nn_381_;
  wire nn_382_;
  wire nn_383_;
  wire nn_384_;
  wire nn_385_;
  wire nn_386_;
  wire nn_387_;
  wire nn_388_;
  wire nn_389_;
  wire nn_390_;
  wire nn_391_;
  wire nn_392_;
  wire nn_393_;
  wire nn_394_;
  wire nn_395_;
  wire nn_396_;
  wire nn_397_;
  wire nn_398_;
  wire nn_399_;
  wire nn_400_;
  wire nn_401_;
  wire nn_402_;
  wire nn_403_;
  wire nn_404_;
  wire nn_405_;
  wire nn_406_;
  wire nn_407_;
  wire nn_408_;
  wire nn_409_;
  wire nn_410_;
  wire nn_411_;
  wire nn_412_;
  wire nn_413_;
  wire nn_414_;
  wire nn_415_;
  wire nn_416_;
  wire nn_417_;
  wire nn_418_;
  wire nn_419_;
  wire nn_420_;
  wire nn_421_;
  wire nn_422_;
  wire nn_423_;
  wire nn_424_;
  wire nn_425_;
  wire nn_426_;
  wire nn_427_;
  wire nn_428_;
  wire nn_429_;
  wire nn_430_;
  wire nn_431_;
  wire nn_432_;
  wire nn_433_;
  wire nn_434_;
  wire nn_435_;
  wire nn_436_;
  wire nn_437_;
  wire nn_438_;
  wire nn_439_;
  wire nn_440_;
  wire nn_441_;
  wire nn_442_;
  wire nn_443_;
  wire nn_444_;
  wire nn_445_;
  wire nn_446_;
  wire nn_447_;
  wire nn_448_;
  wire nn_449_;
  wire nn_450_;
  wire nn_451_;
  wire nn_452_;
  wire nn_453_;
  wire nn_454_;
  wire nn_455_;
  wire nn_456_;
  wire nn_457_;
  wire nn_458_;
  wire nn_459_;
  wire nn_460_;
  wire nn_461_;
  wire nn_462_;
  wire nn_463_;
  wire nn_464_;
  wire nn_465_;
  wire nn_466_;
  wire nn_467_;
  wire nn_468_;
  wire nn_469_;
  wire nn_470_;
  wire nn_471_;
  wire nn_472_;
  wire nn_473_;
  wire nn_474_;
  wire nn_475_;
  wire nn_476_;
  wire nn_477_;
  wire nn_478_;
  wire nn_479_;
  wire nn_480_;
  wire nn_481_;
  wire nn_482_;
  wire nn_483_;
  wire nn_484_;
  wire nn_485_;
  wire nn_486_;
  wire nn_487_;
  wire nn_488_;
  wire nn_489_;
  wire nn_490_;
  wire nn_491_;
  wire nn_492_;
  wire nn_493_;
  wire nn_494_;
  wire nn_495_;
  wire nn_496_;
  wire nn_497_;
  wire nn_498_;
  wire nn_499_;
  wire nn_500_;
  wire nn_501_;
  wire nn_502_;
  wire nn_503_;
  wire nn_504_;
  wire nn_505_;
  wire nn_506_;
  wire nn_507_;
  wire nn_508_;
  wire nn_509_;
  wire nn_510_;
  wire nn_511_;
  wire nn_512_;
  wire nn_513_;
  wire nn_514_;
  wire nn_515_;
  wire nn_516_;
  wire nn_517_;
  wire nn_518_;
  wire nn_519_;
  wire nn_520_;
  wire nn_521_;
  wire nn_522_;
  wire nn_523_;
  wire nn_524_;
  wire nn_525_;
  wire nn_526_;
  wire nn_527_;
  wire nn_528_;
  wire nn_529_;
  wire nn_530_;
  wire nn_531_;
  wire nn_532_;
  wire nn_533_;
  wire nn_534_;
  wire nn_535_;
  wire nn_536_;
  wire nn_537_;
  wire nn_538_;
  wire nn_539_;
  wire nn_540_;
  input bn0;
  input bn1;
  input bn2;
  input bn3;
  input bn4;
  input bn5;
  input bn6;
  input bn7;
  input bn8;
  input bn9;
  input bn10;
  input bn11;
  input bn12;
  input bn13;
  input bn14;
  input bn15;
  input bn16;
  input bn17;
  input bn18;
  input bn19;
  input bn20;
  input bn21;
  input bn22;
  input bn23;
  input bn24;
  input bn25;
  input bn26;
  input bn27;
  input bn28;
  input bn29;
  input bn30;
  input bn31;
  input rn0;
  input rn1;
  input rn2;
  input rn3;
  input rn4;
  input rn5;
  input rn6;
  input rn7;
  input rn8;
  input rn9;
  input rn10;
  input rn11;
  input rn12;
  input rn13;
  input rn14;
  input rn15;
  input rn16;
  input rn17;
  input rn18;
  input rn19;
  input rn20;
  input rn21;
  input rn22;
  input rn23;
  input rn24;
  input rn25;
  input rn26;
  input rn27;
  input rn28;
  input rn29;
  input rn30;
  input rn31;
  output s;

  and_bi gg_0_ (
      .a(nn_63_),
      .b(nn_387_),
      .q(nn_534_)
  );

  or_bi gg_1_ (
      .a(nn_495_),
      .b(nn_466_),
      .q(nn_385_)
  );

  or_bb gg_2_ (
      .a(nn_302_),
      .b(nn_366_),
      .q(nn_535_)
  );

  bfr gg_3_ (
      .a(nn_248_),
      .q(nn_507_)
  );

  bfr gg_4_ (
      .a(nn_0_),
      .q(nn_166_)
  );

  maj_bib gg_5_ (
      .a(nn_178_),
      .b(nn_449_),
      .c(nn_298_),
      .q(nn_440_)
  );

  or_bb gg_6_ (
      .a(nn_25_),
      .b(nn_99_),
      .q(nn_290_)
  );

  and_bi gg_7_ (
      .a(nn_226_),
      .b(nn_297_),
      .q(nn_343_)
  );

  spl2 gg_8_ (
      .a (nn_82_),
      .q0(nn_513_),
      .q1(nn_487_)
  );

  bfr gg_9_ (
      .a(nn_141_),
      .q(nn_344_)
  );

  spl2 gg_10_ (
      .a (bn16),
      .q0(nn_199_),
      .q1(nn_177_)
  );

  bfr gg_11_ (
      .a(nn_127_),
      .q(nn_226_)
  );

  bfr gg_12_ (
      .a(nn_445_),
      .q(nn_503_)
  );

  bfr gg_13_ (
      .a(nn_313_),
      .q(nn_278_)
  );

  bfr gg_14_ (
      .a(nn_439_),
      .q(nn_336_)
  );

  spl3L gg_15_ (
      .a (bn17),
      .q0(nn_101_),
      .q1(nn_27_),
      .q2(nn_88_)
  );

  bfr gg_16_ (
      .a(nn_102_),
      .q(nn_24_)
  );

  spl2 gg_17_ (
      .a (rn28),
      .q0(nn_104_),
      .q1(nn_6_)
  );

  bfr gg_18_ (
      .a(nn_150_),
      .q(nn_415_)
  );

  bfr gg_19_ (
      .a(nn_214_),
      .q(nn_529_)
  );

  bfr gg_20_ (
      .a(nn_507_),
      .q(nn_337_)
  );

  bfr gg_21_ (
      .a(nn_186_),
      .q(nn_523_)
  );

  and_bi gg_22_ (
      .a(nn_325_),
      .b(nn_484_),
      .q(nn_11_)
  );

  and_bi gg_23_ (
      .a(nn_263_),
      .b(nn_199_),
      .q(nn_12_)
  );

  or_bb gg_24_ (
      .a(nn_79_),
      .b(nn_52_),
      .q(nn_13_)
  );

  and_bb gg_25_ (
      .a(nn_209_),
      .b(nn_360_),
      .q(nn_81_)
  );

  spl2 gg_26_ (
      .a (bn6),
      .q0(nn_434_),
      .q1(nn_393_)
  );

  bfr gg_27_ (
      .a(nn_32_),
      .q(nn_346_)
  );

  bfr gg_28_ (
      .a(nn_503_),
      .q(nn_477_)
  );

  bfr gg_29_ (
      .a(nn_100_),
      .q(nn_69_)
  );

  bfr gg_30_ (
      .a(nn_101_),
      .q(nn_200_)
  );

  spl2 gg_31_ (
      .a (bn18),
      .q0(nn_84_),
      .q1(nn_60_)
  );

  bfr gg_32_ (
      .a(nn_104_),
      .q(nn_137_)
  );

  bfr gg_33_ (
      .a(nn_489_),
      .q(nn_469_)
  );

  bfr gg_34_ (
      .a(nn_274_),
      .q(nn_219_)
  );

  and_bi gg_35_ (
      .a(nn_16_),
      .b(nn_352_),
      .q(nn_481_)
  );

  spl3L gg_36_ (
      .a (rn23),
      .q0(nn_54_),
      .q1(nn_424_),
      .q2(nn_486_)
  );

  spl2 gg_37_ (
      .a (rn21),
      .q0(nn_121_),
      .q1(nn_83_)
  );

  or_bi gg_38_ (
      .a(nn_91_),
      .b(nn_184_),
      .q(nn_505_)
  );

  and_bi gg_39_ (
      .a(nn_369_),
      .b(nn_15_),
      .q(nn_20_)
  );

  and_bi gg_40_ (
      .a(nn_359_),
      .b(nn_512_),
      .q(nn_506_)
  );

  or_bi gg_41_ (
      .a(nn_332_),
      .b(nn_121_),
      .q(nn_96_)
  );

  bfr gg_42_ (
      .a(nn_8_),
      .q(nn_496_)
  );

  bfr gg_43_ (
      .a(nn_65_),
      .q(nn_75_)
  );

  spl2 gg_44_ (
      .a (rn2),
      .q0(nn_203_),
      .q1(nn_184_)
  );

  bfr gg_45_ (
      .a(nn_67_),
      .q(nn_9_)
  );

  spl2 gg_46_ (
      .a (rn18),
      .q0(nn_301_),
      .q1(nn_270_)
  );

  bfr gg_47_ (
      .a(nn_210_),
      .q(nn_349_)
  );

  bfr gg_48_ (
      .a(nn_532_),
      .q(nn_245_)
  );

  and_bi gg_49_ (
      .a(nn_174_),
      .b(nn_433_),
      .q(nn_517_)
  );

  and_ib gg_50_ (
      .a(nn_292_),
      .b(nn_478_),
      .q(nn_156_)
  );

  or_bb gg_51_ (
      .a(nn_136_),
      .b(nn_278_),
      .q(nn_41_)
  );

  spl2 gg_52_ (
      .a (nn_156_),
      .q0(nn_23_),
      .q1(nn_8_)
  );

  bfr gg_53_ (
      .a(nn_140_),
      .q(nn_416_)
  );

  bfr gg_54_ (
      .a(nn_9_),
      .q(nn_476_)
  );

  or_bb gg_55_ (
      .a(nn_86_),
      .b(nn_164_),
      .q(nn_134_)
  );

  or_bb gg_56_ (
      .a(nn_461_),
      .b(nn_416_),
      .q(nn_49_)
  );

  spl2 gg_57_ (
      .a (nn_222_),
      .q0(nn_532_),
      .q1(nn_209_)
  );

  bfr gg_58_ (
      .a(nn_307_),
      .q(nn_428_)
  );

  bfr gg_59_ (
      .a(nn_526_),
      .q(nn_158_)
  );

  or_bb gg_60_ (
      .a(nn_142_),
      .b(nn_223_),
      .q(nn_57_)
  );

  or_bi gg_61_ (
      .a(nn_434_),
      .b(nn_154_),
      .q(nn_58_)
  );

  and_bi gg_62_ (
      .a(nn_6_),
      .b(nn_197_),
      .q(nn_59_)
  );

  spl2 gg_63_ (
      .a (bn2),
      .q0(nn_131_),
      .q1(nn_91_)
  );

  bfr gg_64_ (
      .a(nn_155_),
      .q(nn_217_)
  );

  bfr gg_65_ (
      .a(nn_523_),
      .q(nn_240_)
  );

  or_bb gg_66_ (
      .a(nn_148_),
      .b(nn_42_),
      .q(nn_71_)
  );

  or_bi gg_67_ (
      .a(nn_483_),
      .b(nn_176_),
      .q(nn_72_)
  );

  and_bi gg_68_ (
      .a(nn_356_),
      .b(nn_5_),
      .q(nn_524_)
  );

  and_bi gg_69_ (
      .a(nn_259_),
      .b(nn_88_),
      .q(nn_526_)
  );

  spl2 gg_70_ (
      .a (bn22),
      .q0(nn_175_),
      .q1(nn_143_)
  );

  bfr gg_71_ (
      .a(nn_54_),
      .q(nn_255_)
  );

  bfr gg_72_ (
      .a(nn_213_),
      .q(nn_38_)
  );

  bfr gg_73_ (
      .a(nn_240_),
      .q(nn_225_)
  );

  bfr gg_74_ (
      .a(nn_21_),
      .q(nn_46_)
  );

  or_bb gg_75_ (
      .a(nn_415_),
      .b(nn_260_),
      .q(nn_384_)
  );

  and_bi gg_76_ (
      .a(nn_486_),
      .b(nn_94_),
      .q(nn_80_)
  );

  bfr gg_77_ (
      .a(nn_504_),
      .q(nn_55_)
  );

  bfr gg_78_ (
      .a(nn_193_),
      .q(nn_56_)
  );

  bfr gg_79_ (
      .a(nn_39_),
      .q(nn_10_)
  );

  or_bb gg_80_ (
      .a(nn_217_),
      .b(nn_171_),
      .q(nn_413_)
  );

  and_bi gg_81_ (
      .a(nn_237_),
      .b(nn_426_),
      .q(nn_19_)
  );

  and_ib gg_82_ (
      .a(nn_464_),
      .b(nn_4_),
      .q(nn_412_)
  );

  spl2 gg_83_ (
      .a (nn_354_),
      .q0(nn_297_),
      .q1(nn_261_)
  );

  bfr gg_84_ (
      .a(nn_314_),
      .q(nn_66_)
  );

  bfr gg_85_ (
      .a(nn_482_),
      .q(nn_473_)
  );

  spl2 gg_86_ (
      .a (bn3),
      .q0(nn_31_),
      .q1(nn_17_)
  );

  bfr gg_87_ (
      .a(nn_221_),
      .q(nn_76_)
  );

  or_bb gg_88_ (
      .a(nn_162_),
      .b(nn_180_),
      .q(nn_92_)
  );

  or_bb gg_89_ (
      .a(nn_321_),
      .b(nn_284_),
      .q(nn_127_)
  );

  maj_bbi gg_90_ (
      .a(nn_392_),
      .b(nn_235_),
      .c(nn_26_),
      .q(nn_454_)
  );

  bfr gg_91_ (
      .a(nn_385_),
      .q(nn_401_)
  );

  or_bb gg_92_ (
      .a(nn_282_),
      .b(nn_130_),
      .q(nn_363_)
  );

  bfr gg_93_ (
      .a(nn_200_),
      .q(nn_64_)
  );

  bfr gg_94_ (
      .a(nn_137_),
      .q(nn_26_)
  );

  spl2 gg_95_ (
      .a (bn30),
      .q0(nn_305_),
      .q1(nn_272_)
  );

  bfr gg_96_ (
      .a(nn_66_),
      .q(nn_528_)
  );

  maj_bib gg_97_ (
      .a(nn_153_),
      .b(nn_195_),
      .c(nn_491_),
      .q(nn_459_)
  );

  or_bb gg_98_ (
      .a(nn_331_),
      .b(nn_454_),
      .q(nn_441_)
  );

  spl2 gg_99_ (
      .a (rn14),
      .q0(nn_244_),
      .q1(nn_207_)
  );

  spl2 gg_100_ (
      .a (rn16),
      .q0(nn_263_),
      .q1(nn_238_)
  );

  spl2 gg_101_ (
      .a (rn20),
      .q0(nn_210_),
      .q1(nn_521_)
  );

  spl2 gg_102_ (
      .a (rn10),
      .q0(nn_35_),
      .q1(nn_15_)
  );

  bfr gg_103_ (
      .a(nn_76_),
      .q(nn_97_)
  );

  or_bi gg_104_ (
      .a(nn_30_),
      .b(nn_427_),
      .q(nn_40_)
  );

  maj_bib gg_105_ (
      .a(nn_513_),
      .b(nn_435_),
      .c(nn_514_),
      .q(nn_442_)
  );

  bfr gg_106_ (
      .a(nn_299_),
      .q(nn_311_)
  );

  or_bi gg_107_ (
      .a(nn_31_),
      .b(nn_151_),
      .q(nn_48_)
  );

  and_bi gg_108_ (
      .a(nn_68_),
      .b(nn_456_),
      .q(nn_439_)
  );

  or_bb gg_109_ (
      .a(nn_190_),
      .b(nn_218_),
      .q(nn_1_)
  );

  bfr gg_110_ (
      .a(nn_349_),
      .q(nn_7_)
  );

  bfr gg_111_ (
      .a(nn_38_),
      .q(nn_95_)
  );

  or_bb gg_112_ (
      .a(nn_538_),
      .b(nn_215_),
      .q(nn_135_)
  );

  and_bb gg_113_ (
      .a(nn_23_),
      .b(nn_338_),
      .q(nn_136_)
  );

  bfr gg_114_ (
      .a(nn_119_),
      .q(nn_105_)
  );

  bfr gg_115_ (
      .a(nn_134_),
      .q(nn_341_)
  );

  bfr gg_116_ (
      .a(nn_46_),
      .q(nn_274_)
  );

  and_bi gg_117_ (
      .a(nn_2_),
      .b(nn_243_),
      .q(nn_140_)
  );

  and_bi gg_118_ (
      .a(nn_181_),
      .b(nn_175_),
      .q(nn_73_)
  );

  spl2 gg_119_ (
      .a (nn_161_),
      .q0(nn_294_),
      .q1(nn_260_)
  );

  bfr gg_120_ (
      .a(nn_185_),
      .q(nn_111_)
  );

  bfr gg_121_ (
      .a(nn_55_),
      .q(nn_112_)
  );

  bfr gg_122_ (
      .a(nn_95_),
      .q(nn_281_)
  );

  bfr gg_123_ (
      .a(nn_56_),
      .q(nn_113_)
  );

  bfr gg_124_ (
      .a(nn_335_),
      .q(nn_114_)
  );

  bfr gg_125_ (
      .a(nn_10_),
      .q(nn_115_)
  );

  and_bi gg_126_ (
      .a(nn_230_),
      .b(nn_281_),
      .q(nn_142_)
  );

  or_bb gg_127_ (
      .a(nn_529_),
      .b(nn_146_),
      .q(nn_474_)
  );

  or_bb gg_128_ (
      .a(nn_188_),
      .b(nn_98_),
      .q(nn_77_)
  );

  spl2 gg_129_ (
      .a (nn_135_),
      .q0(nn_322_),
      .q1(nn_292_)
  );

  spl2 gg_130_ (
      .a (nn_96_),
      .q0(nn_381_),
      .q1(nn_360_)
  );

  spl2 gg_131_ (
      .a (bn21),
      .q0(nn_332_),
      .q1(nn_304_)
  );

  spl3L gg_132_ (
      .a (bn31),
      .q0(nn_249_),
      .q1(nn_205_),
      .q2(nn_268_)
  );

  bfr gg_133_ (
      .a(nn_105_),
      .q(nn_159_)
  );

  bfr gg_134_ (
      .a(nn_257_),
      .q(nn_276_)
  );

  bfr gg_135_ (
      .a(nn_47_),
      .q(nn_125_)
  );

  and_bb gg_136_ (
      .a(nn_241_),
      .b(nn_97_),
      .q(nn_148_)
  );

  maj_bib gg_137_ (
      .a(nn_367_),
      .b(nn_388_),
      .c(nn_24_),
      .q(nn_525_)
  );

  spl2 gg_138_ (
      .a (rn6),
      .q0(nn_154_),
      .q1(nn_132_)
  );

  bfr gg_139_ (
      .a(nn_255_),
      .q(nn_455_)
  );

  bfr gg_140_ (
      .a(nn_111_),
      .q(nn_110_)
  );

  bfr gg_141_ (
      .a(nn_232_),
      .q(nn_98_)
  );

  bfr gg_142_ (
      .a(nn_113_),
      .q(nn_538_)
  );

  spl2 gg_143_ (
      .a (nn_12_),
      .q0(nn_3_),
      .q1(nn_519_)
  );

  bfr gg_144_ (
      .a(nn_118_),
      .q(nn_138_)
  );

  and_bi gg_145_ (
      .a(nn_244_),
      .b(nn_368_),
      .q(nn_161_)
  );

  bfr gg_146_ (
      .a(nn_246_),
      .q(nn_371_)
  );

  and_bi gg_147_ (
      .a(nn_144_),
      .b(nn_208_),
      .q(nn_171_)
  );

  or_bb gg_148_ (
      .a(nn_147_),
      .b(nn_276_),
      .q(nn_307_)
  );

  or_ib gg_149_ (
      .a(nn_337_),
      .b(nn_258_),
      .q(nn_173_)
  );

  maj_bib gg_150_ (
      .a(nn_381_),
      .b(nn_145_),
      .c(nn_7_),
      .q(nn_216_)
  );

  spl2 gg_151_ (
      .a (bn24),
      .q0(nn_236_),
      .q1(nn_198_)
  );

  bfr gg_152_ (
      .a(nn_249_),
      .q(nn_374_)
  );

  bfr gg_153_ (
      .a(nn_138_),
      .q(nn_478_)
  );

  or_bb gg_154_ (
      .a(nn_252_),
      .b(nn_266_),
      .q(nn_139_)
  );

  or_bb gg_155_ (
      .a(nn_407_),
      .b(nn_329_),
      .q(nn_334_)
  );

  and_bi gg_156_ (
      .a(nn_272_),
      .b(nn_432_),
      .q(nn_180_)
  );

  or_bi gg_157_ (
      .a(nn_124_),
      .b(nn_521_),
      .q(nn_222_)
  );

  spl3L gg_158_ (
      .a (bn13),
      .q0(nn_233_),
      .q1(nn_174_),
      .q2(nn_285_)
  );

  spl2 gg_159_ (
      .a (rn7),
      .q0(nn_456_),
      .q1(nn_427_)
  );

  spl3L gg_160_ (
      .a (rn27),
      .q0(nn_286_),
      .q1(nn_295_),
      .q2(nn_358_)
  );

  spl2 gg_161_ (
      .a (bn20),
      .q0(nn_287_),
      .q1(nn_124_)
  );

  and_bi gg_162_ (
      .a(nn_421_),
      .b(nn_87_),
      .q(nn_187_)
  );

  and_bi gg_163_ (
      .a(nn_465_),
      .b(nn_198_),
      .q(nn_82_)
  );

  spl2 gg_164_ (
      .a (bn1),
      .q0(nn_144_),
      .q1(nn_123_)
  );

  spl2 gg_165_ (
      .a (rn22),
      .q0(nn_181_),
      .q1(nn_152_)
  );

  spl3L gg_166_ (
      .a (bn19),
      .q0(nn_299_),
      .q1(nn_485_),
      .q2(nn_512_)
  );

  spl2 gg_167_ (
      .a (rn24),
      .q0(nn_494_),
      .q1(nn_465_)
  );

  bfr gg_168_ (
      .a(nn_341_),
      .q(nn_160_)
  );

  and_bi gg_169_ (
      .a(nn_269_),
      .b(nn_22_),
      .q(nn_126_)
  );

  and_bi gg_170_ (
      .a(nn_304_),
      .b(nn_83_),
      .q(nn_193_)
  );

  bfr gg_171_ (
      .a(nn_285_),
      .q(nn_418_)
  );

  bfr gg_172_ (
      .a(nn_286_),
      .q(nn_317_)
  );

  spl2 gg_173_ (
      .a (rn5),
      .q0(nn_520_),
      .q1(nn_493_)
  );

  bfr gg_174_ (
      .a(nn_287_),
      .q(nn_399_)
  );

  bfr gg_175_ (
      .a(nn_112_),
      .q(nn_167_)
  );

  bfr gg_176_ (
      .a(nn_80_),
      .q(nn_99_)
  );

  bfr gg_177_ (
      .a(nn_253_),
      .q(nn_407_)
  );

  bfr gg_178_ (
      .a(nn_114_),
      .q(nn_168_)
  );

  and_bi gg_179_ (
      .a(nn_189_),
      .b(nn_159_),
      .q(nn_314_)
  );

  or_bb gg_180_ (
      .a(nn_409_),
      .b(nn_291_),
      .q(nn_194_)
  );

  spl2 gg_181_ (
      .a (nn_453_),
      .q0(nn_206_),
      .q1(nn_182_)
  );

  spl2 gg_182_ (
      .a (bn10),
      .q0(nn_396_),
      .q1(nn_369_)
  );

  spl3L gg_183_ (
      .a (bn23),
      .q0(nn_310_),
      .q1(nn_70_),
      .q2(nn_94_)
  );

  bfr gg_184_ (
      .a(nn_311_),
      .q(nn_14_)
  );

  bfr gg_185_ (
      .a(nn_390_),
      .q(nn_410_)
  );

  bfr gg_186_ (
      .a(nn_125_),
      .q(nn_179_)
  );

  bfr gg_187_ (
      .a(nn_212_),
      .q(nn_522_)
  );

  bfr gg_188_ (
      .a(nn_438_),
      .q(nn_0_)
  );

  or_ib gg_189_ (
      .a(nn_280_),
      .b(nn_300_),
      .q(nn_204_)
  );

  spl2 gg_190_ (
      .a (nn_518_),
      .q0(nn_480_),
      .q1(nn_450_)
  );

  spl3L gg_191_ (
      .a (rn31),
      .q0(nn_389_),
      .q1(nn_357_),
      .q2(nn_246_)
  );

  spl3L gg_192_ (
      .a (bn9),
      .q0(nn_316_),
      .q1(nn_356_),
      .q2(nn_422_)
  );

  and_bi gg_193_ (
      .a(nn_467_),
      .b(nn_394_),
      .q(nn_117_)
  );

  or_bb gg_194_ (
      .a(nn_290_),
      .b(nn_44_),
      .q(nn_215_)
  );

  bfr gg_195_ (
      .a(nn_522_),
      .q(nn_283_)
  );

  bfr gg_196_ (
      .a(nn_251_),
      .q(nn_429_)
  );

  and_bi gg_197_ (
      .a(nn_425_),
      .b(nn_36_),
      .q(nn_150_)
  );

  spl2 gg_198_ (
      .a (nn_126_),
      .q0(nn_490_),
      .q1(nn_461_)
  );

  bfr gg_199_ (
      .a(nn_418_),
      .q(nn_195_)
  );

  bfr gg_200_ (
      .a(nn_412_),
      .q(nn_191_)
  );

  or_bb gg_201_ (
      .a(nn_320_),
      .b(nn_344_),
      .q(nn_230_)
  );

  and_bi gg_202_ (
      .a(bn0),
      .b(rn0),
      .q(nn_155_)
  );

  and_bi gg_203_ (
      .a(nn_35_),
      .b(nn_396_),
      .q(nn_231_)
  );

  or_ib gg_204_ (
      .a(nn_308_),
      .b(nn_319_),
      .q(nn_232_)
  );

  spl2 gg_205_ (
      .a (bn14),
      .q0(nn_368_),
      .q1(nn_330_)
  );

  bfr gg_206_ (
      .a(nn_441_),
      .q(nn_201_)
  );

  bfr gg_207_ (
      .a(nn_139_),
      .q(nn_202_)
  );

  bfr gg_208_ (
      .a(nn_527_),
      .q(nn_250_)
  );

  or_bb gg_209_ (
      .a(nn_327_),
      .b(nn_157_),
      .q(nn_241_)
  );

  and_bi gg_210_ (
      .a(nn_205_),
      .b(nn_357_),
      .q(nn_162_)
  );

  spl2 gg_211_ (
      .a (bn26),
      .q0(nn_22_),
      .q1(nn_2_)
  );

  spl3L gg_212_ (
      .a (bn25),
      .q0(nn_466_),
      .q1(nn_394_),
      .q2(nn_348_)
  );

  bfr gg_213_ (
      .a(nn_403_),
      .q(nn_211_)
  );

  bfr gg_214_ (
      .a(nn_191_),
      .q(nn_50_)
  );

  bfr gg_215_ (
      .a(nn_315_),
      .q(nn_157_)
  );

  and_bi gg_216_ (
      .a(nn_463_),
      .b(nn_233_),
      .q(nn_172_)
  );

  spl2 gg_217_ (
      .a (bn28),
      .q0(nn_339_),
      .q1(nn_197_)
  );

  spl3L gg_218_ (
      .a (rn17),
      .q0(nn_259_),
      .q1(nn_234_),
      .q2(nn_340_)
  );

  bfr gg_219_ (
      .a(nn_201_),
      .q(nn_470_)
  );

  bfr gg_220_ (
      .a(nn_160_),
      .q(nn_220_)
  );

  or_bb gg_221_ (
      .a(nn_487_),
      .b(nn_165_),
      .q(nn_335_)
  );

  or_bb gg_222_ (
      .a(nn_328_),
      .b(nn_342_),
      .q(nn_32_)
  );

  maj_bib gg_223_ (
      .a(nn_3_),
      .b(nn_64_),
      .c(nn_293_),
      .q(nn_373_)
  );

  bfr gg_224_ (
      .a(nn_167_),
      .q(nn_227_)
  );

  bfr gg_225_ (
      .a(nn_168_),
      .q(nn_228_)
  );

  bfr gg_226_ (
      .a(nn_169_),
      .q(nn_229_)
  );

  or_bb gg_227_ (
      .a(nn_334_),
      .b(nn_353_),
      .q(nn_257_)
  );

  or_bb gg_228_ (
      .a(nn_261_),
      .b(nn_408_),
      .q(nn_258_)
  );

  spl2 gg_229_ (
      .a (nn_501_),
      .q0(nn_397_),
      .q1(nn_370_)
  );

  bfr gg_230_ (
      .a(nn_339_),
      .q(nn_457_)
  );

  bfr gg_231_ (
      .a(nn_340_),
      .q(nn_458_)
  );

  spl2 gg_232_ (
      .a (bn4),
      .q0(nn_510_),
      .q1(nn_483_)
  );

  spl2 gg_233_ (
      .a (rn4),
      .q0(nn_196_),
      .q1(nn_176_)
  );

  bfr gg_234_ (
      .a(nn_374_),
      .q(nn_242_)
  );

  bfr gg_235_ (
      .a(nn_179_),
      .q(nn_239_)
  );

  bfr gg_236_ (
      .a(nn_309_),
      .q(nn_44_)
  );

  bfr gg_237_ (
      .a(nn_115_),
      .q(nn_169_)
  );

  and_bi gg_238_ (
      .a(nn_510_),
      .b(nn_196_),
      .q(nn_266_)
  );

  and_bi gg_239_ (
      .a(nn_511_),
      .b(nn_361_),
      .q(nn_267_)
  );

  or_bb gg_240_ (
      .a(nn_343_),
      .b(nn_53_),
      .q(nn_119_)
  );

  bfr gg_241_ (
      .a(nn_348_),
      .q(nn_498_)
  );

  spl3L gg_242_ (
      .a (rn19),
      .q0(nn_380_),
      .q1(nn_296_),
      .q2(nn_359_)
  );

  bfr gg_243_ (
      .a(nn_437_),
      .q(nn_67_)
  );

  bfr gg_244_ (
      .a(nn_229_),
      .q(nn_163_)
  );

  bfr gg_245_ (
      .a(nn_457_),
      .q(nn_235_)
  );

  bfr gg_246_ (
      .a(nn_458_),
      .q(nn_293_)
  );

  spl3L gg_247_ (
      .a (bn11),
      .q0(nn_479_),
      .q1(nn_426_),
      .q2(nn_390_)
  );

  spl2 gg_248_ (
      .a (bn29),
      .q0(nn_303_),
      .q1(nn_271_)
  );

  and_bb gg_249_ (
      .a(nn_326_),
      .b(nn_528_),
      .q(s)
  );

  or_bb gg_250_ (
      .a(nn_477_),
      .b(nn_378_),
      .q(nn_39_)
  );

  bfr gg_251_ (
      .a(nn_317_),
      .q(nn_323_)
  );

  bfr gg_252_ (
      .a(nn_380_),
      .q(nn_375_)
  );

  bfr gg_253_ (
      .a(nn_399_),
      .q(nn_145_)
  );

  bfr gg_254_ (
      .a(nn_106_),
      .q(nn_185_)
  );

  bfr gg_255_ (
      .a(nn_275_),
      .q(nn_256_)
  );

  bfr gg_256_ (
      .a(nn_172_),
      .q(nn_282_)
  );

  or_bb gg_257_ (
      .a(nn_372_),
      .b(nn_383_),
      .q(nn_315_)
  );

  and_bi gg_258_ (
      .a(nn_479_),
      .b(nn_262_),
      .q(nn_214_)
  );

  and_ib gg_259_ (
      .a(nn_74_),
      .b(nn_471_),
      .q(nn_291_)
  );

  bfr gg_260_ (
      .a(nn_488_),
      .q(nn_37_)
  );

  bfr gg_261_ (
      .a(nn_410_),
      .q(nn_449_)
  );

  bfr gg_262_ (
      .a(nn_202_),
      .q(nn_264_)
  );

  bfr gg_263_ (
      .a(nn_250_),
      .q(nn_265_)
  );

  and_bi gg_264_ (
      .a(nn_60_),
      .b(nn_270_),
      .q(nn_300_)
  );

  or_bb gg_265_ (
      .a(nn_90_),
      .b(nn_109_),
      .q(nn_79_)
  );

  and_bi gg_266_ (
      .a(nn_395_),
      .b(nn_303_),
      .q(nn_254_)
  );

  spl3L gg_267_ (
      .a (rn11),
      .q0(nn_262_),
      .q1(nn_237_),
      .q2(nn_419_)
  );

  bfr gg_268_ (
      .a(nn_211_),
      .q(nn_273_)
  );

  or_bb gg_269_ (
      .a(nn_384_),
      .b(nn_345_),
      .q(nn_78_)
  );

  and_bb gg_270_ (
      .a(nn_225_),
      .b(nn_405_),
      .q(nn_248_)
  );

  or_bb gg_271_ (
      .a(nn_386_),
      .b(nn_406_),
      .q(nn_309_)
  );

  spl2 gg_272_ (
      .a (nn_379_),
      .q0(nn_133_),
      .q1(nn_90_)
  );

  bfr gg_273_ (
      .a(nn_264_),
      .q(nn_42_)
  );

  bfr gg_274_ (
      .a(nn_194_),
      .q(nn_338_)
  );

  bfr gg_275_ (
      .a(nn_220_),
      .q(nn_279_)
  );

  bfr gg_276_ (
      .a(nn_265_),
      .q(nn_530_)
  );

  maj_bib gg_277_ (
      .a(nn_62_),
      .b(nn_129_),
      .c(nn_455_),
      .q(nn_120_)
  );

  bfr gg_278_ (
      .a(nn_371_),
      .q(nn_423_)
  );

  bfr gg_279_ (
      .a(nn_227_),
      .q(nn_288_)
  );

  bfr gg_280_ (
      .a(nn_228_),
      .q(nn_289_)
  );

  bfr gg_281_ (
      .a(nn_149_),
      .q(nn_164_)
  );

  and_bb gg_282_ (
      .a(nn_420_),
      .b(nn_414_),
      .q(nn_320_)
  );

  and_bi gg_283_ (
      .a(nn_177_),
      .b(nn_238_),
      .q(nn_319_)
  );

  spl2 gg_284_ (
      .a (nn_1_),
      .q0(nn_74_),
      .q1(nn_33_)
  );

  spl3L gg_285_ (
      .a (rn25),
      .q0(nn_495_),
      .q1(nn_467_),
      .q2(nn_443_)
  );

  bfr gg_286_ (
      .a(nn_310_),
      .q(nn_533_)
  );

  bfr gg_287_ (
      .a(nn_239_),
      .q(nn_402_)
  );

  bfr gg_288_ (
      .a(nn_279_),
      .q(nn_223_)
  );

  bfr gg_289_ (
      .a(nn_192_),
      .q(nn_508_)
  );

  or_ib gg_290_ (
      .a(nn_50_),
      .b(nn_430_),
      .q(nn_326_)
  );

  and_bb gg_291_ (
      .a(nn_413_),
      .b(nn_431_),
      .q(nn_327_)
  );

  and_bi gg_292_ (
      .a(nn_85_),
      .b(nn_493_),
      .q(nn_252_)
  );

  and_bi gg_293_ (
      .a(nn_61_),
      .b(nn_422_),
      .q(nn_253_)
  );

  bfr gg_294_ (
      .a(nn_316_),
      .q(nn_539_)
  );

  bfr gg_295_ (
      .a(nn_499_),
      .q(nn_306_)
  );

  bfr gg_296_ (
      .a(nn_289_),
      .q(nn_408_)
  );

  bfr gg_297_ (
      .a(nn_373_),
      .q(nn_312_)
  );

  bfr gg_298_ (
      .a(nn_402_),
      .q(nn_536_)
  );

  and_bi gg_299_ (
      .a(nn_295_),
      .b(nn_34_),
      .q(nn_342_)
  );

  and_bb gg_300_ (
      .a(nn_245_),
      .b(nn_216_),
      .q(nn_118_)
  );

  bfr gg_301_ (
      .a(nn_256_),
      .q(nn_318_)
  );

  or_bb gg_302_ (
      .a(nn_451_),
      .b(nn_336_),
      .q(nn_353_)
  );

  or_bb gg_303_ (
      .a(nn_452_),
      .b(nn_51_),
      .q(nn_213_)
  );

  or_bb gg_304_ (
      .a(nn_182_),
      .b(nn_470_),
      .q(nn_354_)
  );

  and_ib gg_305_ (
      .a(nn_397_),
      .b(nn_347_),
      .q(nn_321_)
  );

  bfr gg_306_ (
      .a(nn_443_),
      .q(nn_502_)
  );

  spl2 gg_307_ (
      .a (rn3),
      .q0(nn_151_),
      .q1(nn_128_)
  );

  bfr gg_308_ (
      .a(nn_312_),
      .q(nn_471_)
  );

  bfr gg_309_ (
      .a(nn_404_),
      .q(nn_345_)
  );

  or_bi gg_310_ (
      .a(nn_296_),
      .b(nn_485_),
      .q(nn_280_)
  );

  or_bb gg_311_ (
      .a(nn_460_),
      .b(nn_110_),
      .q(nn_365_)
  );

  bfr gg_312_ (
      .a(nn_498_),
      .q(nn_435_)
  );

  spl2 gg_313_ (
      .a (bn5),
      .q0(nn_122_),
      .q1(nn_85_)
  );

  bfr gg_314_ (
      .a(nn_273_),
      .q(nn_333_)
  );

  bfr gg_315_ (
      .a(nn_318_),
      .q(nn_409_)
  );

  bfr gg_316_ (
      .a(nn_117_),
      .q(nn_165_)
  );

  maj_bib gg_317_ (
      .a(nn_480_),
      .b(nn_14_),
      .c(nn_324_),
      .q(nn_275_)
  );

  spl3L gg_318_ (
      .a (rn15),
      .q0(nn_488_),
      .q1(nn_352_),
      .q2(nn_425_)
  );

  spl2 gg_319_ (
      .a (rn12),
      .q0(nn_421_),
      .q1(nn_387_)
  );

  bfr gg_320_ (
      .a(nn_447_),
      .q(nn_224_)
  );

  spl2 gg_321_ (
      .a (nn_173_),
      .q0(nn_492_),
      .q1(nn_464_)
  );

  spl2 gg_322_ (
      .a (nn_187_),
      .q0(nn_153_),
      .q1(nn_130_)
  );

  or_bb gg_323_ (
      .a(nn_322_),
      .b(nn_531_),
      .q(nn_21_)
  );

  bfr gg_324_ (
      .a(nn_375_),
      .q(nn_324_)
  );

  bfr gg_325_ (
      .a(nn_288_),
      .q(nn_350_)
  );

  and_ib gg_326_ (
      .a(nn_116_),
      .b(nn_537_),
      .q(nn_378_)
  );

  bfr gg_327_ (
      .a(nn_459_),
      .q(nn_351_)
  );

  and_bi gg_328_ (
      .a(nn_131_),
      .b(nn_203_),
      .q(nn_383_)
  );

  or_bi gg_329_ (
      .a(nn_234_),
      .b(nn_27_),
      .q(nn_308_)
  );

  spl2 gg_330_ (
      .a (nn_247_),
      .q0(nn_170_),
      .q1(nn_147_)
  );

  spl2 gg_331_ (
      .a (nn_267_),
      .q0(nn_367_),
      .q1(nn_329_)
  );

  bfr gg_332_ (
      .a(nn_37_),
      .q(nn_382_)
  );

  bfr gg_333_ (
      .a(nn_508_),
      .q(nn_251_)
  );

  or_bi gg_334_ (
      .a(nn_122_),
      .b(nn_520_),
      .q(nn_47_)
  );

  or_bb gg_335_ (
      .a(nn_474_),
      .b(nn_469_),
      .q(nn_247_)
  );

  or_bb gg_336_ (
      .a(nn_363_),
      .b(nn_224_),
      .q(nn_149_)
  );

  and_bi gg_337_ (
      .a(nn_389_),
      .b(nn_268_),
      .q(nn_398_)
  );

  bfr gg_338_ (
      .a(nn_29_),
      .q(nn_45_)
  );

  bfr gg_339_ (
      .a(nn_350_),
      .q(nn_107_)
  );

  bfr gg_340_ (
      .a(nn_351_),
      .q(nn_537_)
  );

  bfr gg_341_ (
      .a(nn_306_),
      .q(nn_18_)
  );

  or_bb gg_342_ (
      .a(nn_481_),
      .b(nn_500_),
      .q(nn_404_)
  );

  and_bi gg_343_ (
      .a(nn_283_),
      .b(nn_370_),
      .q(nn_405_)
  );

  and_bi gg_344_ (
      .a(nn_143_),
      .b(nn_152_),
      .q(nn_406_)
  );

  spl2 gg_345_ (
      .a (nn_231_),
      .q0(nn_178_),
      .q1(nn_146_)
  );

  bfr gg_346_ (
      .a(nn_77_),
      .q(nn_43_)
  );

  bfr gg_347_ (
      .a(nn_355_),
      .q(nn_376_)
  );

  bfr gg_348_ (
      .a(nn_81_),
      .q(nn_377_)
  );

  and_bi gg_349_ (
      .a(nn_93_),
      .b(nn_358_),
      .q(nn_328_)
  );

  spl3L gg_350_ (
      .a (bn15),
      .q0(nn_36_),
      .q1(nn_16_),
      .q2(nn_28_)
  );

  bfr gg_351_ (
      .a(nn_497_),
      .q(nn_100_)
  );

  bfr gg_352_ (
      .a(nn_120_),
      .q(nn_192_)
  );

  or_bb gg_353_ (
      .a(nn_476_),
      .b(nn_509_),
      .q(nn_420_)
  );

  bfr gg_354_ (
      .a(nn_533_),
      .q(nn_129_)
  );

  or_bb gg_355_ (
      .a(nn_515_),
      .b(nn_107_),
      .q(nn_430_)
  );

  and_bb gg_356_ (
      .a(nn_505_),
      .b(nn_516_),
      .q(nn_431_)
  );

  or_bb gg_357_ (
      .a(nn_277_),
      .b(nn_450_),
      .q(nn_190_)
  );

  or_bi gg_358_ (
      .a(nn_492_),
      .b(nn_475_),
      .q(nn_189_)
  );

  bfr gg_359_ (
      .a(nn_539_),
      .q(nn_388_)
  );

  spl3L gg_360_ (
      .a (rn9),
      .q0(nn_61_),
      .q1(nn_5_),
      .q2(nn_540_)
  );

  bfr gg_361_ (
      .a(nn_419_),
      .q(nn_103_)
  );

  bfr gg_362_ (
      .a(nn_448_),
      .q(nn_106_)
  );

  bfr gg_363_ (
      .a(nn_333_),
      .q(nn_400_)
  );

  bfr gg_364_ (
      .a(nn_473_),
      .q(nn_212_)
  );

  maj_bib gg_365_ (
      .a(nn_133_),
      .b(nn_242_),
      .c(nn_423_),
      .q(nn_448_)
  );

  bfr gg_366_ (
      .a(nn_440_),
      .q(nn_411_)
  );

  or_bb gg_367_ (
      .a(nn_517_),
      .b(nn_534_),
      .q(nn_447_)
  );

  bfr gg_368_ (
      .a(nn_204_),
      .q(nn_218_)
  );

  spl2 gg_369_ (
      .a (rn8),
      .q0(nn_511_),
      .q1(nn_484_)
  );

  bfr gg_370_ (
      .a(nn_506_),
      .q(nn_277_)
  );

  or_bb gg_371_ (
      .a(nn_158_),
      .b(nn_519_),
      .q(nn_188_)
  );

  and_bi gg_372_ (
      .a(nn_17_),
      .b(nn_128_),
      .q(nn_372_)
  );

  or_bb gg_373_ (
      .a(nn_524_),
      .b(nn_11_),
      .q(nn_451_)
  );

  and_ib gg_374_ (
      .a(nn_170_),
      .b(nn_108_),
      .q(nn_452_)
  );

  or_bb gg_375_ (
      .a(nn_530_),
      .b(nn_13_),
      .q(nn_453_)
  );

  spl2 gg_376_ (
      .a (nn_78_),
      .q0(nn_116_),
      .q1(nn_86_)
  );

  bfr gg_377_ (
      .a(nn_502_),
      .q(nn_514_)
  );

  spl2 gg_378_ (
      .a (rn26),
      .q0(nn_269_),
      .q1(nn_243_)
  );

  bfr gg_379_ (
      .a(nn_535_),
      .q(nn_438_)
  );

  and_bi gg_380_ (
      .a(nn_393_),
      .b(nn_132_),
      .q(nn_499_)
  );

  maj_bib gg_381_ (
      .a(nn_294_),
      .b(nn_75_),
      .c(nn_382_),
      .q(nn_364_)
  );

  and_bi gg_382_ (
      .a(nn_462_),
      .b(nn_305_),
      .q(nn_379_)
  );

  and_bi gg_383_ (
      .a(nn_166_),
      .b(nn_206_),
      .q(nn_460_)
  );

  bfr gg_384_ (
      .a(nn_417_),
      .q(nn_4_)
  );

  spl2 gg_385_ (
      .a (nn_73_),
      .q0(nn_62_),
      .q1(nn_25_)
  );

  spl3L gg_386_ (
      .a (bn27),
      .q0(nn_497_),
      .q1(nn_34_),
      .q2(nn_93_)
  );

  bfr gg_387_ (
      .a(nn_540_),
      .q(nn_102_)
  );

  bfr gg_388_ (
      .a(nn_442_),
      .q(nn_436_)
  );

  bfr gg_389_ (
      .a(nn_18_),
      .q(nn_437_)
  );

  and_bi gg_390_ (
      .a(nn_70_),
      .b(nn_424_),
      .q(nn_386_)
  );

  spl2 gg_391_ (
      .a (bn12),
      .q0(nn_87_),
      .q1(nn_63_)
  );

  bfr gg_392_ (
      .a(nn_376_),
      .q(nn_444_)
  );

  bfr gg_393_ (
      .a(nn_364_),
      .q(nn_445_)
  );

  bfr gg_394_ (
      .a(nn_377_),
      .q(nn_446_)
  );

  or_bi gg_395_ (
      .a(nn_494_),
      .b(nn_236_),
      .q(nn_482_)
  );

  bfr gg_396_ (
      .a(nn_89_),
      .q(nn_331_)
  );

  spl3L gg_397_ (
      .a (rn13),
      .q0(nn_463_),
      .q1(nn_433_),
      .q2(nn_29_)
  );

  spl2 gg_398_ (
      .a (rn1),
      .q0(nn_208_),
      .q1(nn_183_)
  );

  bfr gg_399_ (
      .a(nn_436_),
      .q(nn_347_)
  );

  spl2 gg_400_ (
      .a (bn7),
      .q0(nn_68_),
      .q1(nn_30_)
  );

  spl2 gg_401_ (
      .a (rn30),
      .q0(nn_462_),
      .q1(nn_432_)
  );

  bfr gg_402_ (
      .a(nn_398_),
      .q(nn_109_)
  );

  bfr gg_403_ (
      .a(nn_444_),
      .q(nn_284_)
  );

  bfr gg_404_ (
      .a(nn_446_),
      .q(nn_531_)
  );

  or_bb gg_405_ (
      .a(nn_19_),
      .b(nn_20_),
      .q(nn_489_)
  );

  bfr gg_406_ (
      .a(nn_45_),
      .q(nn_491_)
  );

  bfr gg_407_ (
      .a(nn_400_),
      .q(nn_468_)
  );

  bfr gg_408_ (
      .a(nn_525_),
      .q(nn_391_)
  );

  bfr gg_409_ (
      .a(nn_401_),
      .q(nn_186_)
  );

  and_bi gg_410_ (
      .a(nn_330_),
      .b(nn_207_),
      .q(nn_500_)
  );

  or_bb gg_411_ (
      .a(nn_346_),
      .b(nn_49_),
      .q(nn_501_)
  );

  bfr gg_412_ (
      .a(nn_92_),
      .q(nn_52_)
  );

  bfr gg_413_ (
      .a(nn_411_),
      .q(nn_472_)
  );

  or_bi gg_414_ (
      .a(nn_41_),
      .b(nn_219_),
      .q(nn_475_)
  );

  bfr gg_415_ (
      .a(nn_28_),
      .q(nn_65_)
  );

  bfr gg_416_ (
      .a(nn_468_),
      .q(nn_414_)
  );

  bfr gg_417_ (
      .a(nn_391_),
      .q(nn_108_)
  );

  spl2 gg_418_ (
      .a (bn8),
      .q0(nn_361_),
      .q1(nn_325_)
  );

  bfr gg_419_ (
      .a(nn_428_),
      .q(nn_141_)
  );

  and_bb gg_420_ (
      .a(nn_536_),
      .b(nn_71_),
      .q(nn_509_)
  );

  and_bb gg_421_ (
      .a(nn_48_),
      .b(nn_72_),
      .q(nn_221_)
  );

  maj_bib gg_422_ (
      .a(nn_490_),
      .b(nn_69_),
      .c(nn_323_),
      .q(nn_355_)
  );

  spl2 gg_423_ (
      .a (nn_254_),
      .q0(nn_392_),
      .q1(nn_366_)
  );

  spl2 gg_424_ (
      .a (rn29),
      .q0(nn_395_),
      .q1(nn_362_)
  );

  bfr gg_425_ (
      .a(nn_472_),
      .q(nn_51_)
  );

  bfr gg_426_ (
      .a(nn_429_),
      .q(nn_313_)
  );

  and_bi gg_427_ (
      .a(nn_57_),
      .b(nn_163_),
      .q(nn_515_)
  );

  or_bi gg_428_ (
      .a(nn_123_),
      .b(nn_183_),
      .q(nn_516_)
  );

  and_bb gg_429_ (
      .a(nn_40_),
      .b(nn_58_),
      .q(nn_403_)
  );

  or_bb gg_430_ (
      .a(nn_33_),
      .b(nn_43_),
      .q(nn_504_)
  );

  and_bi gg_431_ (
      .a(nn_301_),
      .b(nn_84_),
      .q(nn_518_)
  );

  and_bi gg_432_ (
      .a(nn_271_),
      .b(nn_362_),
      .q(nn_527_)
  );

  bfr gg_433_ (
      .a(nn_496_),
      .q(nn_417_)
  );

  spl2 gg_434_ (
      .a (nn_59_),
      .q0(nn_89_),
      .q1(nn_302_)
  );

  bfr gg_435_ (
      .a(nn_103_),
      .q(nn_298_)
  );

  bfr gg_436_ (
      .a(nn_365_),
      .q(nn_53_)
  );

endmodule
