module full_adder (
    a_0,
    a_1,
    a_2,
    a_3,
    a_4,
    a_5,
    a_6,
    a_7,
    b_0,
    b_1,
    b_2,
    b_3,
    b_4,
    b_5,
    b_6,
    b_7,
    cin,
    s_0,
    s_1,
    s_2,
    s_3,
    s_4,
    s_5,
    s_6,
    s_7,
    cout
);
  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;
  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  input cin;
  output s_0;
  output s_1;
  output s_2;
  output s_3;
  output s_4;
  output s_5;
  output s_6;
  output s_7;
  output cout;
  wire _w_447;
  wire _w_446;
  wire _w_445;
  wire _w_444;
  wire _w_441;
  wire _w_440;
  wire _w_439;
  wire _w_438;
  wire _w_435;
  wire _w_433;
  wire _w_431;
  wire _w_425;
  wire _w_424;
  wire _w_421;
  wire _w_419;
  wire _w_416;
  wire _w_412;
  wire _w_411;
  wire _w_409;
  wire _w_408;
  wire _w_401;
  wire _w_399;
  wire _w_398;
  wire _w_395;
  wire _w_393;
  wire _w_392;
  wire _w_390;
  wire _w_394;
  wire _w_388;
  wire _w_386;
  wire _w_385;
  wire _w_384;
  wire _w_383;
  wire _w_375;
  wire _w_372;
  wire _w_371;
  wire _w_370;
  wire _w_402;
  wire _w_368;
  wire _w_400;
  wire _w_367;
  wire _w_366;
  wire _w_389;
  wire _w_363;
  wire _w_361;
  wire _w_360;
  wire _w_358;
  wire _w_355;
  wire _w_354;
  wire _w_348;
  wire _w_429;
  wire _w_347;
  wire _w_346;
  wire _w_345;
  wire _w_343;
  wire _w_342;
  wire _w_341;
  wire _w_340;
  wire _w_338;
  wire _w_337;
  wire _w_417;
  wire _w_335;
  wire _w_334;
  wire _w_329;
  wire _w_350;
  wire _w_327;
  wire _w_427;
  wire _w_423;
  wire _w_326;
  wire _w_325;
  wire _w_324;
  wire _w_323;
  wire _w_322;
  wire _w_320;
  wire _w_318;
  wire _w_317;
  wire _w_316;
  wire _w_314;
  wire _w_313;
  wire _w_405;
  wire _w_311;
  wire _w_365;
  wire _w_310;
  wire _w_307;
  wire _w_304;
  wire _w_303;
  wire _w_426;
  wire _w_302;
  wire _w_300;
  wire _w_362;
  wire _w_298;
  wire _w_297;
  wire _w_296;
  wire _w_406;
  wire _w_294;
  wire _w_293;
  wire _w_292;
  wire _w_321;
  wire _w_287;
  wire _w_286;
  wire _w_413;
  wire _w_285;
  wire _w_283;
  wire _w_280;
  wire _w_277;
  wire _w_276;
  wire _w_275;
  wire _w_274;
  wire _w_272;
  wire _w_271;
  wire _w_269;
  wire _w_268;
  wire _w_266;
  wire _w_264;
  wire _w_261;
  wire _w_260;
  wire _w_379;
  wire _w_258;
  wire _w_257;
  wire _w_259;
  wire n24_2;
  wire _w_436;
  wire n25_5;
  wire _w_336;
  wire n24_6;
  wire _w_332;
  wire _w_253;
  wire n52_2;
  wire n28_4;
  wire n74_1;
  wire _w_418;
  wire n42_2;
  wire n42_1;
  wire n56;
  wire _w_403;
  wire a_1__2;
  wire n42_0;
  wire _w_279;
  wire n43_2;
  wire _w_443;
  wire n43_0;
  wire _w_377;
  wire n46_2;
  wire _w_265;
  wire n21;
  wire _w_437;
  wire _w_282;
  wire n46_0;
  wire n23_4;
  wire a_0__0;
  wire _w_284;
  wire n53_0;
  wire n53;
  wire n74_0;
  wire n28_0;
  wire _w_263;
  wire n49_1;
  wire _w_380;
  wire n84_1;
  wire n78;
  wire n36;
  wire n39_3;
  wire n84_0;
  wire n86;
  wire b_4__4;
  wire n85;
  wire _w_404;
  wire a_5__0;
  wire _w_319;
  wire n79;
  wire _w_378;
  wire n42_3;
  wire n26;
  wire n75;
  wire _w_369;
  wire n22;
  wire n74;
  wire b_6__4;
  wire _w_434;
  wire n25_0;
  wire n70;
  wire n20_3;
  wire n66;
  wire _w_374;
  wire n21_1;
  wire n64;
  wire n63;
  wire n61;
  wire _w_306;
  wire b_1__3;
  wire n58;
  wire n40;
  wire n47;
  wire n46;
  wire n82;
  wire b_7__1;
  wire _w_428;
  wire n43;
  wire _w_301;
  wire n42;
  wire _w_414;
  wire _w_262;
  wire a_4__2;
  wire a_2__0;
  wire n52_0;
  wire b_6__1;
  wire n46_1;
  wire n80_0;
  wire _w_312;
  wire n41;
  wire _w_364;
  wire _w_305;
  wire n60;
  wire _w_291;
  wire n52_1;
  wire n35;
  wire n22_0;
  wire _w_382;
  wire n72;
  wire n76;
  wire n48;
  wire n33;
  wire _w_255;
  wire n24_5;
  wire _w_289;
  wire n23_6;
  wire _w_359;
  wire n25_2;
  wire n80_1;
  wire n52;
  wire _w_309;
  wire _w_270;
  wire n28;
  wire n25;
  wire n19;
  wire n22_6;
  wire _w_430;
  wire _w_407;
  wire a_4__1;
  wire n20;
  wire _w_391;
  wire n18;
  wire _w_381;
  wire n24_4;
  wire a_1__1;
  wire n39;
  wire _w_254;
  wire _w_415;
  wire n68;
  wire n28_1;
  wire n39_2;
  wire n38;
  wire a_5__3;
  wire _w_357;
  wire _w_349;
  wire n31;
  wire _w_288;
  wire n49_0;
  wire n24_1;
  wire n32;
  wire n25_1;
  wire a_0__2;
  wire _w_295;
  wire n34;
  wire n24_3;
  wire n28_2;
  wire _w_330;
  wire n24;
  wire b_5__2;
  wire n43_1;
  wire _w_397;
  wire n23;
  wire n27;
  wire n21_3;
  wire n24_0;
  wire _w_333;
  wire n37;
  wire n24_7;
  wire n44;
  wire n69;
  wire c_1;
  wire n34_0;
  wire n80;
  wire n68_1;
  wire _w_308;
  wire n34_1;
  wire n20_4;
  wire n34_3;
  wire n49;
  wire n22_1;
  wire n22_3;
  wire a_5__2;
  wire _w_267;
  wire a_5__1;
  wire n22_4;
  wire n22_5;
  wire _w_353;
  wire n20_1;
  wire n20_2;
  wire b_1__4;
  wire _w_281;
  wire a_0__4;
  wire a_0__5;
  wire n20_5;
  wire a_0__1;
  wire n22_2;
  wire n39_0;
  wire n39_1;
  wire a_6__2;
  wire n68_0;
  wire _w_396;
  wire n30;
  wire n38_0;
  wire a_4__0;
  wire _w_299;
  wire n37_0;
  wire n45;
  wire n37_1;
  wire n67;
  wire n51;
  wire _w_256;
  wire a_3__2;
  wire n50;
  wire n37_2;
  wire _w_432;
  wire _w_331;
  wire n29;
  wire n37_3;
  wire _w_328;
  wire n20_0;
  wire n37_4;
  wire _w_387;
  wire c_0;
  wire c_2;
  wire n28_3;
  wire b_6__0;
  wire _w_278;
  wire b_6__2;
  wire _w_373;
  wire b_2__0;
  wire b_6__3;
  wire b_6__5;
  wire _w_352;
  wire b_5__1;
  wire b_5__3;
  wire _w_351;
  wire b_5__4;
  wire _w_356;
  wire b_7__0;
  wire b_5__0;
  wire b_4__0;
  wire b_4__1;
  wire b_4__2;
  wire n23_3;
  wire n23_7;
  wire b_4__3;
  wire _w_410;
  wire n25_4;
  wire b_4__5;
  wire b_3__0;
  wire b_3__1;
  wire n53_1;
  wire b_2__1;
  wire a_2__1;
  wire b_2__2;
  wire b_1__0;
  wire _w_290;
  wire b_1__1;
  wire n34_2;
  wire n23_2;
  wire b_1__2;
  wire b_0__0;
  wire _w_422;
  wire _w_376;
  wire _w_252;
  wire n25_3;
  wire b_0__2;
  wire a_6__3;
  wire b_0__3;
  wire _w_442;
  wire b_0__4;
  wire _w_344;
  wire n81;
  wire b_3__2;
  wire a_7__0;
  wire _w_315;
  wire a_1__0;
  wire n73;
  wire a_7__1;
  wire n18_0;
  wire a_6__0;
  wire a_6__1;
  wire n23_0;
  wire _w_339;
  wire _w_249;
  wire n23_1;
  wire n23_5;
  wire n23_9;
  wire a_5__4;
  wire n84;
  wire a_3__0;
  wire a_3__1;
  wire n23_8;
  wire a_2__2;
  wire a_4__3;
  wire n49_2;
  wire n38_1;
  wire a_1__3;
  wire a_1__4;
  wire n21_0;
  wire n21_2;
  wire _w_420;
  wire b_0__1;
  wire n21_4;
  wire n54;
  wire n21_5;
  wire _w_273;
  wire n18_1;
  wire a_0__3;
  wire n21_6;
  wire _w_251;
  wire _w_250;

  bfr _b_325 (
      .a(_w_444),
      .q(_w_445)
  );
  bfr _b_322 (
      .a(_w_441),
      .q(_w_442)
  );
  bfr _b_321 (
      .a(_w_440),
      .q(_w_441)
  );
  bfr _b_319 (
      .a(_w_438),
      .q(_w_439)
  );
  bfr _b_317 (
      .a(b_6),
      .q(_w_437)
  );
  bfr _b_312 (
      .a(_w_431),
      .q(_w_432)
  );
  bfr _b_311 (
      .a(_w_430),
      .q(_w_431)
  );
  bfr _b_309 (
      .a(_w_428),
      .q(_w_429)
  );
  bfr _b_307 (
      .a(_w_426),
      .q(_w_419)
  );
  bfr _b_304 (
      .a(_w_423),
      .q(_w_424)
  );
  bfr _b_302 (
      .a(_w_421),
      .q(_w_422)
  );
  bfr _b_300 (
      .a(b_4),
      .q(_w_420)
  );
  bfr _b_298 (
      .a(_w_417),
      .q(_w_418)
  );
  bfr _b_296 (
      .a(b_3),
      .q(_w_416)
  );
  bfr _b_291 (
      .a(_w_410),
      .q(_w_399)
  );
  bfr _b_290 (
      .a(_w_409),
      .q(_w_410)
  );
  bfr _b_315 (
      .a(_w_434),
      .q(_w_435)
  );
  bfr _b_289 (
      .a(_w_408),
      .q(_w_409)
  );
  bfr _b_288 (
      .a(_w_407),
      .q(_w_408)
  );
  bfr _b_287 (
      .a(_w_406),
      .q(_w_407)
  );
  bfr _b_286 (
      .a(_w_405),
      .q(_w_406)
  );
  bfr _b_285 (
      .a(_w_404),
      .q(_w_405)
  );
  bfr _b_282 (
      .a(_w_401),
      .q(_w_402)
  );
  bfr _b_281 (
      .a(_w_400),
      .q(_w_401)
  );
  bfr _b_279 (
      .a(_w_398),
      .q(_w_390)
  );
  bfr _b_278 (
      .a(_w_397),
      .q(_w_398)
  );
  bfr _b_277 (
      .a(_w_396),
      .q(_w_397)
  );
  bfr _b_272 (
      .a(_w_391),
      .q(_w_392)
  );
  bfr _b_269 (
      .a(_w_388),
      .q(_w_389)
  );
  bfr _b_268 (
      .a(_w_387),
      .q(_w_388)
  );
  bfr _b_267 (
      .a(_w_386),
      .q(_w_387)
  );
  bfr _b_264 (
      .a(_w_383),
      .q(_w_384)
  );
  bfr _b_327 (
      .a(_w_446),
      .q(_w_447)
  );
  bfr _b_261 (
      .a(_w_380),
      .q(_w_381)
  );
  bfr _b_260 (
      .a(_w_379),
      .q(_w_380)
  );
  bfr _b_323 (
      .a(_w_442),
      .q(_w_443)
  );
  bfr _b_259 (
      .a(a_3),
      .q(_w_379)
  );
  bfr _b_258 (
      .a(_w_377),
      .q(_w_375)
  );
  bfr _b_257 (
      .a(_w_376),
      .q(_w_377)
  );
  spl2 a_1__s_0 (
      .a (_w_374),
      .q0(a_1__0),
      .q1(a_1__1)
  );
  or_bb g41 (
      .a(n20_3),
      .b(n34_2),
      .q(n41)
  );
  bfr _b_164 (
      .a(_w_283),
      .q(_w_284)
  );
  bfr _b_256 (
      .a(a_2),
      .q(_w_376)
  );
  spl3L g23_s_3 (
      .a (n23_6),
      .q0(n23_7),
      .q1(n23_8),
      .q2(_w_372)
  );
  bfr _b_263 (
      .a(a_4),
      .q(_w_383)
  );
  spl2 g23_s_1 (
      .a (n23_0),
      .q0(n23_3),
      .q1(n23_4)
  );
  spl3L b_2__s_0 (
      .a (_w_412),
      .q0(b_2__0),
      .q1(b_2__1),
      .q2(_w_370)
  );
  bfr _b_316 (
      .a(_w_435),
      .q(_w_427)
  );
  and_bb g73 (
      .a(a_5__1),
      .b(b_5__2),
      .q(n73)
  );
  bfr _b_242 (
      .a(_w_361),
      .q(_w_362)
  );
  bfr _b_328 (
      .a(_w_447),
      .q(_w_436)
  );
  bfr _b_225 (
      .a(_w_344),
      .q(_w_345)
  );
  bfr _b_139 (
      .a(_w_258),
      .q(_w_259)
  );
  bfr _b_173 (
      .a(_w_292),
      .q(_w_293)
  );
  spl2 g38_s_0 (
      .a (n38),
      .q0(n38_0),
      .q1(n38_1)
  );
  spl2 g68_s_0 (
      .a (n68),
      .q0(n43_2),
      .q1(n68_1)
  );
  maj_bbi g59 (
      .a(n37_4),
      .b(n58),
      .c(n38_1),
      .q(_w_354)
  );
  and_bb g52 (
      .a(n49_0),
      .b(n51),
      .q(n52)
  );
  spl3L g23_s_0 (
      .a (n23),
      .q0(n23_0),
      .q1(n23_1),
      .q2(n23_2)
  );
  maj_bbi g45 (
      .a(b_4__5),
      .b(n44),
      .c(n23_2),
      .q(n45)
  );
  spl4L g39_s_0 (
      .a (n39),
      .q0(n39_0),
      .q1(n20_4),
      .q2(n39_2),
      .q3(_w_353)
  );
  bfr _b_186 (
      .a(_w_305),
      .q(_w_306)
  );
  bfr _b_199 (
      .a(_w_318),
      .q(_w_319)
  );
  spl2 b_7__s_0 (
      .a (b_7),
      .q0(b_7__0),
      .q1(b_7__1)
  );
  spl4L g20_s_1 (
      .a (n20_1),
      .q0(n20_2),
      .q1(n20_3),
      .q2(n39_1),
      .q3(n20_5)
  );
  bfr _b_191 (
      .a(_w_310),
      .q(n25_1)
  );
  spl4L g34_s_0 (
      .a (n34),
      .q0(n34_0),
      .q1(n34_1),
      .q2(n34_2),
      .q3(n34_3)
  );
  spl2 a_5__s_1 (
      .a (a_5__2),
      .q0(a_5__3),
      .q1(_w_373)
  );
  spl2 g24_s_1 (
      .a (n24_0),
      .q0(n24_3),
      .q1(_w_350)
  );
  spl4L g25_s_1 (
      .a (n25_1),
      .q0(n25_2),
      .q1(n52_2),
      .q2(n25_4),
      .q3(_w_349)
  );
  bfr _b_262 (
      .a(_w_381),
      .q(_w_378)
  );
  spl3L g52_s_0 (
      .a (n52),
      .q0(n52_0),
      .q1(n53_1),
      .q2(n84_0)
  );
  spl3L g28_s_0 (
      .a (n28),
      .q0(n28_0),
      .q1(n28_1),
      .q2(_w_348)
  );
  bfr _b_280 (
      .a(a_6),
      .q(_w_400)
  );
  spl3L g22_s_2 (
      .a (n22_3),
      .q0(n22_4),
      .q1(n22_5),
      .q2(_w_347)
  );
  spl4L g42_s_0 (
      .a (n42),
      .q0(n42_0),
      .q1(n28_3),
      .q2(n21_6),
      .q3(_w_346)
  );
  spl2 g18_s_0 (
      .a (n18),
      .q0(n18_0),
      .q1(_w_343)
  );
  bfr _b_293 (
      .a(b_2),
      .q(_w_413)
  );
  spl3L g24_s_0 (
      .a (n24),
      .q0(n24_0),
      .q1(n24_1),
      .q2(n24_2)
  );
  bfr _b_190 (
      .a(n50),
      .q(_w_310)
  );
  bfr _b_229 (
      .a(n28_1),
      .q(n28_2)
  );
  bfr _b_236 (
      .a(_w_355),
      .q(_w_356)
  );
  spl2 b_1__s_0 (
      .a (_w_411),
      .q0(b_1__0),
      .q1(b_1__1)
  );
  maj_bbi g44 (
      .a(a_4__3),
      .b(_w_270),
      .c(_w_334),
      .q(n44)
  );
  bfr _b_193 (
      .a(_w_312),
      .q(_w_313)
  );
  bfr _b_204 (
      .a(_w_323),
      .q(a_4__3)
  );
  spl2 g53_s_0 (
      .a (n53),
      .q0(n53_0),
      .q1(_w_341)
  );
  spl2 g74_s_0 (
      .a (n74),
      .q0(n74_0),
      .q1(n46_2)
  );
  bfr _b_239 (
      .a(_w_358),
      .q(_w_359)
  );
  spl2 g80_s_0 (
      .a (n80),
      .q0(n49_2),
      .q1(n80_1)
  );
  bfr _b_314 (
      .a(_w_433),
      .q(_w_434)
  );
  maj_bbb g21 (
      .a(a_2__2),
      .b(b_2__2),
      .c(_w_330),
      .q(n21)
  );
  maj_bbb g85 (
      .a(n25_3),
      .b(n52_2),
      .c(n84_0),
      .q(n85)
  );
  maj_bbi g83 (
      .a(n24_7),
      .b(n82),
      .c(n81),
      .q(_w_338)
  );
  spl2 b_6__s_1 (
      .a (b_6__0),
      .q0(b_6__4),
      .q1(_w_337)
  );
  bfr _b_159 (
      .a(_w_278),
      .q(_w_279)
  );
  spl3L g21_s_1 (
      .a (n21_0),
      .q0(n21_2),
      .q1(n21_3),
      .q2(_w_336)
  );
  maj_bbi g82 (
      .a(n49_2),
      .b(_w_322),
      .c(n24_6),
      .q(n82)
  );
  bfr _b_231 (
      .a(n24_3),
      .q(n24_4)
  );
  bfr _b_243 (
      .a(_w_362),
      .q(_w_363)
  );
  spl4L a_6__s_0 (
      .a (_w_399),
      .q0(a_6__0),
      .q1(a_6__1),
      .q2(a_6__2),
      .q3(_w_335)
  );
  spl2 b_4__s_1 (
      .a (b_4__0),
      .q0(b_4__4),
      .q1(_w_334)
  );
  bfr _b_273 (
      .a(_w_392),
      .q(_w_393)
  );
  bfr _b_219 (
      .a(_w_338),
      .q(_w_339)
  );
  maj_bbb g81 (
      .a(n24_5),
      .b(n49_1),
      .c(n80_1),
      .q(n81)
  );
  spl3L a_2__s_0 (
      .a (_w_375),
      .q0(a_2__0),
      .q1(a_2__1),
      .q2(_w_333)
  );
  bfr _b_136 (
      .a(_w_255),
      .q(_w_256)
  );
  spl2 g20_s_0 (
      .a (n20),
      .q0(n20_0),
      .q1(_w_330)
  );
  bfr _b_151 (
      .a(n22_2),
      .q(n22_3)
  );
  or_bb g78 (
      .a(a_6__1),
      .b(b_6__2),
      .q(n78)
  );
  bfr _b_237 (
      .a(_w_356),
      .q(_w_357)
  );
  maj_bbi g75 (
      .a(n23_7),
      .b(n74_0),
      .c(n46_1),
      .q(n76)
  );
  maj_bbi g71 (
      .a(n22_6),
      .b(n70),
      .c(n69),
      .q(_w_324)
  );
  bfr _b_297 (
      .a(_w_416),
      .q(_w_417)
  );
  bfr _b_208 (
      .a(_w_327),
      .q(_w_328)
  );
  maj_bbi g70 (
      .a(n43_2),
      .b(n68_0),
      .c(_w_347),
      .q(n70)
  );
  spl4L a_4__s_0 (
      .a (_w_382),
      .q0(a_4__0),
      .q1(a_4__1),
      .q2(a_4__2),
      .q3(_w_323)
  );
  maj_bbb g69 (
      .a(n22_4),
      .b(n43_1),
      .c(n68_1),
      .q(n69)
  );
  spl3L g49_s_0 (
      .a (n49),
      .q0(n49_0),
      .q1(n49_1),
      .q2(n24_6)
  );
  bfr _b_294 (
      .a(_w_413),
      .q(_w_414)
  );
  bfr _b_137 (
      .a(_w_256),
      .q(s_3)
  );
  bfr _b_195 (
      .a(_w_314),
      .q(_w_315)
  );
  or_bb g66 (
      .a(a_4__1),
      .b(b_4__2),
      .q(n66)
  );
  spl3L g24_s_2 (
      .a (n24_4),
      .q0(n24_5),
      .q1(n80_0),
      .q2(_w_322)
  );
  maj_bbi g64 (
      .a(n42_1),
      .b(n42_2),
      .c(n21_6),
      .q(n42_3)
  );
  maj_bbi g62 (
      .a(n60),
      .b(n61),
      .c(n39_3),
      .q(_w_311)
  );
  and_bb g67 (
      .a(a_4__2),
      .b(b_4__3),
      .q(n67)
  );
  bfr _b_224 (
      .a(n18_0),
      .q(_w_344)
  );
  bfr _b_253 (
      .a(_w_372),
      .q(n75)
  );
  maj_bbi g61 (
      .a(n34_0),
      .b(n39_2),
      .c(n20_5),
      .q(n39_3)
  );
  bfr _b_201 (
      .a(_w_320),
      .q(_w_321)
  );
  spl3L b_0__s_0 (
      .a (b_0),
      .q0(b_0__0),
      .q1(b_0__1),
      .q2(b_0__2)
  );
  bfr _b_198 (
      .a(_w_317),
      .q(_w_318)
  );
  or_bb g72 (
      .a(a_5__0),
      .b(b_5__1),
      .q(n72)
  );
  bfr _b_131 (
      .a(_w_250),
      .q(_w_251)
  );
  bfr _b_215 (
      .a(b_4__4),
      .q(b_4__5)
  );
  or_bb g55 (
      .a(n18_1),
      .b(n54),
      .q(cout)
  );
  maj_bbb g54 (
      .a(n25_2),
      .b(n52_1),
      .c(n53_1),
      .q(n54)
  );
  spl3L b_1__s_1 (
      .a (b_1__1),
      .q0(b_1__2),
      .q1(b_1__3),
      .q2(n37_0)
  );
  or_bb g53 (
      .a(a_7__1),
      .b(b_7__1),
      .q(_w_296)
  );
  bfr _b_142 (
      .a(_w_261),
      .q(_w_262)
  );
  maj_bbi g87 (
      .a(n25_5),
      .b(n86),
      .c(n85),
      .q(s_7)
  );
  bfr _b_295 (
      .a(_w_414),
      .q(_w_412)
  );
  bfr _b_145 (
      .a(_w_264),
      .q(_w_265)
  );
  and_bi g80 (
      .a(n78),
      .b(n79),
      .q(n80)
  );
  and_bi g84 (
      .a(n53_0),
      .b(_w_343),
      .q(n84)
  );
  spl2 g22_s_0 (
      .a (n22),
      .q0(n22_0),
      .q1(n22_1)
  );
  maj_bbi g40 (
      .a(n20_2),
      .b(n34_1),
      .c(_w_353),
      .q(n40)
  );
  and_bb g49 (
      .a(n46_0),
      .b(n48),
      .q(n49)
  );
  bfr _b_251 (
      .a(b_2__0),
      .q(b_2__2)
  );
  maj_bbi g47 (
      .a(a_5__4),
      .b(b_5__4),
      .c(n23_4),
      .q(n47)
  );
  bfr _b_161 (
      .a(_w_280),
      .q(_w_281)
  );
  spl3L c_s_0 (
      .a (cin),
      .q0(c_0),
      .q1(c_1),
      .q2(_w_332)
  );
  spl3L a_5__s_0 (
      .a (_w_390),
      .q0(a_5__0),
      .q1(a_5__1),
      .q2(a_5__2)
  );
  bfr _b_221 (
      .a(a_0__4),
      .q(a_0__5)
  );
  spl3L a_0__s_1 (
      .a (a_0__2),
      .q0(a_0__3),
      .q1(a_0__4),
      .q2(_w_340)
  );
  maj_bbi g77 (
      .a(n75),
      .b(n76),
      .c(n23_9),
      .q(_w_292)
  );
  and_bi g42 (
      .a(n41),
      .b(n40),
      .q(n42)
  );
  maj_bbb g25 (
      .a(a_6__0),
      .b(b_6__1),
      .c(n24_1),
      .q(n25)
  );
  maj_bbi g60 (
      .a(n20_4),
      .b(n39_1),
      .c(n34_3),
      .q(n61)
  );
  and_bi g34 (
      .a(n32),
      .b(n33),
      .q(n34)
  );
  bfr _b_308 (
      .a(b_5),
      .q(_w_428)
  );
  bfr _b_153 (
      .a(_w_272),
      .q(b_3__2)
  );
  and_bi g39 (
      .a(n38_0),
      .b(n36),
      .q(n39)
  );
  spl3L b_5__s_0 (
      .a (_w_427),
      .q0(b_5__0),
      .q1(b_5__1),
      .q2(b_5__2)
  );
  spl2 g23_s_2 (
      .a (n23_3),
      .q0(n23_5),
      .q1(n23_6)
  );
  bfr _b_227 (
      .a(n42_0),
      .q(n63)
  );
  maj_bbb g38 (
      .a(a_1__3),
      .b(_w_351),
      .c(n37_0),
      .q(n38)
  );
  and_bb g46 (
      .a(n43_0),
      .b(n45),
      .q(n46)
  );
  maj_bbb g37 (
      .a(a_0__1),
      .b(b_0__2),
      .c(_w_332),
      .q(n37)
  );
  maj_bbi g76 (
      .a(n23_8),
      .b(n46_2),
      .c(n74_1),
      .q(n23_9)
  );
  bfr _b_148 (
      .a(_w_267),
      .q(_w_268)
  );
  bfr _b_217 (
      .a(n21_3),
      .q(n21_4)
  );
  maj_bbb g36 (
      .a(a_1__0),
      .b(b_1__0),
      .c(n35),
      .q(_w_290)
  );
  bfr _b_141 (
      .a(_w_260),
      .q(_w_261)
  );
  bfr _b_181 (
      .a(_w_300),
      .q(_w_301)
  );
  maj_bbi g35 (
      .a(a_0__0),
      .b(b_0__1),
      .c(c_1),
      .q(n35)
  );
  maj_bbi g57 (
      .a(a_0__5),
      .b(n56),
      .c(n37_2),
      .q(_w_274)
  );
  bfr _b_305 (
      .a(_w_424),
      .q(_w_425)
  );
  bfr _b_299 (
      .a(_w_418),
      .q(_w_415)
  );
  bfr _b_169 (
      .a(_w_288),
      .q(_w_289)
  );
  bfr _b_180 (
      .a(_w_299),
      .q(_w_300)
  );
  bfr _b_326 (
      .a(_w_445),
      .q(_w_446)
  );
  spl4L b_6__s_0 (
      .a (_w_436),
      .q0(b_6__0),
      .q1(b_6__1),
      .q2(b_6__2),
      .q3(b_6__3)
  );
  or_bb g31 (
      .a(n29),
      .b(n30),
      .q(n31)
  );
  and_bi g30 (
      .a(n28_0),
      .b(_w_336),
      .q(n30)
  );
  spl3L a_1__s_1 (
      .a (a_1__1),
      .q0(a_1__2),
      .q1(_w_371),
      .q2(_w_351)
  );
  spl2 g37_s_1 (
      .a (n37_1),
      .q0(n37_3),
      .q1(_w_331)
  );
  bfr _b_170 (
      .a(_w_289),
      .q(s_0)
  );
  and_bi g29 (
      .a(n21_2),
      .b(_w_348),
      .q(n29)
  );
  bfr _b_133 (
      .a(_w_252),
      .q(_w_253)
  );
  and_bi g28 (
      .a(n26),
      .b(n27),
      .q(n28)
  );
  and_bb g27 (
      .a(a_3__1),
      .b(_w_271),
      .q(n27)
  );
  bfr _b_324 (
      .a(_w_443),
      .q(_w_444)
  );
  or_bb g26 (
      .a(a_3__0),
      .b(b_3__1),
      .q(n26)
  );
  bfr _b_275 (
      .a(_w_394),
      .q(_w_395)
  );
  maj_bbi g86 (
      .a(n52_0),
      .b(n84_1),
      .c(_w_349),
      .q(n86)
  );
  bfr _b_165 (
      .a(_w_284),
      .q(_w_285)
  );
  spl3L b_3__s_0 (
      .a (_w_415),
      .q0(b_3__0),
      .q1(b_3__1),
      .q2(_w_271)
  );
  maj_bbi g51 (
      .a(b_6__5),
      .b(_w_309),
      .c(n25_0),
      .q(n51)
  );
  spl2 g21_s_0 (
      .a (n21),
      .q0(n21_0),
      .q1(n21_1)
  );
  bfr _b_196 (
      .a(_w_315),
      .q(_w_316)
  );
  bfr _b_203 (
      .a(n80_0),
      .q(n24_7)
  );
  spl3L a_0__s_0 (
      .a (a_0),
      .q0(a_0__0),
      .q1(a_0__1),
      .q2(a_0__2)
  );
  maj_bbb g24 (
      .a(a_5__3),
      .b(_w_273),
      .c(n23_1),
      .q(n24)
  );
  bfr _b_144 (
      .a(_w_263),
      .q(_w_264)
  );
  bfr _b_222 (
      .a(_w_341),
      .q(_w_342)
  );
  maj_bbb g23 (
      .a(a_4__0),
      .b(b_4__1),
      .c(n22_1),
      .q(n23)
  );
  spl2 g22_s_1 (
      .a (n22_0),
      .q0(n22_2),
      .q1(_w_270)
  );
  bfr _b_283 (
      .a(_w_402),
      .q(_w_403)
  );
  and_bi g68 (
      .a(n66),
      .b(n67),
      .q(n68)
  );
  bfr _b_245 (
      .a(_w_364),
      .q(_w_365)
  );
  bfr _b_266 (
      .a(_w_385),
      .q(_w_386)
  );
  spl2 g25_s_0 (
      .a (n25),
      .q0(n50),
      .q1(_w_309)
  );
  bfr _b_168 (
      .a(_w_287),
      .q(_w_288)
  );
  and_bb g43 (
      .a(n31),
      .b(_w_346),
      .q(n43)
  );
  maj_bbi g63 (
      .a(n21_5),
      .b(n28_4),
      .c(n28_3),
      .q(n64)
  );
  spl3L g37_s_0 (
      .a (n37),
      .q0(a_1__3),
      .q1(n37_1),
      .q2(n37_2)
  );
  bfr _b_246 (
      .a(_w_365),
      .q(_w_366)
  );
  maj_bbi g58 (
      .a(a_1__4),
      .b(b_1__4),
      .c(_w_331),
      .q(n58)
  );
  bfr _b_143 (
      .a(_w_262),
      .q(_w_263)
  );
  bfr _b_197 (
      .a(_w_316),
      .q(_w_317)
  );
  bfr _b_162 (
      .a(_w_281),
      .q(_w_282)
  );
  or_bb g32 (
      .a(a_2__0),
      .b(b_2__1),
      .q(n32)
  );
  and_bb g19 (
      .a(a_0__3),
      .b(b_0__4),
      .q(n19)
  );
  bfr _b_301 (
      .a(_w_420),
      .q(_w_421)
  );
  and_bb g33 (
      .a(a_2__1),
      .b(_w_370),
      .q(n33)
  );
  and_bb g18 (
      .a(a_7__0),
      .b(b_7__0),
      .q(_w_257)
  );
  spl2 b_0__s_1 (
      .a (b_0__0),
      .q0(b_0__3),
      .q1(b_0__4)
  );
  and_bb g79 (
      .a(a_6__2),
      .b(b_6__3),
      .q(n79)
  );
  bfr _b_130 (
      .a(_w_249),
      .q(_w_250)
  );
  spl2 g84_s_0 (
      .a (n84),
      .q0(n25_3),
      .q1(n84_1)
  );
  maj_bbb g20 (
      .a(a_1__2),
      .b(b_1__3),
      .c(n19),
      .q(n20)
  );
  spl2 g21_s_2 (
      .a (n21_4),
      .q0(n21_5),
      .q1(n42_2)
  );
  bfr _b_202 (
      .a(_w_321),
      .q(s_2)
  );
  bfr _b_212 (
      .a(n37_3),
      .q(n37_4)
  );
  bfr _b_132 (
      .a(_w_251),
      .q(_w_252)
  );
  bfr _b_134 (
      .a(_w_253),
      .q(_w_254)
  );
  bfr _b_135 (
      .a(_w_254),
      .q(_w_255)
  );
  bfr _b_140 (
      .a(_w_259),
      .q(_w_260)
  );
  bfr _b_265 (
      .a(_w_384),
      .q(_w_385)
  );
  bfr _b_146 (
      .a(_w_265),
      .q(_w_266)
  );
  bfr _b_147 (
      .a(_w_266),
      .q(_w_267)
  );
  spl3L g46_s_0 (
      .a (n46),
      .q0(n46_0),
      .q1(n46_1),
      .q2(n74_1)
  );
  bfr _b_149 (
      .a(_w_268),
      .q(_w_269)
  );
  maj_bbi g50 (
      .a(a_6__3),
      .b(_w_350),
      .c(_w_337),
      .q(n25_0)
  );
  maj_bbi g65 (
      .a(n63),
      .b(n64),
      .c(n42_3),
      .q(_w_249)
  );
  bfr _b_216 (
      .a(_w_335),
      .q(a_6__3)
  );
  bfr _b_150 (
      .a(_w_269),
      .q(n18)
  );
  spl2 b_5__s_1 (
      .a (b_5__0),
      .q0(b_5__3),
      .q1(_w_273)
  );
  bfr _b_154 (
      .a(b_5__3),
      .q(b_5__4)
  );
  bfr _b_313 (
      .a(_w_432),
      .q(_w_433)
  );
  bfr _b_292 (
      .a(b_1),
      .q(_w_411)
  );
  bfr _b_152 (
      .a(b_3__0),
      .q(_w_272)
  );
  bfr _b_172 (
      .a(_w_291),
      .q(n36)
  );
  bfr _b_155 (
      .a(_w_274),
      .q(_w_275)
  );
  bfr _b_156 (
      .a(_w_275),
      .q(_w_276)
  );
  bfr _b_138 (
      .a(_w_257),
      .q(_w_258)
  );
  bfr _b_157 (
      .a(_w_276),
      .q(_w_277)
  );
  spl3L g43_s_0 (
      .a (n43),
      .q0(n43_0),
      .q1(n43_1),
      .q2(n68_0)
  );
  bfr _b_187 (
      .a(_w_306),
      .q(_w_307)
  );
  bfr _b_207 (
      .a(_w_326),
      .q(_w_327)
  );
  bfr _b_158 (
      .a(_w_277),
      .q(_w_278)
  );
  maj_bbi g48 (
      .a(n23_5),
      .b(n47),
      .c(n24_2),
      .q(n48)
  );
  bfr _b_163 (
      .a(_w_282),
      .q(_w_283)
  );
  bfr _b_166 (
      .a(_w_285),
      .q(_w_286)
  );
  bfr _b_174 (
      .a(_w_293),
      .q(_w_294)
  );
  bfr _b_271 (
      .a(a_5),
      .q(_w_391)
  );
  bfr _b_179 (
      .a(_w_298),
      .q(_w_299)
  );
  bfr _b_175 (
      .a(_w_294),
      .q(_w_295)
  );
  bfr _b_255 (
      .a(a_1),
      .q(_w_374)
  );
  bfr _b_176 (
      .a(_w_295),
      .q(s_5)
  );
  bfr _b_177 (
      .a(_w_296),
      .q(_w_297)
  );
  bfr _b_250 (
      .a(_w_369),
      .q(a_3__2)
  );
  bfr _b_320 (
      .a(_w_439),
      .q(_w_440)
  );
  bfr _b_182 (
      .a(_w_301),
      .q(_w_302)
  );
  bfr _b_183 (
      .a(_w_302),
      .q(_w_303)
  );
  bfr _b_184 (
      .a(_w_303),
      .q(_w_304)
  );
  bfr _b_185 (
      .a(_w_304),
      .q(_w_305)
  );
  bfr _b_310 (
      .a(_w_429),
      .q(_w_430)
  );
  bfr _b_238 (
      .a(_w_357),
      .q(_w_358)
  );
  bfr _b_188 (
      .a(_w_307),
      .q(_w_308)
  );
  bfr _b_178 (
      .a(_w_297),
      .q(_w_298)
  );
  bfr _b_189 (
      .a(_w_308),
      .q(n53)
  );
  and_bi g74 (
      .a(n72),
      .b(n73),
      .q(_w_352)
  );
  bfr _b_192 (
      .a(_w_311),
      .q(_w_312)
  );
  bfr _b_171 (
      .a(_w_290),
      .q(_w_291)
  );
  bfr _b_194 (
      .a(_w_313),
      .q(_w_314)
  );
  spl4L b_4__s_0 (
      .a (_w_419),
      .q0(b_4__0),
      .q1(b_4__1),
      .q2(b_4__2),
      .q3(b_4__3)
  );
  bfr _b_200 (
      .a(_w_319),
      .q(_w_320)
  );
  bfr _b_235 (
      .a(_w_354),
      .q(_w_355)
  );
  bfr _b_167 (
      .a(_w_286),
      .q(_w_287)
  );
  bfr _b_205 (
      .a(_w_324),
      .q(_w_325)
  );
  bfr _b_206 (
      .a(_w_325),
      .q(_w_326)
  );
  bfr _b_270 (
      .a(_w_389),
      .q(_w_382)
  );
  spl2 g28_s_1 (
      .a (n28_2),
      .q0(n42_1),
      .q1(n28_4)
  );
  maj_bbb g22 (
      .a(a_3__2),
      .b(b_3__2),
      .c(n21_1),
      .q(n22)
  );
  bfr _b_160 (
      .a(_w_279),
      .q(_w_280)
  );
  bfr _b_210 (
      .a(_w_329),
      .q(s_4)
  );
  bfr _b_211 (
      .a(n20_0),
      .q(n20_1)
  );
  bfr _b_306 (
      .a(_w_425),
      .q(_w_426)
  );
  bfr _b_213 (
      .a(c_0),
      .q(c_2)
  );
  bfr _b_276 (
      .a(_w_395),
      .q(_w_396)
  );
  bfr _b_214 (
      .a(_w_333),
      .q(a_2__2)
  );
  bfr _b_218 (
      .a(b_6__4),
      .q(b_6__5)
  );
  spl2 a_7__s_0 (
      .a (a_7),
      .q0(a_7__0),
      .q1(a_7__1)
  );
  bfr _b_220 (
      .a(_w_339),
      .q(s_6)
  );
  bfr _b_230 (
      .a(n25_4),
      .q(n25_5)
  );
  bfr _b_241 (
      .a(_w_360),
      .q(_w_361)
  );
  bfr _b_226 (
      .a(_w_345),
      .q(n18_1)
  );
  bfr _b_247 (
      .a(_w_366),
      .q(_w_367)
  );
  maj_bbi g56 (
      .a(b_0__3),
      .b(c_2),
      .c(_w_340),
      .q(n56)
  );
  bfr _b_228 (
      .a(n22_5),
      .q(n22_6)
  );
  bfr _b_232 (
      .a(_w_371),
      .q(a_1__4)
  );
  bfr _b_233 (
      .a(_w_352),
      .q(n74)
  );
  bfr _b_318 (
      .a(_w_437),
      .q(_w_438)
  );
  bfr _b_234 (
      .a(n39_0),
      .q(n60)
  );
  bfr _b_240 (
      .a(_w_359),
      .q(_w_360)
  );
  bfr _b_244 (
      .a(_w_363),
      .q(_w_364)
  );
  bfr _b_223 (
      .a(_w_342),
      .q(n52_1)
  );
  bfr _b_249 (
      .a(_w_368),
      .q(_w_369)
  );
  bfr _b_284 (
      .a(_w_403),
      .q(_w_404)
  );
  bfr _b_248 (
      .a(_w_367),
      .q(s_1)
  );
  bfr _b_274 (
      .a(_w_393),
      .q(_w_394)
  );
  spl3L a_3__s_0 (
      .a (_w_378),
      .q0(a_3__0),
      .q1(a_3__1),
      .q2(_w_368)
  );
  bfr _b_209 (
      .a(_w_328),
      .q(_w_329)
  );
  bfr _b_252 (
      .a(b_1__2),
      .q(b_1__4)
  );
  bfr _b_303 (
      .a(_w_422),
      .q(_w_423)
  );
  bfr _b_254 (
      .a(_w_373),
      .q(a_5__4)
  );
endmodule
