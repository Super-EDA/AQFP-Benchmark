module comparator (a_0,a_1,a_2,a_3,a_4,a_5,a_6,a_7,b_0,b_1,b_2,b_3,b_4,b_5,b_6,b_7,q);
  input a_0,a_1,a_2,a_3,a_4,a_5,a_6,a_7,b_0,b_1,b_2,b_3,b_4,b_5,b_6,b_7;
  output q;
  wire _w_96,_w_97,_w_92,_w_90,_w_88,_w_86,_w_83,_w_82,a_3_1,a_3_0,a_7_2,a_7_0,_w_94,a_4_0,a_5_2,a_6_3,_w_85,a_6_2,b_2_1,b_2_0,b_3_1,b_3_0,n35,_w_98,b_6_2,a_4_3,a_5_0,n26,n33,n39,b_7_0,a_6_1,b_4_1,b_5_2,n24,b_7_2,_w_87,a_2_1,a_2_0,_w_91,n23_1,b_7_1,n17,n18,n19,n20,b_4_0,n21,b_6_3,n23,n37,_w_81,a_4_2,a_6_0,b_4_3,a_5_1,n23_0,n25,n27,a_4_1,n28,_w_93,n42,n38,n29,n41,_w_89,n30,n32,a_7_1,b_6_0,_w_95,n22,n34,n36,_w_84,n40,b_6_1,n31,b_5_0,b_5_1,b_4_2;

  bfr _b_61(.a(b_3),.q(_w_98));
  bfr _b_60(.a(b_1),.q(_w_97));
  bfr _b_59(.a(a_3),.q(_w_96));
  and_bi g17(.a(a_6_0),.b(b_6_1),.q(b_7_2));
  maj_bbi g29(.a(a_4_2),.b(b_4_3),.c(b_4_2),.q(n29));
  maj_bbi g20(.a(a_6_2),.b(b_6_3),.c(b_6_2),.q(n20));
  maj_bbi g22(.a(n19),.b(n21),.c(a_6_3),.q(n22));
  or_bb g23(.a(n20),.b(n22),.q(n23));
  and_bi g24(.a(a_4_0),.b(b_4_1),.q(b_5_2));
  or_bb g40(.a(n23_1),.b(n39),.q(n40));
  and_bi g42(.a(n41),.b(n27),.q(n42));
  maj_bbi g25(.a(a_5_2),.b(n24),.c(b_5_2),.q(_w_90));
  bfr _b_57(.a(_w_94),.q(n18));
  and_bi g28(.a(a_5_0),.b(_w_85),.q(b_4_2));
  or_bb g41(.a(n32),.b(n40),.q(n41));
  maj_bbi g31(.a(n28),.b(n30),.c(a_4_3),.q(n31));
  and_bi g21(.a(b_7_0),.b(_w_82),.q(n21));
  or_bb g32(.a(n29),.b(n31),.q(_w_88));
  and_bi g38(.a(b_3_0),.b(a_3_1),.q(n38));
  maj_bbi g18(.a(a_7_2),.b(n17),.c(b_7_2),.q(_w_92));
  and_bi g33(.a(b_0),.b(a_0),.q(_w_95));
  maj_bbi g35(.a(b_2_1),.b(n34),.c(a_2_1),.q(n35));
  maj_bbi g34(.a(_w_97),.b(n33),.c(_w_95),.q(a_2_1));
  bfr _b_48(.a(b_5_1),.q(n24));
  and_bi g36(.a(a_2_0),.b(_w_84),.q(n36));
  spl2 b_6_s_1(.a(b_6_0),.q0(n19),.q1(b_6_3));
  maj_bbi g37(.a(a_3_0),.b(n36),.c(b_3_1),.q(n37));
  spl2 a_6_s_1(.a(a_6_1),.q0(a_6_2),.q1(a_6_3));
  maj_bbi g39(.a(n35),.b(n38),.c(n37),.q(_w_87));
  bfr _b_44(.a(_w_81),.q(n34));
  bfr _b_56(.a(_w_93),.q(_w_94));
  spl2 g23_s_0(.a(n23),.q0(n23_0),.q1(n39));
  spl3L b_7_s_0(.a(b_7),.q0(b_7_0),.q1(b_7_1),.q2(_w_86));
  inv inv_n42(.a(n42),.q(q));
  spl2 b_6_s_0(.a(b_6),.q0(b_6_0),.q1(b_6_1));
  spl3L b_5_s_0(.a(b_5),.q0(b_5_0),.q1(b_5_1),.q2(_w_85));
  or_bb g27(.a(n18),.b(n26),.q(n27));
  spl2 a_3_s_0(.a(_w_96),.q0(a_3_0),.q1(a_3_1));
  spl2 b_4_s_0(.a(b_4),.q0(b_4_0),.q1(b_4_1));
  spl2 b_3_s_0(.a(_w_98),.q0(b_3_0),.q1(b_3_1));
  and_bi g26(.a(n25),.b(n23_0),.q(n26));
  bfr _b_47(.a(b_2_0),.q(b_2_1));
  and_bi g19(.a(a_7_0),.b(_w_86),.q(b_6_2));
  spl2 b_2_s_0(.a(b_2),.q0(b_2_0),.q1(_w_84));
  spl2 a_6_s_0(.a(a_6),.q0(a_6_0),.q1(a_6_1));
  spl3L a_5_s_0(.a(a_5),.q0(a_5_0),.q1(a_5_1),.q2(_w_83));
  spl2 a_4_s_1(.a(a_4_1),.q0(a_4_2),.q1(a_4_3));
  bfr _b_51(.a(_w_88),.q(_w_89));
  spl3L a_7_s_0(.a(a_7),.q0(a_7_0),.q1(a_7_1),.q2(_w_82));
  bfr _b_52(.a(_w_89),.q(n32));
  spl2 a_4_s_0(.a(a_4),.q0(a_4_0),.q1(a_4_1));
  spl2 a_2_s_0(.a(a_2),.q0(a_2_0),.q1(_w_81));
  spl2 b_4_s_1(.a(b_4_0),.q0(n28),.q1(b_4_3));
  bfr _b_45(.a(a_7_1),.q(a_7_2));
  bfr _b_46(.a(a_5_1),.q(a_5_2));
  bfr _b_55(.a(_w_92),.q(_w_93));
  bfr _b_49(.a(b_7_1),.q(n17));
  bfr _b_50(.a(_w_87),.q(n23_1));
  bfr _b_53(.a(_w_90),.q(_w_91));
  and_bi g30(.a(b_5_0),.b(_w_83),.q(n30));
  bfr _b_54(.a(_w_91),.q(n25));
  bfr _b_58(.a(a_1),.q(n33));
endmodule
