module adder_8 (a_0_,a_1_,a_2_,a_3_,a_4_,a_5_,a_6_,a_7_,b_0_,b_1_,b_2_,b_3_,b_4_,b_5_,b_6_,b_7_,c,cout,s_0_,s_1_,s_2_,s_3_,s_4_,s_5_,s_6_,s_7_);
  input a_0_,a_1_,a_2_,a_3_,a_4_,a_5_,a_6_,a_7_,b_0_,b_1_,b_2_,b_3_,b_4_,b_5_,b_6_,b_7_,c;
  output cout,s_0_,s_1_,s_2_,s_3_,s_4_,s_5_,s_6_,s_7_;
  wire _w_447,_w_446,_w_445,_w_444,_w_441,_w_440,_w_439,_w_438,_w_435,_w_433,_w_431,_w_425,_w_424,_w_421,_w_419,_w_416,_w_412,_w_411,_w_409,_w_408,_w_401,_w_399,_w_398,_w_395,_w_393,_w_392,_w_390,_w_394,_w_388,_w_386,_w_385,_w_384,_w_383,_w_375,_w_372,_w_371,_w_370,_w_402,_w_368,_w_400,_w_367,_w_366,_w_389,_w_363,_w_361,_w_360,_w_358,_w_355,_w_354,_w_348,_w_429,_w_347,_w_346,_w_345,_w_343,_w_342,_w_341,_w_340,_w_338,_w_337,_w_417,_w_335,_w_334,_w_329,_w_350,_w_327,_w_427,_w_423,_w_326,_w_325,_w_324,_w_323,_w_322,_w_320,_w_318,_w_317,_w_316,_w_314,_w_313,_w_405,_w_311,_w_365,_w_310,_w_307,_w_304,_w_303,_w_426,_w_302,_w_300,_w_362,_w_298,_w_297,_w_296,_w_406,_w_294,_w_293,_w_292,_w_321,_w_287,_w_286,_w_413,_w_285,_w_283,_w_280,_w_277,_w_276,_w_275,_w_274,_w_272,_w_271,_w_269,_w_268,_w_266,_w_264,_w_261,_w_260,_w_379,_w_258,_w_257,_w_259,n24_2,_w_436,n25_5,_w_336,n24_6,_w_332,_w_253,n52_2,n28_4,n74_1,_w_418,n42_2,n42_1,n56,_w_403,a_1__2,n42_0,_w_279,n43_2,_w_443,n43_0,_w_377,n46_2,_w_265,n21,_w_437,_w_282,n46_0,n23_4,a_0__0,_w_284,n53_0,n53,n74_0,n28_0,_w_263,n49_1,_w_380,n84_1,n78,n36,n39_3,n84_0,n86,b_4__4,n85,_w_404,a_5__0,_w_319,n79,_w_378,n42_3,n26,n75,_w_369,n22,n74,b_6__4,_w_434,n25_0,n70,n20_3,n66,_w_374,n21_1,n64,n63,n61,_w_306,b_1__3,n58,n40,n47,n46,n82,b_7__1,_w_428,n43,_w_301,n42,_w_414,_w_262,a_4__2,a_2__0,n52_0,b_6__1,n46_1,n80_0,_w_312,n41,_w_364,_w_305,n60,_w_291,n52_1,n35,n22_0,_w_382,n72,n76,n48,n33,_w_255,n24_5,_w_289,n23_6,_w_359,n25_2,n80_1,n52,_w_309,_w_270,n28,n25,n19,n22_6,_w_430,_w_407,a_4__1,n20,_w_391,n18,_w_381,n24_4,a_1__1,n39,_w_254,_w_415,n68,n28_1,n39_2,n38,a_5__3,_w_357,_w_349,n31,_w_288,n49_0,n24_1,n32,n25_1,a_0__2,_w_295,n34,n24_3,n28_2,_w_330,n24,b_5__2,n43_1,_w_397,n23,n27,n21_3,n24_0,_w_333,n37,n24_7,n44,n69,c_1,n34_0,n80,n68_1,_w_308,n34_1,n20_4,n34_3,n49,n22_1,n22_3,a_5__2,_w_267,a_5__1,n22_4,n22_5,_w_353,n20_1,n20_2,b_1__4,_w_281,a_0__4,a_0__5,n20_5,a_0__1,n22_2,n39_0,n39_1,a_6__2,n68_0,_w_396,n30,n38_0,a_4__0,_w_299,n37_0,n45,n37_1,n67,n51,_w_256,a_3__2,n50,n37_2,_w_432,_w_331,n29,n37_3,_w_328,n20_0,n37_4,_w_387,c_0,c_2,n28_3,b_6__0,_w_278,b_6__2,_w_373,b_2__0,b_6__3,b_6__5,_w_352,b_5__1,b_5__3,_w_351,b_5__4,_w_356,b_7__0,b_5__0,b_4__0,b_4__1,b_4__2,n23_3,n23_7,b_4__3,_w_410,n25_4,b_4__5,b_3__0,b_3__1,n53_1,b_2__1,a_2__1,b_2__2,b_1__0,_w_290,b_1__1,n34_2,n23_2,b_1__2,b_0__0,_w_422,_w_376,_w_252,n25_3,b_0__2,a_6__3,b_0__3,_w_442,b_0__4,_w_344,n81,b_3__2,a_7__0,_w_315,a_1__0,n73,a_7__1,n18_0,a_6__0,a_6__1,n23_0,_w_339,_w_249,n23_1,n23_5,n23_9,a_5__4,n84,a_3__0,a_3__1,n23_8,a_2__2,a_4__3,n49_2,n38_1,a_1__3,a_1__4,n21_0,n21_2,_w_420,b_0__1,n21_4,n54,n21_5,_w_273,n18_1,a_0__3,n21_6,_w_251,_w_250;

  bfr _b_325(.a(_w_444),.q(_w_445));
  bfr _b_322(.a(_w_441),.q(_w_442));
  bfr _b_321(.a(_w_440),.q(_w_441));
  bfr _b_319(.a(_w_438),.q(_w_439));
  bfr _b_317(.a(b_6_),.q(_w_437));
  bfr _b_312(.a(_w_431),.q(_w_432));
  bfr _b_311(.a(_w_430),.q(_w_431));
  bfr _b_309(.a(_w_428),.q(_w_429));
  bfr _b_307(.a(_w_426),.q(_w_419));
  bfr _b_304(.a(_w_423),.q(_w_424));
  bfr _b_302(.a(_w_421),.q(_w_422));
  bfr _b_300(.a(b_4_),.q(_w_420));
  bfr _b_298(.a(_w_417),.q(_w_418));
  bfr _b_296(.a(b_3_),.q(_w_416));
  bfr _b_291(.a(_w_410),.q(_w_399));
  bfr _b_290(.a(_w_409),.q(_w_410));
  bfr _b_315(.a(_w_434),.q(_w_435));
  bfr _b_289(.a(_w_408),.q(_w_409));
  bfr _b_288(.a(_w_407),.q(_w_408));
  bfr _b_287(.a(_w_406),.q(_w_407));
  bfr _b_286(.a(_w_405),.q(_w_406));
  bfr _b_285(.a(_w_404),.q(_w_405));
  bfr _b_282(.a(_w_401),.q(_w_402));
  bfr _b_281(.a(_w_400),.q(_w_401));
  bfr _b_279(.a(_w_398),.q(_w_390));
  bfr _b_278(.a(_w_397),.q(_w_398));
  bfr _b_277(.a(_w_396),.q(_w_397));
  bfr _b_272(.a(_w_391),.q(_w_392));
  bfr _b_269(.a(_w_388),.q(_w_389));
  bfr _b_268(.a(_w_387),.q(_w_388));
  bfr _b_267(.a(_w_386),.q(_w_387));
  bfr _b_264(.a(_w_383),.q(_w_384));
  bfr _b_327(.a(_w_446),.q(_w_447));
  bfr _b_261(.a(_w_380),.q(_w_381));
  bfr _b_260(.a(_w_379),.q(_w_380));
  bfr _b_323(.a(_w_442),.q(_w_443));
  bfr _b_259(.a(a_3_),.q(_w_379));
  bfr _b_258(.a(_w_377),.q(_w_375));
  bfr _b_257(.a(_w_376),.q(_w_377));
  spl2 a_1__s_0(.a(_w_374),.q0(a_1__0),.q1(a_1__1));
  or_bb g41(.a(n20_3),.b(n34_2),.q(n41));
  bfr _b_164(.a(_w_283),.q(_w_284));
  bfr _b_256(.a(a_2_),.q(_w_376));
  spl3L g23_s_3(.a(n23_6),.q0(n23_7),.q1(n23_8),.q2(_w_372));
  bfr _b_263(.a(a_4_),.q(_w_383));
  spl2 g23_s_1(.a(n23_0),.q0(n23_3),.q1(n23_4));
  spl3L b_2__s_0(.a(_w_412),.q0(b_2__0),.q1(b_2__1),.q2(_w_370));
  bfr _b_316(.a(_w_435),.q(_w_427));
  and_bb g73(.a(a_5__1),.b(b_5__2),.q(n73));
  bfr _b_242(.a(_w_361),.q(_w_362));
  bfr _b_328(.a(_w_447),.q(_w_436));
  bfr _b_225(.a(_w_344),.q(_w_345));
  bfr _b_139(.a(_w_258),.q(_w_259));
  bfr _b_173(.a(_w_292),.q(_w_293));
  spl2 g38_s_0(.a(n38),.q0(n38_0),.q1(n38_1));
  spl2 g68_s_0(.a(n68),.q0(n43_2),.q1(n68_1));
  maj_bbi g59(.a(n37_4),.b(n58),.c(n38_1),.q(_w_354));
  and_bb g52(.a(n49_0),.b(n51),.q(n52));
  spl3L g23_s_0(.a(n23),.q0(n23_0),.q1(n23_1),.q2(n23_2));
  maj_bbi g45(.a(b_4__5),.b(n44),.c(n23_2),.q(n45));
  spl4L g39_s_0(.a(n39),.q0(n39_0),.q1(n20_4),.q2(n39_2),.q3(_w_353));
  bfr _b_186(.a(_w_305),.q(_w_306));
  bfr _b_199(.a(_w_318),.q(_w_319));
  spl2 b_7__s_0(.a(b_7_),.q0(b_7__0),.q1(b_7__1));
  spl4L g20_s_1(.a(n20_1),.q0(n20_2),.q1(n20_3),.q2(n39_1),.q3(n20_5));
  bfr _b_191(.a(_w_310),.q(n25_1));
  spl4L g34_s_0(.a(n34),.q0(n34_0),.q1(n34_1),.q2(n34_2),.q3(n34_3));
  spl2 a_5__s_1(.a(a_5__2),.q0(a_5__3),.q1(_w_373));
  spl2 g24_s_1(.a(n24_0),.q0(n24_3),.q1(_w_350));
  spl4L g25_s_1(.a(n25_1),.q0(n25_2),.q1(n52_2),.q2(n25_4),.q3(_w_349));
  bfr _b_262(.a(_w_381),.q(_w_378));
  spl3L g52_s_0(.a(n52),.q0(n52_0),.q1(n53_1),.q2(n84_0));
  spl3L g28_s_0(.a(n28),.q0(n28_0),.q1(n28_1),.q2(_w_348));
  bfr _b_280(.a(a_6_),.q(_w_400));
  spl3L g22_s_2(.a(n22_3),.q0(n22_4),.q1(n22_5),.q2(_w_347));
  spl4L g42_s_0(.a(n42),.q0(n42_0),.q1(n28_3),.q2(n21_6),.q3(_w_346));
  spl2 g18_s_0(.a(n18),.q0(n18_0),.q1(_w_343));
  bfr _b_293(.a(b_2_),.q(_w_413));
  spl3L g24_s_0(.a(n24),.q0(n24_0),.q1(n24_1),.q2(n24_2));
  bfr _b_190(.a(n50),.q(_w_310));
  bfr _b_229(.a(n28_1),.q(n28_2));
  bfr _b_236(.a(_w_355),.q(_w_356));
  spl2 b_1__s_0(.a(_w_411),.q0(b_1__0),.q1(b_1__1));
  maj_bbi g44(.a(a_4__3),.b(_w_270),.c(_w_334),.q(n44));
  bfr _b_193(.a(_w_312),.q(_w_313));
  bfr _b_204(.a(_w_323),.q(a_4__3));
  spl2 g53_s_0(.a(n53),.q0(n53_0),.q1(_w_341));
  spl2 g74_s_0(.a(n74),.q0(n74_0),.q1(n46_2));
  bfr _b_239(.a(_w_358),.q(_w_359));
  spl2 g80_s_0(.a(n80),.q0(n49_2),.q1(n80_1));
  bfr _b_314(.a(_w_433),.q(_w_434));
  maj_bbb g21(.a(a_2__2),.b(b_2__2),.c(_w_330),.q(n21));
  maj_bbb g85(.a(n25_3),.b(n52_2),.c(n84_0),.q(n85));
  maj_bbi g83(.a(n24_7),.b(n82),.c(n81),.q(_w_338));
  spl2 b_6__s_1(.a(b_6__0),.q0(b_6__4),.q1(_w_337));
  bfr _b_159(.a(_w_278),.q(_w_279));
  spl3L g21_s_1(.a(n21_0),.q0(n21_2),.q1(n21_3),.q2(_w_336));
  maj_bbi g82(.a(n49_2),.b(_w_322),.c(n24_6),.q(n82));
  bfr _b_231(.a(n24_3),.q(n24_4));
  bfr _b_243(.a(_w_362),.q(_w_363));
  spl4L a_6__s_0(.a(_w_399),.q0(a_6__0),.q1(a_6__1),.q2(a_6__2),.q3(_w_335));
  spl2 b_4__s_1(.a(b_4__0),.q0(b_4__4),.q1(_w_334));
  bfr _b_273(.a(_w_392),.q(_w_393));
  bfr _b_219(.a(_w_338),.q(_w_339));
  maj_bbb g81(.a(n24_5),.b(n49_1),.c(n80_1),.q(n81));
  spl3L a_2__s_0(.a(_w_375),.q0(a_2__0),.q1(a_2__1),.q2(_w_333));
  bfr _b_136(.a(_w_255),.q(_w_256));
  spl2 g20_s_0(.a(n20),.q0(n20_0),.q1(_w_330));
  bfr _b_151(.a(n22_2),.q(n22_3));
  or_bb g78(.a(a_6__1),.b(b_6__2),.q(n78));
  bfr _b_237(.a(_w_356),.q(_w_357));
  maj_bbi g75(.a(n23_7),.b(n74_0),.c(n46_1),.q(n76));
  maj_bbi g71(.a(n22_6),.b(n70),.c(n69),.q(_w_324));
  bfr _b_297(.a(_w_416),.q(_w_417));
  bfr _b_208(.a(_w_327),.q(_w_328));
  maj_bbi g70(.a(n43_2),.b(n68_0),.c(_w_347),.q(n70));
  spl4L a_4__s_0(.a(_w_382),.q0(a_4__0),.q1(a_4__1),.q2(a_4__2),.q3(_w_323));
  maj_bbb g69(.a(n22_4),.b(n43_1),.c(n68_1),.q(n69));
  spl3L g49_s_0(.a(n49),.q0(n49_0),.q1(n49_1),.q2(n24_6));
  bfr _b_294(.a(_w_413),.q(_w_414));
  bfr _b_137(.a(_w_256),.q(s_3_));
  bfr _b_195(.a(_w_314),.q(_w_315));
  or_bb g66(.a(a_4__1),.b(b_4__2),.q(n66));
  spl3L g24_s_2(.a(n24_4),.q0(n24_5),.q1(n80_0),.q2(_w_322));
  maj_bbi g64(.a(n42_1),.b(n42_2),.c(n21_6),.q(n42_3));
  maj_bbi g62(.a(n60),.b(n61),.c(n39_3),.q(_w_311));
  and_bb g67(.a(a_4__2),.b(b_4__3),.q(n67));
  bfr _b_224(.a(n18_0),.q(_w_344));
  bfr _b_253(.a(_w_372),.q(n75));
  maj_bbi g61(.a(n34_0),.b(n39_2),.c(n20_5),.q(n39_3));
  bfr _b_201(.a(_w_320),.q(_w_321));
  spl3L b_0__s_0(.a(b_0_),.q0(b_0__0),.q1(b_0__1),.q2(b_0__2));
  bfr _b_198(.a(_w_317),.q(_w_318));
  or_bb g72(.a(a_5__0),.b(b_5__1),.q(n72));
  bfr _b_131(.a(_w_250),.q(_w_251));
  bfr _b_215(.a(b_4__4),.q(b_4__5));
  or_bb g55(.a(n18_1),.b(n54),.q(cout));
  maj_bbb g54(.a(n25_2),.b(n52_1),.c(n53_1),.q(n54));
  spl3L b_1__s_1(.a(b_1__1),.q0(b_1__2),.q1(b_1__3),.q2(n37_0));
  or_bb g53(.a(a_7__1),.b(b_7__1),.q(_w_296));
  bfr _b_142(.a(_w_261),.q(_w_262));
  maj_bbi g87(.a(n25_5),.b(n86),.c(n85),.q(s_7_));
  bfr _b_295(.a(_w_414),.q(_w_412));
  bfr _b_145(.a(_w_264),.q(_w_265));
  and_bi g80(.a(n78),.b(n79),.q(n80));
  and_bi g84(.a(n53_0),.b(_w_343),.q(n84));
  spl2 g22_s_0(.a(n22),.q0(n22_0),.q1(n22_1));
  maj_bbi g40(.a(n20_2),.b(n34_1),.c(_w_353),.q(n40));
  and_bb g49(.a(n46_0),.b(n48),.q(n49));
  bfr _b_251(.a(b_2__0),.q(b_2__2));
  maj_bbi g47(.a(a_5__4),.b(b_5__4),.c(n23_4),.q(n47));
  bfr _b_161(.a(_w_280),.q(_w_281));
  spl3L c_s_0(.a(c),.q0(c_0),.q1(c_1),.q2(_w_332));
  spl3L a_5__s_0(.a(_w_390),.q0(a_5__0),.q1(a_5__1),.q2(a_5__2));
  bfr _b_221(.a(a_0__4),.q(a_0__5));
  spl3L a_0__s_1(.a(a_0__2),.q0(a_0__3),.q1(a_0__4),.q2(_w_340));
  maj_bbi g77(.a(n75),.b(n76),.c(n23_9),.q(_w_292));
  and_bi g42(.a(n41),.b(n40),.q(n42));
  maj_bbb g25(.a(a_6__0),.b(b_6__1),.c(n24_1),.q(n25));
  maj_bbi g60(.a(n20_4),.b(n39_1),.c(n34_3),.q(n61));
  and_bi g34(.a(n32),.b(n33),.q(n34));
  bfr _b_308(.a(b_5_),.q(_w_428));
  bfr _b_153(.a(_w_272),.q(b_3__2));
  and_bi g39(.a(n38_0),.b(n36),.q(n39));
  spl3L b_5__s_0(.a(_w_427),.q0(b_5__0),.q1(b_5__1),.q2(b_5__2));
  spl2 g23_s_2(.a(n23_3),.q0(n23_5),.q1(n23_6));
  bfr _b_227(.a(n42_0),.q(n63));
  maj_bbb g38(.a(a_1__3),.b(_w_351),.c(n37_0),.q(n38));
  and_bb g46(.a(n43_0),.b(n45),.q(n46));
  maj_bbb g37(.a(a_0__1),.b(b_0__2),.c(_w_332),.q(n37));
  maj_bbi g76(.a(n23_8),.b(n46_2),.c(n74_1),.q(n23_9));
  bfr _b_148(.a(_w_267),.q(_w_268));
  bfr _b_217(.a(n21_3),.q(n21_4));
  maj_bbb g36(.a(a_1__0),.b(b_1__0),.c(n35),.q(_w_290));
  bfr _b_141(.a(_w_260),.q(_w_261));
  bfr _b_181(.a(_w_300),.q(_w_301));
  maj_bbi g35(.a(a_0__0),.b(b_0__1),.c(c_1),.q(n35));
  maj_bbi g57(.a(a_0__5),.b(n56),.c(n37_2),.q(_w_274));
  bfr _b_305(.a(_w_424),.q(_w_425));
  bfr _b_299(.a(_w_418),.q(_w_415));
  bfr _b_169(.a(_w_288),.q(_w_289));
  bfr _b_180(.a(_w_299),.q(_w_300));
  bfr _b_326(.a(_w_445),.q(_w_446));
  spl4L b_6__s_0(.a(_w_436),.q0(b_6__0),.q1(b_6__1),.q2(b_6__2),.q3(b_6__3));
  or_bb g31(.a(n29),.b(n30),.q(n31));
  and_bi g30(.a(n28_0),.b(_w_336),.q(n30));
  spl3L a_1__s_1(.a(a_1__1),.q0(a_1__2),.q1(_w_371),.q2(_w_351));
  spl2 g37_s_1(.a(n37_1),.q0(n37_3),.q1(_w_331));
  bfr _b_170(.a(_w_289),.q(s_0_));
  and_bi g29(.a(n21_2),.b(_w_348),.q(n29));
  bfr _b_133(.a(_w_252),.q(_w_253));
  and_bi g28(.a(n26),.b(n27),.q(n28));
  and_bb g27(.a(a_3__1),.b(_w_271),.q(n27));
  bfr _b_324(.a(_w_443),.q(_w_444));
  or_bb g26(.a(a_3__0),.b(b_3__1),.q(n26));
  bfr _b_275(.a(_w_394),.q(_w_395));
  maj_bbi g86(.a(n52_0),.b(n84_1),.c(_w_349),.q(n86));
  bfr _b_165(.a(_w_284),.q(_w_285));
  spl3L b_3__s_0(.a(_w_415),.q0(b_3__0),.q1(b_3__1),.q2(_w_271));
  maj_bbi g51(.a(b_6__5),.b(_w_309),.c(n25_0),.q(n51));
  spl2 g21_s_0(.a(n21),.q0(n21_0),.q1(n21_1));
  bfr _b_196(.a(_w_315),.q(_w_316));
  bfr _b_203(.a(n80_0),.q(n24_7));
  spl3L a_0__s_0(.a(a_0_),.q0(a_0__0),.q1(a_0__1),.q2(a_0__2));
  maj_bbb g24(.a(a_5__3),.b(_w_273),.c(n23_1),.q(n24));
  bfr _b_144(.a(_w_263),.q(_w_264));
  bfr _b_222(.a(_w_341),.q(_w_342));
  maj_bbb g23(.a(a_4__0),.b(b_4__1),.c(n22_1),.q(n23));
  spl2 g22_s_1(.a(n22_0),.q0(n22_2),.q1(_w_270));
  bfr _b_283(.a(_w_402),.q(_w_403));
  and_bi g68(.a(n66),.b(n67),.q(n68));
  bfr _b_245(.a(_w_364),.q(_w_365));
  bfr _b_266(.a(_w_385),.q(_w_386));
  spl2 g25_s_0(.a(n25),.q0(n50),.q1(_w_309));
  bfr _b_168(.a(_w_287),.q(_w_288));
  and_bb g43(.a(n31),.b(_w_346),.q(n43));
  maj_bbi g63(.a(n21_5),.b(n28_4),.c(n28_3),.q(n64));
  spl3L g37_s_0(.a(n37),.q0(a_1__3),.q1(n37_1),.q2(n37_2));
  bfr _b_246(.a(_w_365),.q(_w_366));
  maj_bbi g58(.a(a_1__4),.b(b_1__4),.c(_w_331),.q(n58));
  bfr _b_143(.a(_w_262),.q(_w_263));
  bfr _b_197(.a(_w_316),.q(_w_317));
  bfr _b_162(.a(_w_281),.q(_w_282));
  or_bb g32(.a(a_2__0),.b(b_2__1),.q(n32));
  and_bb g19(.a(a_0__3),.b(b_0__4),.q(n19));
  bfr _b_301(.a(_w_420),.q(_w_421));
  and_bb g33(.a(a_2__1),.b(_w_370),.q(n33));
  and_bb g18(.a(a_7__0),.b(b_7__0),.q(_w_257));
  spl2 b_0__s_1(.a(b_0__0),.q0(b_0__3),.q1(b_0__4));
  and_bb g79(.a(a_6__2),.b(b_6__3),.q(n79));
  bfr _b_130(.a(_w_249),.q(_w_250));
  spl2 g84_s_0(.a(n84),.q0(n25_3),.q1(n84_1));
  maj_bbb g20(.a(a_1__2),.b(b_1__3),.c(n19),.q(n20));
  spl2 g21_s_2(.a(n21_4),.q0(n21_5),.q1(n42_2));
  bfr _b_202(.a(_w_321),.q(s_2_));
  bfr _b_212(.a(n37_3),.q(n37_4));
  bfr _b_132(.a(_w_251),.q(_w_252));
  bfr _b_134(.a(_w_253),.q(_w_254));
  bfr _b_135(.a(_w_254),.q(_w_255));
  bfr _b_140(.a(_w_259),.q(_w_260));
  bfr _b_265(.a(_w_384),.q(_w_385));
  bfr _b_146(.a(_w_265),.q(_w_266));
  bfr _b_147(.a(_w_266),.q(_w_267));
  spl3L g46_s_0(.a(n46),.q0(n46_0),.q1(n46_1),.q2(n74_1));
  bfr _b_149(.a(_w_268),.q(_w_269));
  maj_bbi g50(.a(a_6__3),.b(_w_350),.c(_w_337),.q(n25_0));
  maj_bbi g65(.a(n63),.b(n64),.c(n42_3),.q(_w_249));
  bfr _b_216(.a(_w_335),.q(a_6__3));
  bfr _b_150(.a(_w_269),.q(n18));
  spl2 b_5__s_1(.a(b_5__0),.q0(b_5__3),.q1(_w_273));
  bfr _b_154(.a(b_5__3),.q(b_5__4));
  bfr _b_313(.a(_w_432),.q(_w_433));
  bfr _b_292(.a(b_1_),.q(_w_411));
  bfr _b_152(.a(b_3__0),.q(_w_272));
  bfr _b_172(.a(_w_291),.q(n36));
  bfr _b_155(.a(_w_274),.q(_w_275));
  bfr _b_156(.a(_w_275),.q(_w_276));
  bfr _b_138(.a(_w_257),.q(_w_258));
  bfr _b_157(.a(_w_276),.q(_w_277));
  spl3L g43_s_0(.a(n43),.q0(n43_0),.q1(n43_1),.q2(n68_0));
  bfr _b_187(.a(_w_306),.q(_w_307));
  bfr _b_207(.a(_w_326),.q(_w_327));
  bfr _b_158(.a(_w_277),.q(_w_278));
  maj_bbi g48(.a(n23_5),.b(n47),.c(n24_2),.q(n48));
  bfr _b_163(.a(_w_282),.q(_w_283));
  bfr _b_166(.a(_w_285),.q(_w_286));
  bfr _b_174(.a(_w_293),.q(_w_294));
  bfr _b_271(.a(a_5_),.q(_w_391));
  bfr _b_179(.a(_w_298),.q(_w_299));
  bfr _b_175(.a(_w_294),.q(_w_295));
  bfr _b_255(.a(a_1_),.q(_w_374));
  bfr _b_176(.a(_w_295),.q(s_5_));
  bfr _b_177(.a(_w_296),.q(_w_297));
  bfr _b_250(.a(_w_369),.q(a_3__2));
  bfr _b_320(.a(_w_439),.q(_w_440));
  bfr _b_182(.a(_w_301),.q(_w_302));
  bfr _b_183(.a(_w_302),.q(_w_303));
  bfr _b_184(.a(_w_303),.q(_w_304));
  bfr _b_185(.a(_w_304),.q(_w_305));
  bfr _b_310(.a(_w_429),.q(_w_430));
  bfr _b_238(.a(_w_357),.q(_w_358));
  bfr _b_188(.a(_w_307),.q(_w_308));
  bfr _b_178(.a(_w_297),.q(_w_298));
  bfr _b_189(.a(_w_308),.q(n53));
  and_bi g74(.a(n72),.b(n73),.q(_w_352));
  bfr _b_192(.a(_w_311),.q(_w_312));
  bfr _b_171(.a(_w_290),.q(_w_291));
  bfr _b_194(.a(_w_313),.q(_w_314));
  spl4L b_4__s_0(.a(_w_419),.q0(b_4__0),.q1(b_4__1),.q2(b_4__2),.q3(b_4__3));
  bfr _b_200(.a(_w_319),.q(_w_320));
  bfr _b_235(.a(_w_354),.q(_w_355));
  bfr _b_167(.a(_w_286),.q(_w_287));
  bfr _b_205(.a(_w_324),.q(_w_325));
  bfr _b_206(.a(_w_325),.q(_w_326));
  bfr _b_270(.a(_w_389),.q(_w_382));
  spl2 g28_s_1(.a(n28_2),.q0(n42_1),.q1(n28_4));
  maj_bbb g22(.a(a_3__2),.b(b_3__2),.c(n21_1),.q(n22));
  bfr _b_160(.a(_w_279),.q(_w_280));
  bfr _b_210(.a(_w_329),.q(s_4_));
  bfr _b_211(.a(n20_0),.q(n20_1));
  bfr _b_306(.a(_w_425),.q(_w_426));
  bfr _b_213(.a(c_0),.q(c_2));
  bfr _b_276(.a(_w_395),.q(_w_396));
  bfr _b_214(.a(_w_333),.q(a_2__2));
  bfr _b_218(.a(b_6__4),.q(b_6__5));
  spl2 a_7__s_0(.a(a_7_),.q0(a_7__0),.q1(a_7__1));
  bfr _b_220(.a(_w_339),.q(s_6_));
  bfr _b_230(.a(n25_4),.q(n25_5));
  bfr _b_241(.a(_w_360),.q(_w_361));
  bfr _b_226(.a(_w_345),.q(n18_1));
  bfr _b_247(.a(_w_366),.q(_w_367));
  maj_bbi g56(.a(b_0__3),.b(c_2),.c(_w_340),.q(n56));
  bfr _b_228(.a(n22_5),.q(n22_6));
  bfr _b_232(.a(_w_371),.q(a_1__4));
  bfr _b_233(.a(_w_352),.q(n74));
  bfr _b_318(.a(_w_437),.q(_w_438));
  bfr _b_234(.a(n39_0),.q(n60));
  bfr _b_240(.a(_w_359),.q(_w_360));
  bfr _b_244(.a(_w_363),.q(_w_364));
  bfr _b_223(.a(_w_342),.q(n52_1));
  bfr _b_249(.a(_w_368),.q(_w_369));
  bfr _b_284(.a(_w_403),.q(_w_404));
  bfr _b_248(.a(_w_367),.q(s_1_));
  bfr _b_274(.a(_w_393),.q(_w_394));
  spl3L a_3__s_0(.a(_w_378),.q0(a_3__0),.q1(a_3__1),.q2(_w_368));
  bfr _b_209(.a(_w_328),.q(_w_329));
  bfr _b_252(.a(b_1__2),.q(b_1__4));
  bfr _b_303(.a(_w_422),.q(_w_423));
  bfr _b_254(.a(_w_373),.q(a_5__4));
endmodule
