module c499 (N1,N101,N105,N109,N113,N117,N121,N125,N129,N13,N130,N131,N132,N133,N134,N135,N136,N137,N17,N21,N25,N29,N33,N37,N41,N45,N49,N5,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N9,N93,N97,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755);
  input N1,N101,N105,N109,N113,N117,N121,N125,N129,N13,N130,N131,N132,N133,N134,N135,N136,N137,N17,N21,N25,N29,N33,N37,N41,N45,N49,N5,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N9,N93,N97;
  output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755;
  wire _w_1977,_w_1975,_w_1973,_w_1970,_w_1967,_w_1965,_w_1964,_w_1960,_w_1959,_w_1952,_w_1951,_w_1948,_w_1946,_w_1941,_w_1971,_w_1939,_w_1936,_w_1934,_w_1933,_w_1956,_w_1929,_w_1925,_w_1924,_w_1923,_w_1921,_w_1919,_w_1917,_w_1915,_w_1913,_w_1909,_w_1906,_w_1904,_w_1903,_w_1902,_w_1899,_w_1898,_w_1897,_w_1895,_w_1888,_w_1886,_w_1885,_w_1883,_w_1882,_w_1881,_w_1880,_w_1879,_w_1877,_w_1875,_w_1874,_w_1872,_w_1920,_w_1870,_w_1869,_w_1867,_w_1865,_w_1914,_w_1863,_w_1862,_w_1861,_w_1859,_w_1858,_w_1852,_w_1851,_w_1850,_w_1849,_w_1848,_w_1846,_w_1845,_w_1844,_w_1842,_w_1841,_w_1840,_w_1838,_w_1836,_w_1828,_w_1827,_w_1826,_w_1825,_w_1824,_w_1820,_w_1819,_w_1818,_w_1811,_w_1808,_w_1804,_w_1835,_w_1803,_w_1802,_w_1801,_w_1795,_w_1794,_w_1793,_w_1792,_w_1790,_w_1789,_w_1787,_w_1785,_w_1873,_w_1853,_w_1784,_w_1783,_w_1782,_w_1777,_w_1776,_w_1775,_w_1774,_w_1772,_w_1771,_w_1770,_w_1768,_w_1766,_w_1763,_w_1762,_w_1760,_w_1759,_w_1758,_w_1757,_w_1752,_w_1747,_w_1963,_w_1745,_w_1737,_w_1893,_w_1733,_w_1725,_w_1722,_w_1721,_w_1720,_w_1719,_w_1717,_w_1716,_w_1812,_w_1712,_w_1711,_w_1707,_w_1702,_w_1701,_w_1698,_w_1966,_w_1697,_w_1696,_w_1695,_w_1694,_w_1691,_w_1687,_w_1686,_w_1685,_w_1681,_w_1680,_w_1676,_w_1670,_w_1668,_w_1666,_w_1665,_w_1660,_w_1657,_w_1655,_w_1654,_w_1652,_w_1651,_w_1647,_w_1644,_w_1643,_w_1639,_w_1637,_w_1634,_w_1633,_w_1630,_w_1626,_w_1624,_w_1621,_w_1620,_w_1618,_w_1614,_w_1613,_w_1612,_w_1627,_w_1610,_w_1609,_w_1607,_w_1606,_w_1605,_w_1604,_w_1603,_w_1602,_w_1601,_w_1599,_w_1595,_w_1592,_w_1590,_w_1589,_w_1976,_w_1588,_w_1927,_w_1587,_w_1833,_w_1584,_w_1582,_w_1581,_w_1580,_w_1837,_w_1576,_w_1574,_w_1572,_w_1571,_w_1570,_w_1569,_w_1568,_w_1567,_w_1565,_w_1645,_w_1563,_w_1559,_w_1558,_w_1557,_w_1556,_w_1552,_w_1551,_w_1550,_w_1548,_w_1542,_w_1541,_w_1539,_w_1538,_w_1536,_w_1535,_w_1534,_w_1544,_w_1533,_w_1530,_w_1529,_w_1528,_w_1683,_w_1526,_w_1520,_w_1519,_w_1798,_w_1516,_w_1640,_w_1512,_w_1511,_w_1510,_w_1507,_w_1505,_w_1504,_w_1503,_w_1502,_w_1501,_w_1692,_w_1500,_w_1499,_w_1497,_w_1495,_w_1494,_w_1492,_w_1491,_w_1490,_w_1489,_w_1488,_w_1806,_w_1486,_w_1484,_w_1482,_w_1481,_w_1809,_w_1479,_w_1478,_w_1477,_w_1476,_w_1474,_w_1470,_w_1469,_w_1467,_w_1600,_w_1466,_w_1464,_w_1463,_w_1461,_w_1458,_w_1457,_w_1456,_w_1455,_w_1451,_w_1447,_w_1445,_w_1444,_w_1855,_w_1443,_w_1442,_w_1441,_w_1440,_w_1439,_w_1434,_w_1431,_w_1427,_w_1424,_w_1421,_w_1496,_w_1420,_w_1656,_w_1419,_w_1415,_w_1414,_w_1413,_w_1754,_w_1732,_w_1437,_w_1412,_w_1411,_w_1406,_w_1405,_w_1404,_w_1402,_w_1401,_w_1400,_w_1398,_w_1395,_w_1393,_w_1616,_w_1392,_w_1515,_w_1391,_w_1388,_w_1387,_w_1974,_w_1386,_w_1383,_w_1547,_w_1381,_w_1564,_w_1380,_w_1379,_w_1678,_w_1376,_w_1375,_w_1374,_w_1373,_w_1371,_w_1705,_w_1454,_w_1370,_w_1369,_w_1713,_w_1368,_w_1947,_w_1366,_w_1365,_w_1364,_w_1363,_w_1950,_w_1362,_w_1360,_w_1356,_w_1354,_w_1677,_w_1353,_w_1350,_w_1348,_w_1736,_w_1347,_w_1345,_w_1343,_w_1342,_w_1807,_w_1337,_w_1336,_w_1335,_w_1334,_w_1598,_w_1344,_w_1333,_w_1331,_w_1330,_w_1699,_w_1329,_w_1327,_w_1325,_w_1324,_w_1323,_w_1322,_w_1321,_w_1320,_w_1319,_w_1318,_w_1317,_w_1937,_w_1315,_w_1312,_w_1311,_w_1310,_w_1813,_w_1540,_w_1309,_w_1308,_w_1307,_w_1306,_w_1303,_w_1301,_w_1300,_w_1299,_w_1296,_w_1295,_w_1689,_w_1294,_w_1293,_w_1292,_w_1290,_w_1288,_w_1546,_w_1287,_w_1521,_w_1286,_w_1282,_w_1619,_w_1281,_w_1955,_w_1280,_w_1277,_w_1275,_w_1796,_w_1274,_w_1662,_w_1273,_w_1272,_w_1709,_w_1271,_w_1485,_w_1270,_w_1708,_w_1269,_w_1468,_w_1267,_w_1263,_w_1748,_w_1262,_w_1261,_w_1259,_w_1688,_w_1257,_w_1255,_w_1253,_w_1459,_w_1251,_w_1250,_w_1244,_w_1241,_w_1240,_w_1237,_w_1487,_w_1236,_w_1235,_w_1596,_w_1233,_w_1232,_w_1231,_w_1230,_w_1227,_w_1225,_w_1224,_w_1222,_w_1428,_w_1221,_w_1409,_w_1243,_w_1220,_w_1480,_w_1217,_w_1900,_w_1735,_w_1215,_w_1214,_w_1212,_w_1211,_w_1210,_w_1209,_w_1206,_w_1204,_w_1203,_w_1734,_w_1352,_w_1202,_w_1200,_w_1197,_w_1196,_w_1585,_w_1194,_w_1191,_w_1817,_w_1187,_w_1186,_w_1185,_w_1432,_w_1184,_w_1219,_w_1183,_w_1182,_w_1180,_w_1179,_w_1177,_w_1176,_w_1175,_w_1174,_w_1173,_w_1171,_w_1170,_w_1901,_w_1767,_w_1509,_w_1169,_w_1168,_w_1664,_w_1166,_w_1396,_w_1163,_w_1161,_w_1160,_w_1159,_w_1483,_w_1158,_w_1156,_w_1246,_w_1155,_w_1153,_w_1152,_w_1864,_w_1151,_w_1617,_w_1146,_w_1144,_w_1788,_w_1143,_w_1890,_w_1141,_w_1140,_w_1139,_w_1138,_w_1137,_w_1132,_w_1131,_w_1129,_w_1127,_w_1126,_w_1125,_w_1124,_w_1123,_w_1122,_w_1121,_w_1753,_w_1119,_w_1117,_w_1116,_w_1961,_w_1435,_w_1113,_w_1112,_w_1111,_w_1663,_w_1109,n215_1,_w_1816,n253_0,_w_1659,n142,n259_8,_w_1378,n259_7,n259_3,n78_6,_w_1868,_w_1410,n262_1,n148,n137_2,n317_0,n132,n196,n266_1,n144,n269_1,n96,N13_0,_w_1871,N121_1,n278_7,n278_1,n282_1,_w_1843,n294_1,N33_0,n298_0,n42,_w_1942,_w_1473,n304_1,n61,_w_1672,n308_0,n100_2,n358_1,n358_0,n413_0,_w_1710,n259_6,n318_3,_w_1894,_w_1475,_w_1417,n318_0,n335_2,n336_1,n336_0,_w_1912,n281_3,n360_2,n55,n112_1,n379_0,_w_1943,n232,n383_1,n383_0,n395_3,_w_1797,n152_3,n270,n308_1,_w_1653,n395_0,_w_1918,n290,n413_1,n286,n421_0,_w_1256,n275_0,_w_1265,n204,_w_1114,n426,n89,n184_1,n413,_w_1372,_w_1223,n379_1,n406,n316_0,n401,n400,N17_4,n397,_w_1399,N109_2,n340_1,n290_0,_w_1690,n395,_w_1446,n209_4,n391,_w_1646,_w_1149,n389,_w_1276,N37_6,_w_1706,n383,_w_1426,n177,n381,n379,n78,n100,_w_1856,n418,_w_1714,n266,n370,_w_1693,_w_1560,_w_1527,n366,n345,n365,_w_1349,_w_1284,n153_1,_w_1545,n360,n359,n207,n91_1,n357,n356,N109_3,n54_1,N113_1,n422,n348,_w_1377,N45_3,n369,_w_1823,N73_2,_w_1130,n346,n67,_w_1118,n45_1,_w_1433,N101_3,n272_1,n337,n233_3,_w_1147,n44_1,n335,n332,n281_2,n146,N53_7,n244_1,n152_0,n181_4,n328,_w_1096,n327,n209_7,n402,N113_0,n208,_w_1264,n344_0,_w_1761,_w_1493,n79_1,n320,N41_0,_w_1969,n194,N121_4,_w_1506,n278_3,n318,n387,n358,n316,n51,N13_1,n306,n304,n199,N61_5,n341,n301,n66_0,n300,n209_8,n414,n109,n278,n233,_w_1635,n296,n209_2,n371,n292,N85_7,N81_4,n284,n226,n109_3,n269_0,n304_0,n138,N137_3,n283,n268,n282,n281,n280,_w_1723,n302,n182,n327_0,_w_1148,n276,_w_1549,n274,_w_1341,n273,_w_1649,N17_0,n272,n269,n421,n265,_w_1108,n263,n262,n425,n348_1,n221,N117_5,_w_1543,N49_5,n261,_w_1133,n60_0,_w_1834,n259,n215,n194_1,n160_1,_w_1916,n233_0,n257,_w_1932,n91,N21_2,n254,_w_1905,n250,n417_1,_w_1891,n114,N13_4,n224_0,N97_4,n92,n355,n247,_w_1738,n410,N105_7,N17_3,_w_1671,n300_0,_w_1554,n246,N121_2,n244,n128_1,n342,n380,n97_0,_w_1593,n278_0,_w_1724,n323_1,_w_1756,n181_0,n236,N17_5,n240_1,_w_1523,n230,n375,n227,n253_1,n417,_w_1839,N121_6,n153,n93,N113_2,n163_0,n350,n250_1,n291,n86,n70,_w_1907,n65,N5_6,n128_0,n425_0,n275,n412_3,n64,_w_1145,n361,n147,_w_1884,n313,n51_0,_w_1105,n319_1,n263_1,_w_1928,_w_1730,_w_1193,n185_0,N53_2,N25_6,n290_1,n331,_w_1531,n146_3,n340,N33_4,_w_1266,n255,n374,n278_5,_w_1358,n294,n218,_w_1814,_w_1658,n421_1,n134_1,n176,_w_1525,n210,n57,_w_1164,n323,n181_3,n195,n233_5,n335_0,_w_1650,n404,n280_0,n384,n151,N85_2,n53,n280_1,n278_2,_w_1195,N29_3,n79,n264,_w_1436,n52,_w_1968,n152_8,n395_2,n83,_w_1154,n310,n239,_w_1188,_w_1092,_w_1667,_w_1422,n282_0,n321,n249,n50,n221_0,n259_0,n278_8,n312,_w_1764,n47,n74,n169,n298_1,n316_1,N37_1,_w_1095,n82,N1_5,_w_1847,_w_1258,n43,n396_0,n45,n90,_w_1896,_w_1192,n113,n106,n181_6,n194_0,N33_5,N65_5,n278_4,n185_1,_w_1260,n305,_w_1382,n408_0,n54,N49_2,_w_1128,n295,n106_0,n238,_w_1462,n245,n247_1,N41_2,_w_1661,_w_1429,_w_1298,_w_1162,n281_1,n156,_w_1167,n188_1,n369_1,n125_0,_w_1190,n209_6,n122,_w_1213,_w_1460,n336,n209_5,n335_3,N25_3,_w_1810,n169_0,_w_1448,N65_4,n111,N77_5,_w_1586,n263_0,n56,_w_1239,n251,n71,_w_1110,_w_1779,n235_0,_w_1450,n253,n63_2,n191,_w_1471,n45_0,n60,_w_1743,n218_1,_w_1854,n166_1,n340_0,n127,_w_1234,n256,_w_1099,n198,n362,N65_1,n75,_w_1566,n131,N1_4,_w_1780,n388,n172,n131_1,_w_1135,n139,n211_0,n423,N65_6,n68,_w_1518,_w_1648,_w_1438,N57_3,_w_1791,N105_0,_w_1718,n247_0,_w_1632,_w_1181,n360_3,n143_1,_w_1889,n165,N17_7,n385,n367,n58,n412,_w_1328,n240,N77_1,n84,N25_1,_w_1751,_w_1165,_w_1597,n163,n105,_w_1623,n218_0,_w_1248,_w_1727,N93_3,n209_3,_w_1316,n327_1,n164,n69,n143,_w_1061,n308,n46,_w_1314,n48,_w_1778,n277,n76,_w_1561,_w_1684,n143_0,N9_1,n59,n181_5,n299,_w_1304,n211,n192,n88_0,n87,_w_1384,n85,n335_1,n107,n317,n279_0,N9_2,_w_1346,N29_0,n365_0,n160,n81,N105_5,n248,n216,n136,n344,n78_1,n161,N81_7,_w_1822,n235,N97_6,n409,N13_7,n408_1,n94,n117,_w_1769,n197,n124,n314,N117_2,n66,n97,n417_0,n344_1,n360_1,N97_2,_w_1953,n63_0,n425_1,_w_1931,n186,N137_1,n377,n187,N25_0,n112,n242,N137_6,n278_6,n391_1,n281_0,n119,n317_1,n120,n223,N41_1,_w_1673,N25_7,n123,_w_1359,n149,_w_1962,N89_0,n352,n126,_w_1205,_w_1198,n128,n125,_w_1085,n130,n175,N137_7,n224,n82_0,_w_1524,n213_0,n134,n190,n135,n200_1,_w_1498,_w_1103,n118,n235_1,n259_2,_w_1514,n267,n168,_w_1728,n137,n288,n158,n104,n141,_w_1742,_w_1098,_w_1831,_w_1522,n395_1,n205,n79_0,_w_1815,_w_1403,_w_1207,n419,n181_9,_w_1517,_w_1408,n63,_w_1591,_w_1508,n202,n210_1,n298_2,n150,_w_1750,n266_0,n309,N29_5,n110,n333,_w_1397,n152,n243,n359_0,_w_1578,n349,n360_0,n170,_w_1302,n206_0,n154,n178,n157,_w_1741,n184,n396,_w_1385,n193,n75_1,n159,_w_1326,_w_1189,n185,_w_1268,n214,n324,n318_1,n62,n369_0,n162,n60_1,n392,n166,_w_1805,n427,N5_2,_w_1555,_w_1537,N109_7,_w_1060,n167,n98,n387_1,_w_1430,_w_1339,_w_1313,n354,n171,n312_0,_w_1449,n287,_w_1065,n179,n155,n180,_w_1178,n181,_w_1892,n183,N97_7,N25_2,N109_0,n300_1,N37_5,n188,N137_0,n400_0,n200,_w_1978,_w_1746,n222,_w_1944,n189,n44,n129,n373,n201,n181_8,n203,_w_1615,_w_1107,n348_0,n115,n209,n353,N17_1,n212,n88,N49_4,n213,n230_1,N33_7,N93_4,n174,n78_4,n217,n365_1,n219,n220,n225,n299_0,n244_0,n243_0,n97_1,n243_1,_w_1799,N125_7,n230_0,n231,n85_1,n203_0,n227_0,n227_1,n78_0,n78_3,N85_5,n78_5,N85_1,n63_3,n78_7,_w_1091,n78_8,n91_0,_w_1669,n259_4,n169_1,n361_0,n361_1,n210_0,n57_0,n57_1,_w_1945,n94_1,_w_1423,n286_1,_w_1226,n258,N17_6,_w_1821,_w_1453,n77,n404_0,N101_6,n404_1,_w_1765,n94_0,_w_1573,n294_0,N121_7,n233_1,n331_0,n298_3,n233_4,n134_0,n49,n233_6,N117_7,_w_1332,N41_6,n233_7,n240_0,_w_1641,n233_8,n233_11,N97_1,_w_1305,n119_0,N97_3,n318_2,n101,N97_5,N57_0,_w_1860,n78_2,N57_1,n286_0,N77_4,n100_3,N57_2,N57_4,N57_5,N57_6,n109_1,N57_7,n323_0,n72_0,_w_1715,_w_1070,_w_1575,N81_0,N101_4,N81_1,n213_1,_w_1418,n197_0,N81_3,N81_5,N21_3,N81_6,n396_1,_w_1781,n82_1,n54_0,N41_4,n373_0,_w_1800,N41_7,n221_1,n378_0,N61_7,n119_1,_w_1216,_w_1115,n378_2,n378_3,n122_0,n122_1,_w_1208,n116_1,n73,N117_0,N117_1,_w_1622,n393,N117_3,N117_4,_w_1636,_w_1252,N117_6,_w_1247,n125_1,_w_1625,n259_1,N73_1,n140_1,N17_2,n191_0,n191_1,_w_1830,n209_1,n233_9,n146_0,n146_1,_w_1228,n146_2,_w_1452,n75_0,n271,n172_0,n172_1,_w_1297,N85_4,N1_3,_w_1629,N9_0,N53_6,N9_3,_w_1064,N9_4,_w_1355,N9_5,_w_1954,N5_1,n133,N9_6,N9_7,N89_1,N25_4,_w_1949,_w_1150,N89_2,_w_1254,N89_3,N13_5,N89_4,N89_5,N89_6,N89_7,n229,N33_2,_w_1157,N69_0,N69_1,N69_2,N69_3,N69_4,N69_6,_w_1513,n72_2,N69_7,_w_1367,N77_0,n241,N77_2,N77_3,_w_1957,n275_1,N77_6,_w_1704,N73_0,N73_3,n203_2,n319,N73_5,_w_1908,n72_3,N1_1,_w_1425,N73_7,_w_1910,_w_1201,n250_0,n363,n412_0,n272_0,n72,n412_1,_w_1278,_w_1172,_w_1071,n412_2,N61_0,_w_1700,n233_2,N61_1,N61_2,N61_3,N61_4,N61_6,N5_0,n181_1,N5_3,N5_4,N5_5,N5_7,n103,N49_0,_w_1357,n298,N49_1,N49_3,_w_1579,n319_0,N49_6,N49_7,N45_1,_w_1242,N45_2,_w_1390,N45_4,_w_1101,N45_5,N101_2,N45_6,N45_7,_w_1389,N109_1,N105_2,n163_1,N37_0,n206_1,n378,N37_2,N37_4,n387_0,n299_2,n102,N33_1,N1_2,n69_0,_w_1074,N33_3,_w_1749,N33_6,N29_1,n338,N29_2,n312_1,n184_0,N29_4,N73_6,N29_6,N29_7,_w_1887,_w_1829,N105_1,N21_0,N109_5,N21_1,n329,N21_4,n121,_w_1097,_w_1283,N21_5,N21_6,N21_7,n48_0,n48_1,_w_1338,n140,N53_0,_w_1740,_w_1079,N85_0,N85_6,N137_2,_w_1407,N109_6,N137_4,n145,N137_5,N137_8,N93_0,_w_1351,N137_9,n408,n299_1,_w_1674,N101_1,_w_1611,n115_4,n299_3,n69_1,n103_0,_w_1631,_w_1142,_w_1078,_w_1077,n103_1,n157_1,n85_0,_w_1832,_w_1638,N69_5,N53_4,_w_1291,n331_1,N93_1,N93_2,_w_1134,N13_3,N77_7,N93_5,N93_6,N93_7,_w_1930,_w_1628,_w_1465,n405,N13_2,N121_0,_w_1340,_w_1249,n233_10,n152_6,N121_3,N121_5,_w_1229,N41_3,N113_3,N113_4,_w_1394,n203_1,N113_5,_w_1938,_w_1726,N113_6,_w_1102,N113_7,N65_0,n325,N109_4,n400_1,n116,N1_0,n106_1,_w_1594,_w_1245,N45_0,n100_0,N73_4,N1_6,_w_1289,n66_1,N1_7,N105_3,n378_1,n181_2,_w_1731,N105_4,n99,N105_6,_w_1911,_w_1786,N125_5,_w_1120,n256_0,N101_0,N101_5,n175_2,N101_7,_w_1773,_w_1729,n109_0,_w_1532,n115_3,n109_2,n377_0,n112_0,n116_0,_w_1940,n197_1,n175_0,_w_1199,n391_0,n154_0,n175_1,_w_1583,n359_1,n175_3,n279,N53_1,n377_1,n51_1,N53_3,N53_5,_w_1703,n224_1,N25_5,N85_3,n137_1,_w_1935,n137_3,_w_1675,n100_1,N37_3,n140_0,_w_1922,_w_1878,_w_1136,n63_1,n237,n149_0,_w_1739,n149_1,n152_1,n173,n131_0,n152_2,_w_1069,n152_4,n152_5,_w_1279,n152_7,n153_0,_w_1472,n153_2,n72_1,n153_3,n154_1,_w_1577,n228,n80,N65_2,N65_3,_w_1876,_w_1755,N97_0,N65_7,n157_0,n160_0,_w_1682,_w_1084,n166_0,N125_0,n215_0,N125_1,n256_1,_w_1416,n373_1,N125_2,N125_3,N125_6,_w_1958,n178_0,_w_1361,n178_1,_w_1562,n181_7,n137_0,n188_0,n200_0,_w_1972,n44_0,n203_3,_w_1744,n115_0,_w_1238,n115_1,_w_1642,n115_2,n115_5,n234,n115_6,n115_7,_w_1553,n415,n115_8,_w_1285,n279_1,n209_0,n262_0,n212_0,n252,N81_2,n212_1,N13_6,n88_1,n108,_w_1062,_w_1866,_w_1608,_w_1063,_w_1066,_w_1679,_w_1067,_w_1068,_w_1072,_w_1926,_w_1073,_w_1075,_w_1076,_w_1080,_w_1081,_w_1857,N125_4,_w_1082,_w_1218,_w_1083,n95,n398,_w_1086,_w_1087,_w_1088,n259_5,N41_5,_w_1089,n260,_w_1090,_w_1093,n206,N37_7,_w_1094,n211_1,_w_1100,_w_1104,_w_1106;

  bfr _b_1559(.a(N53),.q(_w_1978));
  bfr _b_1556(.a(N33),.q(_w_1975));
  bfr _b_1555(.a(_w_1974),.q(_w_1973));
  bfr _b_1554(.a(N136),.q(_w_1974));
  bfr _b_1553(.a(_w_1972),.q(_w_1971));
  bfr _b_1551(.a(N134),.q(_w_1970));
  bfr _b_1550(.a(_w_1969),.q(_w_1968));
  bfr _b_1546(.a(_w_1965),.q(_w_1964));
  bfr _b_1544(.a(_w_1963),.q(_w_1962));
  bfr _b_1542(.a(N129),.q(_w_1961));
  bfr _b_1539(.a(_w_1958),.q(_w_1959));
  bfr _b_1537(.a(_w_1956),.q(_w_1957));
  bfr _b_1536(.a(_w_1955),.q(_w_1956));
  bfr _b_1535(.a(_w_1954),.q(_w_1955));
  bfr _b_1534(.a(_w_1953),.q(_w_1954));
  bfr _b_1533(.a(_w_1952),.q(_w_1953));
  bfr _b_1541(.a(_w_1960),.q(N105_5));
  bfr _b_1528(.a(_w_1947),.q(_w_1948));
  bfr _b_1526(.a(_w_1945),.q(_w_1946));
  bfr _b_1524(.a(_w_1943),.q(_w_1944));
  bfr _b_1523(.a(_w_1942),.q(_w_1943));
  bfr _b_1522(.a(_w_1941),.q(_w_1942));
  bfr _b_1521(.a(_w_1940),.q(_w_1941));
  bfr _b_1520(.a(_w_1939),.q(_w_1940));
  bfr _b_1519(.a(_w_1938),.q(_w_1939));
  bfr _b_1516(.a(_w_1935),.q(_w_1936));
  bfr _b_1515(.a(_w_1934),.q(_w_1935));
  bfr _b_1513(.a(_w_1932),.q(_w_1933));
  bfr _b_1512(.a(_w_1931),.q(_w_1932));
  bfr _b_1510(.a(_w_1929),.q(_w_1930));
  bfr _b_1509(.a(_w_1928),.q(_w_1929));
  bfr _b_1507(.a(_w_1926),.q(_w_1927));
  bfr _b_1506(.a(_w_1925),.q(_w_1926));
  bfr _b_1504(.a(_w_1923),.q(_w_1924));
  bfr _b_1503(.a(_w_1922),.q(_w_1923));
  bfr _b_1502(.a(_w_1921),.q(_w_1922));
  bfr _b_1500(.a(_w_1919),.q(_w_1920));
  bfr _b_1499(.a(_w_1918),.q(_w_1919));
  bfr _b_1497(.a(_w_1916),.q(_w_1917));
  bfr _b_1496(.a(_w_1915),.q(_w_1916));
  bfr _b_1493(.a(_w_1912),.q(_w_1913));
  bfr _b_1491(.a(_w_1910),.q(_w_1911));
  bfr _b_1489(.a(_w_1908),.q(_w_1909));
  bfr _b_1480(.a(_w_1899),.q(_w_1900));
  bfr _b_1475(.a(_w_1894),.q(_w_1895));
  bfr _b_1474(.a(_w_1893),.q(_w_1894));
  bfr _b_1473(.a(_w_1892),.q(_w_1893));
  bfr _b_1472(.a(_w_1891),.q(_w_1892));
  bfr _b_1471(.a(_w_1890),.q(N89_5));
  bfr _b_1470(.a(_w_1889),.q(_w_1890));
  bfr _b_1468(.a(_w_1887),.q(_w_1888));
  bfr _b_1466(.a(_w_1885),.q(_w_1886));
  bfr _b_1465(.a(_w_1884),.q(_w_1885));
  bfr _b_1463(.a(_w_1882),.q(_w_1883));
  bfr _b_1462(.a(_w_1881),.q(_w_1882));
  bfr _b_1459(.a(_w_1878),.q(_w_1879));
  bfr _b_1458(.a(_w_1877),.q(_w_1878));
  bfr _b_1456(.a(_w_1875),.q(_w_1876));
  bfr _b_1455(.a(_w_1874),.q(_w_1875));
  bfr _b_1454(.a(_w_1873),.q(_w_1874));
  bfr _b_1453(.a(_w_1872),.q(_w_1873));
  bfr _b_1450(.a(_w_1869),.q(_w_1870));
  bfr _b_1449(.a(_w_1868),.q(_w_1869));
  bfr _b_1444(.a(_w_1863),.q(_w_1864));
  bfr _b_1442(.a(_w_1861),.q(_w_1862));
  bfr _b_1461(.a(_w_1880),.q(_w_1881));
  bfr _b_1441(.a(_w_1860),.q(_w_1861));
  bfr _b_1440(.a(_w_1859),.q(_w_1860));
  bfr _b_1433(.a(_w_1852),.q(_w_1853));
  bfr _b_1431(.a(_w_1850),.q(_w_1851));
  bfr _b_1429(.a(_w_1848),.q(_w_1849));
  bfr _b_1427(.a(_w_1846),.q(_w_1847));
  bfr _b_1548(.a(_w_1967),.q(_w_1966));
  bfr _b_1424(.a(_w_1843),.q(N17_5));
  bfr _b_1422(.a(_w_1841),.q(_w_1842));
  bfr _b_1420(.a(_w_1839),.q(_w_1840));
  bfr _b_1419(.a(_w_1838),.q(_w_1839));
  bfr _b_1418(.a(_w_1837),.q(_w_1838));
  bfr _b_1417(.a(_w_1836),.q(_w_1837));
  bfr _b_1412(.a(_w_1831),.q(_w_1832));
  bfr _b_1410(.a(_w_1829),.q(_w_1830));
  bfr _b_1408(.a(_w_1827),.q(_w_1828));
  bfr _b_1407(.a(_w_1826),.q(_w_1827));
  bfr _b_1406(.a(_w_1825),.q(_w_1826));
  bfr _b_1405(.a(_w_1824),.q(_w_1825));
  bfr _b_1404(.a(_w_1823),.q(_w_1824));
  bfr _b_1403(.a(_w_1822),.q(_w_1823));
  bfr _b_1402(.a(_w_1821),.q(_w_1822));
  bfr _b_1399(.a(_w_1818),.q(_w_1819));
  bfr _b_1398(.a(_w_1817),.q(_w_1818));
  bfr _b_1396(.a(_w_1815),.q(_w_1816));
  bfr _b_1394(.a(_w_1813),.q(_w_1814));
  bfr _b_1391(.a(_w_1810),.q(_w_1811));
  bfr _b_1388(.a(_w_1807),.q(_w_1808));
  bfr _b_1387(.a(_w_1806),.q(_w_1807));
  bfr _b_1384(.a(_w_1803),.q(_w_1804));
  bfr _b_1381(.a(_w_1800),.q(_w_1801));
  bfr _b_1380(.a(_w_1799),.q(_w_1800));
  bfr _b_1379(.a(_w_1798),.q(_w_1799));
  bfr _b_1378(.a(_w_1797),.q(_w_1798));
  bfr _b_1377(.a(_w_1796),.q(_w_1797));
  bfr _b_1413(.a(_w_1832),.q(_w_1833));
  bfr _b_1375(.a(_w_1794),.q(_w_1795));
  bfr _b_1374(.a(_w_1793),.q(N21_5));
  bfr _b_1373(.a(_w_1792),.q(_w_1793));
  bfr _b_1371(.a(_w_1790),.q(_w_1791));
  bfr _b_1369(.a(_w_1788),.q(_w_1789));
  bfr _b_1366(.a(_w_1785),.q(_w_1786));
  bfr _b_1364(.a(_w_1783),.q(_w_1784));
  bfr _b_1359(.a(_w_1778),.q(_w_1779));
  bfr _b_1357(.a(_w_1776),.q(_w_1777));
  bfr _b_1356(.a(_w_1775),.q(_w_1776));
  bfr _b_1355(.a(_w_1774),.q(_w_1775));
  bfr _b_1354(.a(_w_1773),.q(_w_1774));
  bfr _b_1352(.a(_w_1771),.q(_w_1772));
  bfr _b_1351(.a(_w_1770),.q(_w_1771));
  bfr _b_1350(.a(_w_1769),.q(N81_5));
  bfr _b_1349(.a(_w_1768),.q(_w_1769));
  bfr _b_1348(.a(_w_1767),.q(_w_1768));
  bfr _b_1347(.a(_w_1766),.q(_w_1767));
  bfr _b_1460(.a(_w_1879),.q(_w_1880));
  bfr _b_1345(.a(_w_1764),.q(_w_1765));
  bfr _b_1341(.a(_w_1760),.q(_w_1761));
  bfr _b_1338(.a(_w_1757),.q(_w_1758));
  bfr _b_1337(.a(_w_1756),.q(_w_1757));
  bfr _b_1336(.a(_w_1755),.q(_w_1756));
  bfr _b_1335(.a(_w_1754),.q(_w_1755));
  bfr _b_1334(.a(_w_1753),.q(_w_1754));
  bfr _b_1330(.a(_w_1749),.q(_w_1750));
  bfr _b_1329(.a(_w_1748),.q(_w_1749));
  bfr _b_1328(.a(_w_1747),.q(_w_1748));
  bfr _b_1325(.a(_w_1744),.q(_w_1745));
  bfr _b_1332(.a(_w_1751),.q(_w_1752));
  bfr _b_1322(.a(_w_1741),.q(_w_1742));
  bfr _b_1321(.a(_w_1740),.q(_w_1741));
  bfr _b_1525(.a(_w_1944),.q(_w_1945));
  bfr _b_1319(.a(_w_1738),.q(_w_1739));
  bfr _b_1317(.a(_w_1736),.q(_w_1737));
  bfr _b_1314(.a(_w_1733),.q(_w_1734));
  bfr _b_1312(.a(_w_1731),.q(_w_1732));
  bfr _b_1397(.a(_w_1816),.q(_w_1817));
  bfr _b_1311(.a(_w_1730),.q(_w_1731));
  bfr _b_1307(.a(_w_1726),.q(_w_1727));
  bfr _b_1306(.a(_w_1725),.q(_w_1726));
  bfr _b_1305(.a(_w_1724),.q(_w_1725));
  bfr _b_1304(.a(_w_1723),.q(_w_1724));
  bfr _b_1303(.a(_w_1722),.q(N97_2));
  bfr _b_1302(.a(_w_1721),.q(_w_1722));
  bfr _b_1301(.a(_w_1720),.q(_w_1721));
  bfr _b_1300(.a(_w_1719),.q(n233_7));
  bfr _b_1298(.a(_w_1717),.q(_w_1718));
  bfr _b_1297(.a(_w_1716),.q(_w_1717));
  bfr _b_1295(.a(_w_1714),.q(_w_1715));
  bfr _b_1294(.a(_w_1713),.q(_w_1714));
  bfr _b_1292(.a(_w_1711),.q(_w_1712));
  bfr _b_1291(.a(_w_1710),.q(_w_1711));
  bfr _b_1290(.a(_w_1709),.q(_w_1710));
  bfr _b_1289(.a(_w_1708),.q(n259_4));
  bfr _b_1514(.a(_w_1933),.q(_w_1934));
  bfr _b_1287(.a(_w_1706),.q(_w_1707));
  bfr _b_1286(.a(_w_1705),.q(_w_1706));
  bfr _b_1283(.a(_w_1702),.q(_w_1703));
  bfr _b_1282(.a(_w_1701),.q(n259_2));
  bfr _b_1327(.a(_w_1746),.q(N57_5));
  bfr _b_1280(.a(_w_1699),.q(_w_1700));
  bfr _b_1279(.a(_w_1698),.q(_w_1699));
  bfr _b_1276(.a(_w_1695),.q(n298_1));
  bfr _b_1274(.a(_w_1693),.q(_w_1694));
  bfr _b_1278(.a(_w_1697),.q(_w_1698));
  bfr _b_1272(.a(_w_1691),.q(_w_1692));
  bfr _b_1268(.a(_w_1687),.q(_w_1688));
  bfr _b_1277(.a(_w_1696),.q(_w_1697));
  bfr _b_1267(.a(_w_1686),.q(_w_1687));
  bfr _b_1264(.a(_w_1683),.q(N753));
  bfr _b_1259(.a(_w_1678),.q(N747));
  bfr _b_1258(.a(_w_1677),.q(N746));
  bfr _b_1255(.a(_w_1674),.q(N740));
  bfr _b_1254(.a(_w_1673),.q(n233_5));
  bfr _b_1251(.a(_w_1670),.q(_w_1671));
  bfr _b_1250(.a(_w_1669),.q(_w_1670));
  bfr _b_1249(.a(_w_1668),.q(_w_1669));
  bfr _b_1248(.a(_w_1667),.q(_w_1668));
  bfr _b_1372(.a(_w_1791),.q(_w_1792));
  bfr _b_1246(.a(_w_1665),.q(_w_1666));
  bfr _b_1245(.a(_w_1664),.q(_w_1665));
  bfr _b_1242(.a(_w_1661),.q(_w_1662));
  bfr _b_1241(.a(_w_1660),.q(_w_1661));
  bfr _b_1239(.a(_w_1658),.q(_w_1659));
  bfr _b_1324(.a(_w_1743),.q(_w_1744));
  bfr _b_1235(.a(_w_1654),.q(_w_1655));
  bfr _b_1234(.a(_w_1653),.q(_w_1654));
  bfr _b_1233(.a(_w_1652),.q(_w_1653));
  bfr _b_1361(.a(_w_1780),.q(_w_1781));
  bfr _b_1232(.a(_w_1651),.q(_w_1652));
  bfr _b_1230(.a(_w_1649),.q(N61_5));
  bfr _b_1229(.a(_w_1648),.q(_w_1649));
  bfr _b_1228(.a(_w_1647),.q(_w_1648));
  bfr _b_1227(.a(_w_1646),.q(_w_1647));
  bfr _b_1370(.a(_w_1789),.q(_w_1790));
  bfr _b_1323(.a(_w_1742),.q(_w_1743));
  bfr _b_1226(.a(_w_1645),.q(_w_1646));
  bfr _b_1224(.a(_w_1643),.q(_w_1644));
  bfr _b_1221(.a(_w_1640),.q(_w_1641));
  bfr _b_1270(.a(_w_1689),.q(n316_1));
  bfr _b_1263(.a(_w_1682),.q(N752));
  bfr _b_1220(.a(_w_1639),.q(_w_1640));
  bfr _b_1219(.a(_w_1638),.q(_w_1639));
  bfr _b_1214(.a(_w_1633),.q(_w_1634));
  bfr _b_1213(.a(_w_1632),.q(_w_1633));
  bfr _b_1265(.a(_w_1684),.q(N754));
  bfr _b_1212(.a(_w_1631),.q(_w_1632));
  bfr _b_1211(.a(_w_1630),.q(_w_1631));
  bfr _b_1207(.a(_w_1626),.q(_w_1627));
  bfr _b_1206(.a(_w_1625),.q(N53_5));
  bfr _b_1205(.a(_w_1624),.q(_w_1625));
  bfr _b_1204(.a(_w_1623),.q(_w_1624));
  bfr _b_1482(.a(_w_1901),.q(_w_1902));
  bfr _b_1203(.a(_w_1622),.q(_w_1623));
  bfr _b_1200(.a(_w_1619),.q(_w_1620));
  bfr _b_1549(.a(N133),.q(_w_1969));
  bfr _b_1199(.a(_w_1618),.q(_w_1619));
  bfr _b_1198(.a(_w_1617),.q(_w_1618));
  bfr _b_1196(.a(_w_1615),.q(_w_1616));
  bfr _b_1193(.a(_w_1612),.q(_w_1613));
  bfr _b_1192(.a(_w_1611),.q(_w_1612));
  bfr _b_1191(.a(_w_1610),.q(_w_1611));
  bfr _b_1190(.a(_w_1609),.q(_w_1610));
  bfr _b_1189(.a(_w_1608),.q(_w_1609));
  bfr _b_1188(.a(_w_1607),.q(_w_1608));
  bfr _b_1187(.a(_w_1606),.q(_w_1607));
  bfr _b_1186(.a(_w_1605),.q(_w_1606));
  bfr _b_1389(.a(_w_1808),.q(_w_1809));
  bfr _b_1183(.a(_w_1602),.q(_w_1603));
  bfr _b_1180(.a(_w_1599),.q(_w_1600));
  bfr _b_1179(.a(_w_1598),.q(_w_1599));
  bfr _b_1177(.a(_w_1596),.q(N69_5));
  bfr _b_1176(.a(_w_1595),.q(_w_1596));
  bfr _b_1174(.a(_w_1593),.q(_w_1594));
  bfr _b_1173(.a(_w_1592),.q(_w_1593));
  bfr _b_1171(.a(_w_1590),.q(_w_1591));
  bfr _b_1169(.a(_w_1588),.q(_w_1589));
  bfr _b_1168(.a(_w_1587),.q(_w_1588));
  bfr _b_1167(.a(_w_1586),.q(_w_1587));
  bfr _b_1166(.a(_w_1585),.q(_w_1586));
  bfr _b_1163(.a(_w_1582),.q(_w_1583));
  bfr _b_1162(.a(_w_1581),.q(_w_1582));
  bfr _b_1159(.a(_w_1578),.q(_w_1579));
  bfr _b_1158(.a(_w_1577),.q(_w_1578));
  bfr _b_1157(.a(_w_1576),.q(_w_1577));
  bfr _b_1156(.a(_w_1575),.q(_w_1576));
  bfr _b_1154(.a(_w_1573),.q(N117_2));
  bfr _b_1153(.a(_w_1572),.q(_w_1573));
  bfr _b_1152(.a(_w_1571),.q(_w_1572));
  bfr _b_1150(.a(_w_1569),.q(n154));
  bfr _b_1148(.a(_w_1567),.q(_w_1568));
  bfr _b_1147(.a(_w_1566),.q(N73_5));
  bfr _b_1146(.a(_w_1565),.q(_w_1566));
  bfr _b_1144(.a(_w_1563),.q(_w_1564));
  bfr _b_1142(.a(_w_1561),.q(_w_1562));
  bfr _b_1141(.a(_w_1560),.q(_w_1561));
  bfr _b_1140(.a(_w_1559),.q(_w_1560));
  bfr _b_1138(.a(_w_1557),.q(_w_1558));
  bfr _b_1137(.a(_w_1556),.q(_w_1557));
  bfr _b_1136(.a(_w_1555),.q(_w_1556));
  bfr _b_1133(.a(_w_1552),.q(_w_1553));
  bfr _b_1132(.a(_w_1551),.q(_w_1552));
  bfr _b_1293(.a(_w_1712),.q(_w_1713));
  bfr _b_1131(.a(_w_1550),.q(_w_1551));
  bfr _b_1129(.a(_w_1548),.q(_w_1549));
  bfr _b_1128(.a(_w_1547),.q(_w_1548));
  bfr _b_1127(.a(_w_1546),.q(_w_1547));
  bfr _b_1124(.a(_w_1543),.q(N748));
  bfr _b_1160(.a(_w_1579),.q(_w_1580));
  bfr _b_1122(.a(_w_1541),.q(_w_1542));
  bfr _b_1120(.a(_w_1539),.q(_w_1540));
  bfr _b_1119(.a(_w_1538),.q(_w_1539));
  bfr _b_1118(.a(_w_1537),.q(_w_1538));
  bfr _b_1116(.a(_w_1535),.q(_w_1536));
  bfr _b_1115(.a(_w_1534),.q(_w_1535));
  bfr _b_1114(.a(_w_1533),.q(_w_1534));
  bfr _b_1113(.a(_w_1532),.q(_w_1533));
  bfr _b_1111(.a(_w_1530),.q(_w_1531));
  bfr _b_1110(.a(_w_1529),.q(_w_1530));
  bfr _b_1109(.a(_w_1528),.q(_w_1529));
  bfr _b_1071(.a(_w_1490),.q(N750));
  spl3L N37_s_0(.a(_w_1976),.q0(N37_0),.q1(N37_1),.q2(_w_1937));
  spl3L N49_s_1(.a(N49_2),.q0(N49_3),.q1(N49_4),.q2(_w_1915));
  spl2 N5_s_2(.a(N5_5),.q0(N5_6),.q1(N5_7));
  bfr _b_1310(.a(_w_1729),.q(_w_1730));
  and_bb g93(.a(N13_4),.b(N9_4),.q(n93));
  spl3L N5_s_1(.a(N5_2),.q0(N5_3),.q1(N5_4),.q2(_w_1891));
  bfr _b_1194(.a(_w_1613),.q(_w_1614));
  spl3L N73_s_0(.a(N73),.q0(N73_0),.q1(N73_1),.q2(N73_2));
  and_bi g199(.a(N117_1),.b(N113_1),.q(n199));
  spl3L N21_s_0(.a(N21),.q0(N21_0),.q1(N21_1),.q2(N21_2));
  bfr _b_1495(.a(_w_1914),.q(N5_5));
  spl3L N77_s_0(.a(N77),.q0(N77_0),.q1(N77_1),.q2(N77_2));
  bfr _b_1112(.a(_w_1531),.q(_w_1532));
  and_bi g206(.a(n205),.b(n204),.q(n206));
  spl3L N5_s_0(.a(N5),.q0(N5_0),.q1(N5_1),.q2(N5_2));
  and_bb g359(.a(n235_1),.b(n358_0),.q(n359));
  spl2 g240_s_0(.a(n240),.q0(n240_0),.q1(n240_1));
  bfr _b_1409(.a(_w_1828),.q(_w_1829));
  spl2 g215_s_0(.a(n215),.q0(n215_0),.q1(n215_1));
  and_bb g369(.a(n115_5),.b(n360_2),.q(n369));
  and_bb g374(.a(N77_6),.b(n373_0),.q(n374));
  bfr _b_914(.a(_w_1333),.q(_w_1334));
  spl2 N69_s_2(.a(N69_5),.q0(N69_6),.q1(N69_7));
  spl2 g206_s_0(.a(n206),.q0(n206_0),.q1(n206_1));
  bfr _b_932(.a(_w_1351),.q(_w_1352));
  spl2 N89_s_2(.a(N89_5),.q0(N89_6),.q1(N89_7));
  and_bi g57(.a(n55),.b(n56),.q(n57));
  bfr _b_1125(.a(_w_1544),.q(_w_1545));
  spl3L N89_s_1(.a(N89_2),.q0(N89_3),.q1(N89_4),.q2(_w_1868));
  and_bi g62(.a(n57_1),.b(n60_1),.q(n62));
  bfr _b_1077(.a(_w_1496),.q(_w_1497));
  spl2 N9_s_2(.a(N9_5),.q0(N9_6),.q1(N9_7));
  spl3L N9_s_1(.a(N9_2),.q0(N9_3),.q1(N9_4),.q2(_w_1844));
  and_bi g113(.a(n112_0),.b(n91_0),.q(n113));
  and_bi g201(.a(n200_0),.b(n197_0),.q(n201));
  spl2 g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(n140_1));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(n75_1));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  and_bb g367(.a(N69_7),.b(n365_1),.q(n367));
  bfr _b_824(.a(_w_1243),.q(_w_1244));
  spl2 N117_s_2(.a(N117_5),.q0(N117_6),.q1(N117_7));
  and_bi g314(.a(N29_7),.b(n312_1),.q(n314));
  spl2 N41_s_2(.a(N41_5),.q0(N41_6),.q1(N41_7));
  bfr _b_943(.a(_w_1362),.q(_w_1363));
  or_bb g301(.a(N17_6),.b(n300_0),.q(n301));
  spl4L g146_s_0(.a(n146),.q0(n146_0),.q1(n146_1),.q2(n146_2),.q3(n146_3));
  spl3L N41_s_1(.a(N41_2),.q0(N41_3),.q1(N41_4),.q2(_w_1796));
  spl2 g45_s_0(.a(n45),.q0(n45_0),.q1(n45_1));
  spl4L g318_s_0(.a(n318),.q0(n318_0),.q1(n318_1),.q2(n318_2),.q3(n318_3));
  and_bi g248(.a(n244_0),.b(n247_0),.q(n248));
  spl3L N29_s_0(.a(N29),.q0(N29_0),.q1(N29_1),.q2(N29_2));
  spl3L N57_s_0(.a(N57),.q0(N57_0),.q1(N57_1),.q2(N57_2));
  spl2 g131_s_0(.a(n131),.q0(n131_0),.q1(n131_1));
  spl3L N57_s_1(.a(N57_2),.q0(N57_3),.q1(N57_4),.q2(_w_1723));
  and_bi g131(.a(n129),.b(n130),.q(n131));
  spl3L N97_s_0(.a(N97),.q0(N97_0),.q1(N97_1),.q2(_w_1720));
  bfr _b_976(.a(_w_1395),.q(_w_1396));
  spl4L g233_s_4(.a(n233_7),.q0(n233_8),.q1(n233_9),.q2(n233_10),.q3(n233_11));
  spl2 g233_s_3(.a(n233_5),.q0(n233_6),.q1(_w_1716));
  bfr _b_702(.a(_w_1121),.q(_w_1122));
  spl2 g94_s_0(.a(n94),.q0(n94_0),.q1(n94_1));
  bfr _b_1498(.a(_w_1917),.q(_w_1918));
  and_bi g249(.a(n247_1),.b(n244_1),.q(n249));
  spl4L g78_s_2(.a(n78_4),.q0(n78_5),.q1(n78_6),.q2(n78_7),.q3(n78_8));
  bfr _b_924(.a(_w_1343),.q(_w_1344));
  spl2 g78_s_1(.a(n78_2),.q0(n78_3),.q1(_w_1709));
  or_bb g175(.a(n173),.b(n174),.q(n175));
  spl2 g417_s_0(.a(n417),.q0(n417_0),.q1(n417_1));
  bfr _b_740(.a(_w_1159),.q(_w_1160));
  spl2 g227_s_0(.a(n227),.q0(n227_0),.q1(n227_1));
  spl2 g247_s_0(.a(n247),.q0(n247_0),.q1(n247_1));
  and_bi g190(.a(n188_1),.b(n185_1),.q(n190));
  bfr _b_1135(.a(_w_1554),.q(_w_1555));
  bfr _b_700(.a(_w_1119),.q(_w_1120));
  bfr _b_1386(.a(_w_1805),.q(_w_1806));
  bfr _b_1244(.a(_w_1663),.q(_w_1664));
  bfr _b_873(.a(_w_1292),.q(_w_1293));
  spl2 N61_s_2(.a(N61_5),.q0(N61_6),.q1(N61_7));
  spl4L g278_s_2(.a(n278_4),.q0(n278_5),.q1(n278_6),.q2(n278_7),.q3(n278_8));
  spl2 g373_s_0(.a(n373),.q0(n373_0),.q1(n373_1));
  spl2 g279_s_0(.a(n279),.q0(n279_0),.q1(_w_1696));
  bfr _b_1316(.a(_w_1735),.q(_w_1736));
  or_bb g195(.a(N121_0),.b(N125_0),.q(n195));
  bfr _b_1451(.a(_w_1870),.q(_w_1871));
  bfr _b_1393(.a(_w_1812),.q(_w_1813));
  bfr _b_1343(.a(_w_1762),.q(_w_1763));
  bfr _b_795(.a(_w_1214),.q(_w_1215));
  spl2 g266_s_0(.a(n266),.q0(n266_0),.q1(n266_1));
  spl2 g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1));
  spl2 N29_s_2(.a(N29_5),.q0(N29_6),.q1(N29_7));
  bfr _b_782(.a(_w_1201),.q(_w_1202));
  bfr _b_1339(.a(_w_1758),.q(_w_1759));
  and_bi g58(.a(N65_0),.b(N69_0),.q(n58));
  bfr _b_908(.a(_w_1327),.q(_w_1328));
  spl3L N121_s_0(.a(N121),.q0(N121_0),.q1(N121_1),.q2(N121_2));
  bfr _b_1098(.a(_w_1517),.q(_w_1518));
  bfr _b_1106(.a(_w_1525),.q(_w_1526));
  spl2 g316_s_0(.a(n316),.q0(n316_0),.q1(_w_1685));
  bfr _b_990(.a(_w_1409),.q(_w_1410));
  bfr _b_813(.a(_w_1232),.q(_w_1233));
  spl2 g391_s_0(.a(n391),.q0(n391_0),.q1(n391_1));
  spl4L g115_s_2(.a(n115_4),.q0(n115_5),.q1(n115_6),.q2(n115_7),.q3(n115_8));
  bfr _b_1443(.a(_w_1862),.q(_w_1863));
  bfr _b_1216(.a(_w_1635),.q(_w_1636));
  spl4L g259_s_2(.a(n259_4),.q0(n259_5),.q1(n259_6),.q2(n259_7),.q3(n259_8));
  or_bb g310(.a(N25_7),.b(n308_1),.q(n310));
  bfr _b_1123(.a(_w_1542),.q(N29_5));
  and_bb g196(.a(N121_1),.b(N125_1),.q(n196));
  spl2 g400_s_0(.a(n400),.q0(n400_0),.q1(n400_1));
  bfr _b_1477(.a(_w_1896),.q(_w_1897));
  bfr _b_1385(.a(_w_1804),.q(_w_1805));
  bfr _b_659(.a(_w_1078),.q(_w_1079));
  spl2 g421_s_0(.a(n421),.q0(n421_0),.q1(n421_1));
  and_bb g427(.a(N125_7),.b(n425_1),.q(n427));
  and_bb g425(.a(n152_8),.b(n412_3),.q(n425));
  and_bi g424(.a(n423),.b(n422),.q(_w_1684));
  spl2 g122_s_0(.a(n122),.q0(n122_0),.q1(n122_1));
  bfr _b_1068(.a(_w_1487),.q(_w_1488));
  and_bi g420(.a(n418),.b(n419),.q(_w_1683));
  or_bb g418(.a(N117_6),.b(n417_0),.q(n418));
  spl2 g282_s_0(.a(n282),.q0(n282_0),.q1(n282_1));
  bfr _b_787(.a(_w_1206),.q(_w_1207));
  bfr _b_1415(.a(_w_1834),.q(_w_1835));
  bfr _b_942(.a(_w_1361),.q(_w_1362));
  and_bb g415(.a(N113_7),.b(n413_1),.q(n415));
  and_bb g413(.a(n259_8),.b(n412_0),.q(n413));
  or_bb g85(.a(n83),.b(n84),.q(n85));
  and_bi g261(.a(N117_4),.b(N101_4),.q(n261));
  bfr _b_698(.a(_w_1117),.q(_w_1118));
  bfr _b_1240(.a(_w_1659),.q(_w_1660));
  and_bb g398(.a(N97_7),.b(n396_1),.q(n398));
  or_bb g397(.a(N97_6),.b(n396_0),.q(n397));
  bfr _b_1490(.a(_w_1909),.q(_w_1910));
  and_bi g394(.a(n392),.b(n393),.q(_w_1678));
  or_bb g366(.a(N69_6),.b(n365_0),.q(n366));
  spl2 N85_s_2(.a(N85_5),.q0(N85_6),.q1(N85_7));
  and_bi g390(.a(n389),.b(n388),.q(_w_1677));
  or_bb g152(.a(n150),.b(n151),.q(n152));
  and_bb g387(.a(n115_6),.b(n378_2),.q(n387));
  bfr _b_1260(.a(_w_1679),.q(N33_2));
  and_bi g406(.a(N105_7),.b(n404_1),.q(n406));
  bfr _b_691(.a(_w_1110),.q(_w_1111));
  and_bb g378(.a(n213_1),.b(n377_0),.q(n378));
  and_bb g377(.a(n233_6),.b(n358_1),.q(n377));
  spl2 g243_s_0(.a(n243),.q0(n243_0),.q1(n243_1));
  bfr _b_1035(.a(_w_1454),.q(_w_1455));
  spl2 N37_s_2(.a(N37_5),.q0(N37_6),.q1(N37_7));
  and_bi g371(.a(N73_7),.b(n369_1),.q(n371));
  and_bi g61(.a(n60_0),.b(n57_0),.q(n61));
  and_bi g242(.a(N113_4),.b(N97_4),.q(n242));
  bfr _b_957(.a(_w_1376),.q(_w_1377));
  and_bi g370(.a(n369_0),.b(N73_6),.q(n370));
  bfr _b_1033(.a(_w_1452),.q(_w_1453));
  and_bi g368(.a(n366),.b(n367),.q(_w_1675));
  bfr _b_1342(.a(_w_1761),.q(_w_1762));
  and_bb g365(.a(n278_5),.b(n360_1),.q(n365));
  and_bi g272(.a(n270),.b(n271),.q(n272));
  bfr _b_818(.a(_w_1237),.q(_w_1238));
  bfr _b_1552(.a(N135),.q(_w_1972));
  spl3L N105_s_1(.a(N105_2),.q0(N105_3),.q1(N105_4),.q2(_w_1938));
  bfr _b_981(.a(_w_1400),.q(_w_1401));
  or_bb g355(.a(n153_0),.b(n298_0),.q(n355));
  and_bi g121(.a(N93_4),.b(N77_4),.q(n121));
  spl2 g340_s_0(.a(n340),.q0(n340_0),.q1(n340_1));
  bfr _b_934(.a(_w_1353),.q(_w_1354));
  and_bi g354(.a(n352),.b(n353),.q(n354));
  and_bi g326(.a(n324),.b(n325),.q(N733));
  or_bb g283(.a(N1_6),.b(n282_0),.q(n283));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  or_bb g352(.a(n279_0),.b(n316_0),.q(n352));
  or_bb g350(.a(N61_7),.b(n348_1),.q(n350));
  bfr _b_770(.a(_w_1189),.q(_w_1190));
  bfr _b_940(.a(_w_1359),.q(_w_1360));
  and_bb g349(.a(N61_6),.b(n348_0),.q(n349));
  and_bb g373(.a(n152_5),.b(n360_3),.q(n373));
  and_bi g183(.a(N53_4),.b(N37_4),.q(n183));
  and_bi g347(.a(n346),.b(n345),.q(N738));
  and_bi g246(.a(N81_4),.b(N65_4),.q(n246));
  bfr _b_1121(.a(_w_1540),.q(_w_1541));
  bfr _b_695(.a(_w_1114),.q(N125_5));
  and_bb g342(.a(N53_7),.b(n340_1),.q(n342));
  bfr _b_1222(.a(_w_1641),.q(_w_1642));
  spl2 g275_s_0(.a(n275),.q0(n275_0),.q1(n275_1));
  or_bb g255(.a(n100_3),.b(n137_3),.q(n255));
  bfr _b_1425(.a(_w_1844),.q(_w_1845));
  and_bi g339(.a(n337),.b(n338),.q(N736));
  bfr _b_690(.a(_w_1109),.q(_w_1110));
  and_bb g338(.a(N49_7),.b(n336_1),.q(n338));
  and_bb g336(.a(n335_0),.b(n78_8),.q(n336));
  and_bb g335(.a(n298_3),.b(n317_1),.q(n335));
  bfr _b_1269(.a(_w_1688),.q(_w_1689));
  bfr _b_1087(.a(_w_1506),.q(_w_1507));
  bfr _b_1501(.a(_w_1920),.q(_w_1921));
  and_bi g334(.a(n332),.b(n333),.q(N735));
  and_bb g333(.a(N45_7),.b(n331_1),.q(n333));
  or_bb g184(.a(n182),.b(n183),.q(n184));
  bfr _b_1040(.a(_w_1459),.q(_w_1460));
  or_bb g332(.a(N45_6),.b(n331_0),.q(n332));
  and_bi g330(.a(n329),.b(n328),.q(N734));
  bfr _b_1210(.a(_w_1629),.q(_w_1630));
  bfr _b_898(.a(_w_1317),.q(_w_1318));
  and_bb g328(.a(N41_6),.b(n327_0),.q(n328));
  spl2 N97_s_2(.a(N97_5),.q0(N97_6),.q1(N97_7));
  bfr _b_1243(.a(_w_1662),.q(_w_1663));
  or_bb g324(.a(N37_6),.b(n323_0),.q(n324));
  and_bi g405(.a(n404_0),.b(N105_6),.q(n405));
  and_bb g402(.a(N101_7),.b(n400_1),.q(n402));
  bfr _b_1430(.a(_w_1849),.q(_w_1850));
  bfr _b_780(.a(_w_1199),.q(_w_1200));
  spl4L g335_s_0(.a(n335),.q0(n335_0),.q1(n335_1),.q2(n335_2),.q3(n335_3));
  and_bb g327(.a(n181_8),.b(n318_2),.q(n327));
  bfr _b_1092(.a(_w_1511),.q(_w_1512));
  bfr _b_1545(.a(N131),.q(_w_1965));
  spl2 g327_s_0(.a(n327),.q0(n327_0),.q1(n327_1));
  spl2 g169_s_0(.a(n169),.q0(n169_0),.q1(n169_1));
  bfr _b_838(.a(_w_1257),.q(_w_1258));
  and_bi g322(.a(n320),.b(n321),.q(N732));
  and_bb g391(.a(n152_6),.b(n378_3),.q(n391));
  spl3L N53_s_1(.a(N53_2),.q0(N53_3),.q1(N53_4),.q2(_w_1604));
  bfr _b_1217(.a(_w_1636),.q(_w_1637));
  and_bb g361(.a(n259_5),.b(n360_0),.q(n361));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(n250_1));
  spl2 g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1));
  bfr _b_1143(.a(_w_1562),.q(_w_1563));
  and_bb g319(.a(n318_0),.b(n78_7),.q(n319));
  and_bb g312(.a(n233_9),.b(n299_3),.q(n312));
  bfr _b_1281(.a(_w_1700),.q(n279_1));
  and_bi g311(.a(n310),.b(n309),.q(N730));
  or_bb g127(.a(n116_1),.b(n125_1),.q(n127));
  bfr _b_1416(.a(_w_1835),.q(_w_1836));
  spl2 g210_s_0(.a(n210),.q0(n210_0),.q1(_w_1597));
  or_bb g389(.a(N89_7),.b(n387_1),.q(n389));
  and_bi g307(.a(n305),.b(n306),.q(N729));
  bfr _b_1395(.a(_w_1814),.q(_w_1815));
  bfr _b_1151(.a(_w_1570),.q(N755));
  bfr _b_1139(.a(_w_1558),.q(_w_1559));
  and_bi g219(.a(N13_0),.b(N29_0),.q(n219));
  spl2 g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1));
  bfr _b_1530(.a(_w_1949),.q(_w_1950));
  bfr _b_1401(.a(_w_1820),.q(_w_1821));
  bfr _b_692(.a(_w_1111),.q(_w_1112));
  bfr _b_1063(.a(_w_1482),.q(_w_1483));
  spl3L N69_s_1(.a(N69_2),.q0(N69_3),.q1(N69_4),.q2(_w_1574));
  bfr _b_747(.a(_w_1166),.q(_w_1167));
  or_bb g305(.a(N21_6),.b(n304_0),.q(n305));
  spl3L N117_s_0(.a(N117),.q0(N117_0),.q1(N117_1),.q2(_w_1571));
  bfr _b_988(.a(_w_1407),.q(_w_1408));
  bfr _b_1247(.a(_w_1666),.q(_w_1667));
  or_bb g356(.a(n259_3),.b(n278_3),.q(n356));
  bfr _b_944(.a(_w_1363),.q(N25_5));
  bfr _b_970(.a(_w_1389),.q(_w_1390));
  and_bb g383(.a(n278_6),.b(n378_1),.q(n383));
  and_bb g300(.a(n299_0),.b(n78_6),.q(n300));
  or_bb g92(.a(N13_3),.b(N9_3),.q(n92));
  bfr _b_1023(.a(_w_1442),.q(_w_1443));
  bfr _b_867(.a(_w_1286),.q(_w_1287));
  and_bb g379(.a(n259_6),.b(n378_0),.q(n379));
  and_bb g299(.a(n280_1),.b(n298_2),.q(n299));
  or_bb g167(.a(N105_0),.b(N109_0),.q(n167));
  and_bb g417(.a(n278_8),.b(n412_1),.q(n417));
  bfr _b_1045(.a(_w_1464),.q(_w_1465));
  bfr _b_1479(.a(_w_1898),.q(_w_1899));
  spl2 N33_s_2(.a(N33_5),.q0(N33_6),.q1(N33_7));
  and_bi g162(.a(n157_1),.b(n160_1),.q(n162));
  and_bi g158(.a(N9_0),.b(N25_0),.q(n158));
  bfr _b_797(.a(_w_1216),.q(_w_1217));
  and_bi g105(.a(N37_1),.b(N33_1),.q(n105));
  spl4L g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1),.q2(n137_2),.q3(n137_3));
  and_bi g428(.a(n426),.b(n427),.q(_w_1570));
  or_bb g423(.a(N121_7),.b(n421_1),.q(n423));
  bfr _b_1447(.a(_w_1866),.q(_w_1867));
  bfr _b_1073(.a(_w_1492),.q(_w_1493));
  and_bi g155(.a(N41_0),.b(N57_0),.q(n155));
  spl2 g359_s_0(.a(n359),.q0(n359_0),.q1(n359_1));
  bfr _b_714(.a(_w_1133),.q(_w_1134));
  and_bi g289(.a(n287),.b(n288),.q(N725));
  bfr _b_1445(.a(_w_1864),.q(_w_1865));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(n88_1));
  bfr _b_814(.a(_w_1233),.q(_w_1234));
  and_bb g421(.a(n115_8),.b(n412_2),.q(n421));
  and_bb g147(.a(n137_0),.b(n146_0),.q(n147));
  spl3L N37_s_1(.a(N37_2),.q0(N37_3),.q1(N37_4),.q2(_w_1650));
  or_bb g240(.a(n234),.b(n239),.q(n240));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(n112_1));
  and_bi g236(.a(n233_2),.b(n181_4),.q(n236));
  bfr _b_1527(.a(_w_1946),.q(_w_1947));
  bfr _b_1518(.a(_w_1937),.q(N37_2));
  and_bb g282(.a(n281_0),.b(n78_5),.q(n282));
  bfr _b_1145(.a(_w_1564),.q(_w_1565));
  spl2 g269_s_0(.a(n269),.q0(n269_0),.q1(n269_1));
  and_bi g151(.a(n128_1),.b(n149_1),.q(n151));
  spl2 g365_s_0(.a(n365),.q0(n365_0),.q1(n365_1));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(n119_1));
  bfr _b_750(.a(_w_1169),.q(_w_1170));
  and_bb g318(.a(n153_3),.b(n317_0),.q(n318));
  bfr _b_880(.a(_w_1299),.q(_w_1300));
  bfr _b_1130(.a(_w_1549),.q(_w_1550));
  bfr _b_890(.a(_w_1309),.q(N113_5));
  and_bi g144(.a(n143_0),.b(n140_0),.q(n144));
  and_bi g140(.a(n138),.b(n139),.q(n140));
  or_bb g138(.a(N57_3),.b(N61_3),.q(n138));
  or_bb g329(.a(N41_7),.b(n327_1),.q(n329));
  or_bb g88(.a(n86),.b(n87),.q(n88));
  or_bb g137(.a(n135),.b(n136),.q(n137));
  and_bb g154(.a(_w_1964),.b(N137_6),.q(_w_1567));
  or_bb g353(.a(n115_3),.b(n152_3),.q(n353));
  bfr _b_794(.a(_w_1213),.q(_w_1214));
  or_bb g90(.a(n79_1),.b(n88_1),.q(n90));
  and_bi g95(.a(N1_3),.b(N5_3),.q(n95));
  bfr _b_1426(.a(_w_1845),.q(_w_1846));
  spl2 g387_s_0(.a(n387),.q0(n387_0),.q1(n387_1));
  bfr _b_784(.a(_w_1203),.q(_w_1204));
  or_bb g209(.a(n207),.b(n208),.q(n209));
  bfr _b_1275(.a(_w_1694),.q(_w_1695));
  spl2 g116_s_0(.a(n116),.q0(n116_0),.q1(n116_1));
  and_bi g174(.a(n169_1),.b(n172_1),.q(n174));
  bfr _b_1273(.a(_w_1692),.q(_w_1693));
  bfr _b_861(.a(_w_1280),.q(_w_1281));
  or_bb g160(.a(n158),.b(n159),.q(n160));
  spl2 g404_s_0(.a(n404),.q0(n404_0),.q1(n404_1));
  and_bb g254(.a(n100_2),.b(n137_2),.q(n254));
  spl2 g51_s_0(.a(n51),.q0(n51_0),.q1(n51_1));
  bfr _b_1483(.a(_w_1902),.q(_w_1903));
  bfr _b_737(.a(_w_1156),.q(_w_1157));
  and_bb g130(.a(N25_4),.b(N29_4),.q(n130));
  bfr _b_967(.a(_w_1386),.q(N77_5));
  or_bb g129(.a(N25_3),.b(N29_3),.q(n129));
  and_bb g53(.a(n44_1),.b(n51_1),.q(n53));
  and_bb g395(.a(n210_1),.b(n359_1),.q(n395));
  spl3L N73_s_1(.a(N73_2),.q0(N73_3),.q1(N73_4),.q2(_w_1544));
  bfr _b_1117(.a(_w_1536),.q(_w_1537));
  and_bi g187(.a(N21_1),.b(N5_1),.q(n187));
  and_bb g168(.a(N105_1),.b(N109_1),.q(n168));
  and_bi g296(.a(N13_7),.b(n294_1),.q(n296));
  and_bi g128(.a(n127),.b(n126),.q(n128));
  and_bb g193(.a(n184_1),.b(n191_1),.q(n193));
  bfr _b_926(.a(_w_1345),.q(_w_1346));
  and_bb g126(.a(n116_0),.b(n125_0),.q(n126));
  bfr _b_1531(.a(_w_1950),.q(_w_1951));
  or_bb g125(.a(n123),.b(n124),.q(n125));
  bfr _b_696(.a(_w_1115),.q(_w_1116));
  bfr _b_1362(.a(_w_1781),.q(_w_1782));
  bfr _b_1215(.a(_w_1634),.q(_w_1635));
  or_bb g375(.a(N77_7),.b(n373_1),.q(n375));
  and_bi g194(.a(n192),.b(n193),.q(n194));
  and_bi g123(.a(n122_0),.b(n119_0),.q(n123));
  and_bi g399(.a(n397),.b(n398),.q(_w_1543));
  bfr _b_1253(.a(_w_1672),.q(n278_2));
  spl3L N41_s_0(.a(N41),.q0(N41_0),.q1(N41_1),.q2(N41_2));
  and_bb g381(.a(N81_7),.b(n379_1),.q(n381));
  and_bb g325(.a(N37_7),.b(n323_1),.q(n325));
  or_bb g119(.a(n117),.b(n118),.q(n119));
  bfr _b_844(.a(_w_1263),.q(_w_1264));
  bfr _b_1318(.a(_w_1737),.q(_w_1738));
  and_bi g256(.a(n255),.b(n254),.q(n256));
  and_bi g118(.a(N125_4),.b(N109_4),.q(n118));
  or_bb g297(.a(n295),.b(n296),.q(N727));
  spl3L N29_s_1(.a(N29_2),.q0(N29_3),.q1(N29_4),.q2(_w_1519));
  spl2 g312_s_0(.a(n312),.q0(n312_0),.q1(n312_1));
  or_bb g250(.a(n248),.b(n249),.q(n250));
  bfr _b_853(.a(_w_1272),.q(N85_5));
  or_bb g270(.a(n262_0),.b(n269_0),.q(n270));
  and_bi g112(.a(n111),.b(n110),.q(n112));
  and_bi g234(.a(n214),.b(n233_4),.q(n234));
  or_bb g111(.a(n100_1),.b(n109_1),.q(n111));
  spl2 g262_s_0(.a(n262),.q0(n262_0),.q1(n262_1));
  and_bb g110(.a(n100_0),.b(n109_0),.q(n110));
  and_bb g408(.a(n152_7),.b(n395_3),.q(n408));
  and_bi g222(.a(n221_0),.b(n218_0),.q(n222));
  and_bi g220(.a(N29_1),.b(N13_1),.q(n220));
  bfr _b_1201(.a(_w_1620),.q(_w_1621));
  spl2 g348_s_0(.a(n348),.q0(n348_0),.q1(n348_1));
  bfr _b_836(.a(_w_1255),.q(_w_1256));
  and_bi g150(.a(n149_0),.b(n128_0),.q(n150));
  or_bb g63(.a(n61),.b(n62),.q(n63));
  and_bb g164(.a(n154_0),.b(n163_0),.q(n164));
  and_bb g306(.a(N21_7),.b(n304_1),.q(n306));
  bfr _b_1439(.a(_w_1858),.q(_w_1859));
  bfr _b_1363(.a(_w_1782),.q(_w_1783));
  bfr _b_1288(.a(_w_1707),.q(_w_1708));
  bfr _b_1091(.a(_w_1510),.q(_w_1511));
  and_bb g102(.a(N41_4),.b(N45_4),.q(n102));
  spl2 g57_s_0(.a(n57),.q0(n57_0),.q1(n57_1));
  or_bb g337(.a(N49_6),.b(n336_0),.q(n337));
  and_bb g56(.a(N73_1),.b(N77_1),.q(n56));
  bfr _b_1085(.a(_w_1504),.q(_w_1505));
  bfr _b_1042(.a(_w_1461),.q(_w_1462));
  spl2 N73_s_2(.a(N73_5),.q0(N73_6),.q1(N73_7));
  spl2 g233_s_2(.a(n233_3),.q0(n233_4),.q1(_w_1673));
  bfr _b_1043(.a(_w_1462),.q(_w_1463));
  and_bi g135(.a(n134_0),.b(n131_0),.q(n135));
  and_bb g176(.a(n175_0),.b(n63_2),.q(n176));
  and_bi g66(.a(n64),.b(n65),.q(n66));
  or_bb g64(.a(N89_0),.b(N93_0),.q(n64));
  and_bb g321(.a(N33_7),.b(n319_1),.q(n321));
  and_bi g161(.a(n160_0),.b(n157_0),.q(n161));
  bfr _b_1484(.a(_w_1903),.q(_w_1904));
  and_bb g294(.a(n233_8),.b(n281_3),.q(n294));
  and_bi g46(.a(N1_0),.b(N17_0),.q(n46));
  spl2 g244_s_0(.a(n244),.q0(n244_0),.q1(n244_1));
  bfr _b_1170(.a(_w_1589),.q(_w_1590));
  and_bi g42(.a(N33_3),.b(N49_3),.q(n42));
  spl2 g256_s_0(.a(n256),.q0(n256_0),.q1(n256_1));
  spl2 g323_s_0(.a(n323),.q0(n323_0),.q1(n323_1));
  and_bi g91(.a(n90),.b(n89),.q(n91));
  and_bi g313(.a(n312_0),.b(N29_6),.q(n313));
  and_bi g156(.a(N57_1),.b(N41_1),.q(n156));
  bfr _b_1079(.a(_w_1498),.q(_w_1499));
  spl3L N45_s_1(.a(N45_2),.q0(N45_3),.q1(N45_4),.q2(_w_1491));
  and_bi g75(.a(n74),.b(n73),.q(n75));
  spl2 g263_s_0(.a(n263),.q0(n263_0),.q1(n263_1));
  and_bi g217(.a(N61_1),.b(N45_1),.q(n217));
  bfr _b_1414(.a(_w_1833),.q(_w_1834));
  and_bb g73(.a(n63_0),.b(n72_0),.q(n73));
  or_bb g407(.a(n405),.b(n406),.q(_w_1490));
  and_bi g108(.a(n103_1),.b(n106_1),.q(n108));
  and_bi g47(.a(N17_1),.b(N1_1),.q(n47));
  spl2 g413_s_0(.a(n413),.q0(n413_0),.q1(n413_1));
  and_bb g45(.a(_w_1961),.b(N137_0),.q(_w_1489));
  bfr _b_1436(.a(_w_1855),.q(_w_1856));
  bfr _b_701(.a(_w_1120),.q(_w_1121));
  and_bb g385(.a(N85_7),.b(n383_1),.q(n385));
  bfr _b_875(.a(_w_1294),.q(_w_1295));
  and_bi g197(.a(n195),.b(n196),.q(n197));
  spl2 g166_s_0(.a(n166),.q0(n166_0),.q1(n166_1));
  bfr _b_1237(.a(_w_1656),.q(_w_1657));
  or_bb g203(.a(n201),.b(n202),.q(n203));
  bfr _b_713(.a(_w_1132),.q(_w_1133));
  bfr _b_820(.a(_w_1239),.q(_w_1240));
  and_bi g141(.a(N49_0),.b(N53_0),.q(n141));
  and_bi g59(.a(N69_1),.b(N65_1),.q(n59));
  spl3L N33_s_1(.a(N33_2),.q0(N33_3),.q1(N33_4),.q2(_w_1467));
  and_bi g43(.a(N49_4),.b(N33_4),.q(n43));
  and_bi g182(.a(N37_3),.b(N53_3),.q(n182));
  or_bb g191(.a(n189),.b(n190),.q(n191));
  spl4L g395_s_0(.a(n395),.q0(n395_0),.q1(n395_1),.q2(n395_2),.q3(n395_3));
  or_bb g237(.a(n235_0),.b(n236),.q(n237));
  spl2 g253_s_0(.a(n253),.q0(n253_0),.q1(n253_1));
  bfr _b_1423(.a(_w_1842),.q(_w_1843));
  and_bb g396(.a(n259_7),.b(n395_0),.q(n396));
  bfr _b_1432(.a(_w_1851),.q(_w_1852));
  and_bb g393(.a(N93_7),.b(n391_1),.q(n393));
  or_bb g269(.a(n267),.b(n268),.q(n269));
  or_bb g287(.a(N5_6),.b(n286_0),.q(n287));
  bfr _b_1266(.a(_w_1685),.q(_w_1686));
  bfr _b_1172(.a(_w_1591),.q(_w_1592));
  and_bi g49(.a(n45_0),.b(n48_0),.q(n49));
  and_bi g376(.a(n375),.b(n374),.q(_w_1466));
  or_bb g165(.a(n154_1),.b(n163_1),.q(n165));
  bfr _b_999(.a(_w_1418),.q(_w_1419));
  bfr _b_1178(.a(_w_1597),.q(_w_1598));
  spl4L g360_s_0(.a(n360),.q0(n360_0),.q1(n360_1),.q2(n360_2),.q3(n360_3));
  spl2 g383_s_0(.a(n383),.q0(n383_0),.q1(n383_1));
  spl3L N125_s_0(.a(N125),.q0(N125_0),.q1(N125_1),.q2(N125_2));
  and_bb g302(.a(N17_7),.b(n300_1),.q(n302));
  bfr _b_733(.a(_w_1152),.q(_w_1153));
  and_bi g178(.a(n177),.b(n176),.q(n178));
  bfr _b_1434(.a(_w_1853),.q(_w_1854));
  and_bi g186(.a(N5_0),.b(N21_0),.q(n186));
  bfr _b_1025(.a(_w_1444),.q(_w_1445));
  bfr _b_863(.a(_w_1282),.q(_w_1283));
  bfr _b_726(.a(_w_1145),.q(n152_2));
  spl2 g233_s_0(.a(n233),.q0(n233_0),.q1(n233_1));
  bfr _b_1027(.a(_w_1446),.q(_w_1447));
  or_bb g55(.a(N73_0),.b(N77_0),.q(n55));
  and_bi g245(.a(N65_3),.b(N81_3),.q(n245));
  bfr _b_767(.a(_w_1186),.q(_w_1187));
  and_bi g77(.a(n54_1),.b(n75_1),.q(n77));
  bfr _b_1149(.a(_w_1568),.q(_w_1569));
  bfr _b_1086(.a(_w_1505),.q(_w_1506));
  bfr _b_1082(.a(_w_1501),.q(_w_1502));
  bfr _b_1557(.a(N37),.q(_w_1976));
  spl2 g308_s_0(.a(n308),.q0(n308_0),.q1(n308_1));
  and_bb g345(.a(N57_6),.b(n344_0),.q(n345));
  bfr _b_1165(.a(_w_1584),.q(_w_1585));
  or_bb g218(.a(n216),.b(n217),.q(n218));
  spl3L N13_s_1(.a(N13_2),.q0(N13_3),.q1(N13_4),.q2(_w_1442));
  bfr _b_859(.a(_w_1278),.q(_w_1279));
  and_bi g132(.a(N17_3),.b(N21_3),.q(n132));
  spl3L g115_s_0(.a(n115),.q0(n115_0),.q1(n115_1),.q2(_w_1441));
  bfr _b_1231(.a(_w_1650),.q(_w_1651));
  bfr _b_647(.a(_w_1066),.q(n212_1));
  and_bi g83(.a(N73_3),.b(N89_3),.q(n83));
  bfr _b_1467(.a(_w_1886),.q(_w_1887));
  bfr _b_643(.a(_w_1062),.q(_w_1063));
  spl2 N57_s_2(.a(N57_5),.q0(N57_6),.q1(N57_7));
  spl2 g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1));
  spl3L g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1),.q2(_w_1438));
  spl3L N9_s_0(.a(N9),.q0(N9_0),.q1(N9_1),.q2(N9_2));
  spl2 g425_s_0(.a(n425),.q0(n425_0),.q1(n425_1));
  or_bb g414(.a(N113_6),.b(n413_0),.q(n414));
  spl3L N93_s_1(.a(N93_2),.q0(N93_3),.q1(N93_4),.q2(_w_1414));
  and_bb g404(.a(n115_7),.b(n395_2),.q(n404));
  and_bb g308(.a(n181_7),.b(n299_2),.q(n308));
  bfr _b_1134(.a(_w_1553),.q(_w_1554));
  spl2 g317_s_0(.a(n317),.q0(n317_0),.q1(n317_1));
  bfr _b_731(.a(_w_1150),.q(n211_1));
  or_bb g251(.a(n243_0),.b(n250_0),.q(n251));
  or_bb g315(.a(n313),.b(n314),.q(N731));
  spl2 g230_s_0(.a(n230),.q0(n230_0),.q1(n230_1));
  and_bi g298(.a(n152_1),.b(n115_1),.q(n298));
  or_bb g163(.a(n161),.b(n162),.q(n163));
  and_bb g65(.a(N89_1),.b(N93_1),.q(n65));
  and_bi g50(.a(n48_1),.b(n45_1),.q(n50));
  and_bi g84(.a(N89_4),.b(N73_4),.q(n84));
  bfr _b_668(.a(_w_1087),.q(_w_1088));
  bfr _b_746(.a(_w_1165),.q(_w_1166));
  bfr _b_1529(.a(_w_1948),.q(_w_1949));
  and_bb g340(.a(n209_8),.b(n335_1),.q(n340));
  bfr _b_964(.a(_w_1383),.q(_w_1384));
  or_bb g143(.a(n141),.b(n142),.q(n143));
  bfr _b_1181(.a(_w_1600),.q(_w_1601));
  bfr _b_1103(.a(_w_1522),.q(_w_1523));
  spl2 g125_s_0(.a(n125),.q0(n125_0),.q1(n125_1));
  and_bi g265(.a(N85_4),.b(N69_4),.q(n265));
  and_bi g207(.a(n206_0),.b(n194_0),.q(n207));
  and_bb g360(.a(n212_1),.b(n359_0),.q(n360));
  bfr _b_769(.a(_w_1188),.q(_w_1189));
  and_bi g114(.a(n91_1),.b(n112_1),.q(n114));
  bfr _b_1457(.a(_w_1876),.q(_w_1877));
  or_bb g122(.a(n120),.b(n121),.q(n122));
  and_bi g86(.a(n85_0),.b(n82_0),.q(n86));
  spl3L N65_s_0(.a(N65),.q0(N65_0),.q1(N65_1),.q2(N65_2));
  or_bb g134(.a(n132),.b(n133),.q(n134));
  spl4L g72_s_0(.a(n72),.q0(n72_0),.q1(n72_1),.q2(n72_2),.q3(n72_3));
  and_bb g89(.a(n79_0),.b(n88_0),.q(n89));
  bfr _b_652(.a(_w_1071),.q(_w_1072));
  or_bb g52(.a(n44_0),.b(n51_0),.q(n52));
  and_bb g363(.a(N65_7),.b(n361_1),.q(n363));
  and_bi g99(.a(n94_1),.b(n97_1),.q(n99));
  spl4L N137_s_2(.a(N137_3),.q0(N137_6),.q1(N137_7),.q2(N137_8),.q3(N137_9));
  and_bi g76(.a(n75_0),.b(n54_0),.q(n76));
  bfr _b_1271(.a(_w_1690),.q(_w_1691));
  and_bi g107(.a(n106_0),.b(n103_0),.q(n107));
  bfr _b_666(.a(_w_1085),.q(_w_1086));
  bfr _b_832(.a(_w_1251),.q(_w_1252));
  or_bb g100(.a(n98),.b(n99),.q(n100));
  bfr _b_730(.a(_w_1149),.q(_w_1150));
  bfr _b_1256(.a(_w_1675),.q(N741));
  bfr _b_765(.a(_w_1184),.q(_w_1185));
  and_bi g103(.a(n101),.b(n102),.q(n103));
  or_bb g72(.a(n70),.b(n71),.q(n72));
  spl3L N117_s_1(.a(N117_2),.q0(N117_3),.q1(N117_4),.q2(_w_1394));
  spl2 g286_s_0(.a(n286),.q0(n286_0),.q1(n286_1));
  and_bi g208(.a(n194_1),.b(n206_1),.q(n208));
  and_bi g213(.a(n212_0),.b(n181_1),.q(n213));
  and_bi g169(.a(n167),.b(n168),.q(n169));
  and_bi g170(.a(N97_0),.b(N101_0),.q(n170));
  bfr _b_1218(.a(_w_1637),.q(_w_1638));
  and_bb g290(.a(n181_6),.b(n281_2),.q(n290));
  and_bi g285(.a(n283),.b(n284),.q(N724));
  and_bi g171(.a(N101_1),.b(N97_1),.q(n171));
  spl3L N81_s_1(.a(N81_2),.q0(N81_3),.q1(N81_4),.q2(_w_1747));
  spl2 g377_s_0(.a(n377),.q0(n377_0),.q1(n377_1));
  spl3L N53_s_0(.a(_w_1978),.q0(N53_0),.q1(N53_1),.q2(_w_1393));
  bfr _b_1000(.a(_w_1419),.q(_w_1420));
  bfr _b_1340(.a(_w_1759),.q(_w_1760));
  and_bi g173(.a(n172_0),.b(n169_0),.q(n173));
  or_bb g426(.a(N125_6),.b(n425_0),.q(n426));
  bfr _b_882(.a(_w_1301),.q(_w_1302));
  bfr _b_1257(.a(_w_1676),.q(N742));
  and_bb g252(.a(n243_1),.b(n250_1),.q(n252));
  and_bi g179(.a(n178_0),.b(n166_0),.q(n179));
  bfr _b_1344(.a(_w_1763),.q(_w_1764));
  and_bb g317(.a(n240_1),.b(n316_1),.q(n317));
  bfr _b_899(.a(_w_1318),.q(_w_1319));
  and_bi g180(.a(n166_1),.b(n178_1),.q(n180));
  bfr _b_1532(.a(_w_1951),.q(_w_1952));
  bfr _b_1464(.a(_w_1883),.q(_w_1884));
  bfr _b_1309(.a(_w_1728),.q(_w_1729));
  or_bb g82(.a(n80),.b(n81),.q(n82));
  spl2 g221_s_0(.a(n221),.q0(n221_0),.q1(n221_1));
  and_bb g412(.a(n211_1),.b(n377_1),.q(n412));
  bfr _b_915(.a(_w_1334),.q(_w_1335));
  and_bi g216(.a(N45_0),.b(N61_0),.q(n216));
  and_bb g228(.a(n203_2),.b(n72_2),.q(n228));
  or_bb g358(.a(n354),.b(n357),.q(n358));
  spl3L N25_s_0(.a(N25),.q0(N25_0),.q1(N25_1),.q2(N25_2));
  or_bb g346(.a(N57_7),.b(n344_1),.q(n346));
  bfr _b_1517(.a(_w_1936),.q(N49_5));
  and_bi g264(.a(N69_3),.b(N85_3),.q(n264));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(_w_1387));
  and_bb g185(.a(_w_1962),.b(N137_7),.q(n185));
  or_bb g188(.a(n186),.b(n187),.q(n188));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  bfr _b_1313(.a(_w_1732),.q(_w_1733));
  and_bi g241(.a(N97_3),.b(N113_3),.q(n241));
  and_bb g291(.a(N9_6),.b(n290_0),.q(n291));
  bfr _b_1028(.a(_w_1447),.q(_w_1448));
  spl3L N77_s_1(.a(N77_2),.q0(N77_3),.q1(N77_4),.q2(_w_1364));
  bfr _b_849(.a(_w_1268),.q(_w_1269));
  bfr _b_856(.a(_w_1275),.q(_w_1276));
  bfr _b_1029(.a(_w_1448),.q(_w_1449));
  spl2 g143_s_0(.a(n143),.q0(n143_0),.q1(n143_1));
  and_bb g271(.a(n262_1),.b(n269_1),.q(n271));
  spl2 N77_s_2(.a(N77_5),.q0(N77_6),.q1(N77_7));
  and_bi g166(.a(n165),.b(n164),.q(n166));
  and_bb g409(.a(N109_6),.b(n408_0),.q(n409));
  or_bb g320(.a(N33_6),.b(n319_0),.q(n320));
  spl2 g218_s_0(.a(n218),.q0(n218_0),.q1(n218_1));
  and_bb g273(.a(n109_2),.b(n146_2),.q(n273));
  or_bb g200(.a(n198),.b(n199),.q(n200));
  spl3L N85_s_0(.a(N85),.q0(N85_0),.q1(N85_1),.q2(N85_2));
  spl4L g412_s_0(.a(n412),.q0(n412_0),.q1(n412_1),.q2(n412_2),.q3(n412_3));
  or_bb g157(.a(n155),.b(n156),.q(n157));
  and_bb g331(.a(n233_10),.b(n318_3),.q(n331));
  or_bb g380(.a(N81_6),.b(n379_0),.q(n380));
  bfr _b_772(.a(_w_1191),.q(_w_1192));
  and_bi g268(.a(n266_1),.b(n263_1),.q(n268));
  spl2 N45_s_2(.a(N45_5),.q0(N45_6),.q1(N45_7));
  and_bb g244(.a(_w_1968),.b(N137_9),.q(_w_1339));
  spl2 g163_s_0(.a(n163),.q0(n163_0),.q1(n163_1));
  or_bb g292(.a(N9_7),.b(n290_1),.q(n292));
  spl2 g278_s_1(.a(n278_2),.q0(n278_3),.q1(_w_1332));
  bfr _b_684(.a(_w_1103),.q(_w_1104));
  or_bb g392(.a(N93_6),.b(n391_0),.q(n392));
  and_bi g117(.a(N109_3),.b(N125_3),.q(n117));
  bfr _b_912(.a(_w_1331),.q(N49_2));
  and_bi g202(.a(n197_1),.b(n200_1),.q(n202));
  bfr _b_1320(.a(_w_1739),.q(_w_1740));
  spl2 N13_s_2(.a(N13_5),.q0(N13_6),.q1(N13_7));
  bfr _b_1175(.a(_w_1594),.q(_w_1595));
  bfr _b_660(.a(_w_1079),.q(_w_1080));
  or_bb g226(.a(n215_1),.b(n224_1),.q(n226));
  and_bb g400(.a(n278_7),.b(n395_1),.q(n400));
  spl2 g157_s_0(.a(n157),.q0(n157_0),.q1(n157_1));
  and_bi g198(.a(N113_0),.b(N117_0),.q(n198));
  bfr _b_688(.a(_w_1107),.q(_w_1108));
  and_bb g204(.a(n175_2),.b(n203_0),.q(n204));
  bfr _b_1195(.a(_w_1614),.q(_w_1615));
  and_bi g316(.a(n278_1),.b(n259_1),.q(n316));
  bfr _b_760(.a(_w_1179),.q(_w_1180));
  or_bb g372(.a(n370),.b(n371),.q(_w_1676));
  bfr _b_922(.a(_w_1341),.q(_w_1342));
  bfr _b_928(.a(_w_1347),.q(_w_1348));
  and_bi g258(.a(n253_1),.b(n256_1),.q(n258));
  or_bb g106(.a(n104),.b(n105),.q(n106));
  or_bb g115(.a(n113),.b(n114),.q(n115));
  spl2 g272_s_0(.a(n272),.q0(n272_0),.q1(n272_1));
  spl2 N81_s_2(.a(N81_5),.q0(N81_6),.q1(N81_7));
  and_bb g288(.a(N5_7),.b(n286_1),.q(n288));
  spl2 g91_s_0(.a(n91),.q0(n91_0),.q1(n91_1));
  and_bi g295(.a(n294_0),.b(N13_6),.q(n295));
  bfr _b_1083(.a(_w_1502),.q(_w_1503));
  or_bb g74(.a(n63_1),.b(n72_1),.q(n74));
  and_bi g210(.a(n209_0),.b(n78_0),.q(n210));
  and_bi g253(.a(n251),.b(n252),.q(n253));
  and_bi g211(.a(n210_0),.b(n181_0),.q(n211));
  bfr _b_1358(.a(_w_1777),.q(_w_1778));
  bfr _b_706(.a(_w_1125),.q(_w_1126));
  spl3L N49_s_0(.a(_w_1977),.q0(N49_0),.q1(N49_1),.q2(_w_1331));
  bfr _b_754(.a(_w_1173),.q(N101_2));
  bfr _b_1543(.a(N130),.q(_w_1963));
  spl3L g278_s_0(.a(n278),.q0(n278_0),.q1(n278_1),.q2(_w_1672));
  and_bi g70(.a(n69_0),.b(n66_0),.q(n70));
  and_bi g382(.a(n380),.b(n381),.q(_w_1310));
  and_bi g343(.a(n341),.b(n342),.q(N737));
  spl2 g213_s_0(.a(n213),.q0(n213_0),.q1(_w_1285));
  bfr _b_1236(.a(_w_1655),.q(_w_1656));
  and_bi g67(.a(N81_0),.b(N85_0),.q(n67));
  or_bb g214(.a(n211_0),.b(n213_0),.q(n214));
  bfr _b_1360(.a(_w_1779),.q(_w_1780));
  or_bb g384(.a(N85_6),.b(n383_0),.q(n384));
  bfr _b_858(.a(_w_1277),.q(n233_3));
  and_bb g225(.a(n215_0),.b(n224_0),.q(n225));
  bfr _b_1056(.a(_w_1475),.q(_w_1476));
  or_bb g274(.a(n109_3),.b(n146_3),.q(n274));
  spl3L g259_s_0(.a(n259),.q0(n259_0),.q1(n259_1),.q2(_w_1701));
  and_bb g116(.a(_w_1973),.b(N137_5),.q(_w_1278));
  and_bb g215(.a(_w_1966),.b(N137_8),.q(_w_1282));
  bfr _b_790(.a(_w_1209),.q(_w_1210));
  or_bb g221(.a(n219),.b(n220),.q(n221));
  bfr _b_1421(.a(_w_1840),.q(_w_1841));
  bfr _b_1164(.a(_w_1583),.q(_w_1584));
  bfr _b_718(.a(_w_1137),.q(N65_5));
  bfr _b_777(.a(_w_1196),.q(_w_1197));
  spl2 g369_s_0(.a(n369),.q0(n369_0),.q1(n369_1));
  or_bb g229(.a(n203_3),.b(n72_3),.q(n229));
  spl2 g298_s_1(.a(n298_1),.q0(n298_2),.q1(n298_3));
  and_bb g309(.a(N25_6),.b(n308_0),.q(n309));
  or_bb g78(.a(n76),.b(n77),.q(n78));
  bfr _b_1540(.a(_w_1959),.q(_w_1960));
  bfr _b_681(.a(_w_1100),.q(_w_1101));
  and_bi g223(.a(n218_1),.b(n221_1),.q(n223));
  bfr _b_829(.a(_w_1248),.q(_w_1249));
  bfr _b_1061(.a(_w_1480),.q(_w_1481));
  bfr _b_655(.a(_w_1074),.q(_w_1075));
  spl2 N137_s_1(.a(N137_2),.q0(N137_4),.q1(N137_5));
  or_bb g224(.a(n222),.b(n223),.q(n224));
  bfr _b_1155(.a(_w_1574),.q(_w_1575));
  or_bb g192(.a(n184_0),.b(n191_0),.q(n192));
  bfr _b_1100(.a(_w_1519),.q(_w_1520));
  and_bi g227(.a(n226),.b(n225),.q(n227));
  spl2 g233_s_1(.a(n233_1),.q0(n233_2),.q1(_w_1277));
  or_bb g247(.a(n245),.b(n246),.q(n247));
  bfr _b_874(.a(_w_1293),.q(_w_1294));
  spl2 g48_s_0(.a(n48),.q0(n48_0),.q1(n48_1));
  or_bb g259(.a(n257),.b(n258),.q(n259));
  and_bb g344(.a(n181_9),.b(n335_2),.q(n344));
  or_bb g238(.a(n209_3),.b(n78_3),.q(n238));
  spl2 g344_s_0(.a(n344),.q0(n344_0),.q1(n344_1));
  and_bi g212(.a(n78_1),.b(n209_1),.q(n212));
  spl2 g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1));
  and_bi g231(.a(n230_0),.b(n227_0),.q(n231));
  bfr _b_697(.a(_w_1116),.q(_w_1117));
  bfr _b_1024(.a(_w_1443),.q(_w_1444));
  bfr _b_781(.a(_w_1200),.q(N1_5));
  bfr _b_1067(.a(_w_1486),.q(_w_1487));
  and_bi g232(.a(n227_1),.b(n230_1),.q(n232));
  or_bb g233(.a(n231),.b(n232),.q(_w_1275));
  and_bb g304(.a(n209_6),.b(n299_1),.q(n304));
  bfr _b_1018(.a(_w_1437),.q(N745));
  or_bb g243(.a(n241),.b(n242),.q(n243));
  or_bb g177(.a(n175_1),.b(n63_3),.q(n177));
  and_bb g422(.a(N121_6),.b(n421_0),.q(n422));
  bfr _b_959(.a(_w_1378),.q(_w_1379));
  spl2 g331_s_0(.a(n331),.q0(n331_0),.q1(n331_1));
  or_bb g410(.a(N109_7),.b(n408_1),.q(n410));
  bfr _b_807(.a(_w_1226),.q(N113_2));
  or_bb g101(.a(N41_3),.b(N45_3),.q(n101));
  and_bi g260(.a(N101_3),.b(N117_3),.q(n260));
  and_bb g419(.a(N117_7),.b(n417_1),.q(n419));
  and_bi g120(.a(N77_3),.b(N93_3),.q(n120));
  or_bb g262(.a(n260),.b(n261),.q(n262));
  or_bb g97(.a(n95),.b(n96),.q(n97));
  bfr _b_656(.a(_w_1075),.q(_w_1076));
  bfr _b_1481(.a(_w_1900),.q(_w_1901));
  and_bb g263(.a(_w_1970),.b(N137_1),.q(_w_1273));
  bfr _b_657(.a(_w_1076),.q(n209_2));
  bfr _b_984(.a(_w_1403),.q(_w_1404));
  or_bb g341(.a(N53_6),.b(n340_0),.q(n341));
  bfr _b_1047(.a(_w_1466),.q(N743));
  or_bb g60(.a(n58),.b(n59),.q(n60));
  and_bi g267(.a(n263_0),.b(n266_0),.q(n267));
  spl2 g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1));
  bfr _b_1508(.a(_w_1927),.q(_w_1928));
  bfr _b_871(.a(_w_1290),.q(_w_1291));
  or_bb g109(.a(n107),.b(n108),.q(n109));
  and_bi g275(.a(n274),.b(n273),.q(n275));
  bfr _b_1299(.a(_w_1718),.q(_w_1719));
  bfr _b_1262(.a(_w_1681),.q(N751));
  spl2 g153_s_1(.a(n153_1),.q0(n153_2),.q1(n153_3));
  and_bi g104(.a(N33_0),.b(N37_0),.q(n104));
  bfr _b_646(.a(_w_1065),.q(_w_1066));
  and_bi g276(.a(n275_0),.b(n272_0),.q(n276));
  or_bb g278(.a(n276),.b(n277),.q(n278));
  and_bb g280(.a(n240_0),.b(n279_1),.q(n280));
  and_bb g281(.a(n153_2),.b(n280_0),.q(n281));
  bfr _b_1428(.a(_w_1847),.q(_w_1848));
  bfr _b_1376(.a(_w_1795),.q(n181));
  bfr _b_1039(.a(_w_1458),.q(_w_1459));
  and_bi g277(.a(n272_1),.b(n275_1),.q(n277));
  spl2 g194_s_0(.a(n194),.q0(n194_0),.q1(n194_1));
  or_bb g69(.a(n67),.b(n68),.q(n69));
  and_bb g286(.a(n209_5),.b(n281_1),.q(n286));
  spl2 g298_s_0(.a(n298),.q0(n298_0),.q1(_w_1690));
  and_bi g80(.a(N105_3),.b(N121_3),.q(n80));
  spl3L N85_s_1(.a(N85_2),.q0(N85_3),.q1(N85_4),.q2(_w_1250));
  spl2 N65_s_2(.a(N65_5),.q0(N65_6),.q1(N65_7));
  spl4L N137_s_0(.a(N137),.q0(N137_0),.q1(N137_1),.q2(N137_2),.q3(N137_3));
  spl4L g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1),.q2(n299_2),.q3(n299_3));
  spl2 N93_s_2(.a(N93_5),.q0(N93_6),.q1(N93_7));
  spl2 g85_s_0(.a(n85),.q0(n85_0),.q1(n85_1));
  bfr _b_850(.a(_w_1269),.q(_w_1270));
  spl3L N93_s_0(.a(N93),.q0(N93_0),.q1(N93_1),.q2(N93_2));
  spl3L N121_s_1(.a(N121_2),.q0(N121_3),.q1(N121_4),.q2(_w_1227));
  bfr _b_673(.a(_w_1092),.q(_w_1093));
  bfr _b_839(.a(_w_1258),.q(_w_1259));
  spl2 N121_s_2(.a(N121_5),.q0(N121_6),.q1(N121_7));
  bfr _b_641(.a(_w_1060),.q(_w_1061));
  and_bi g364(.a(n362),.b(n363),.q(_w_1674));
  spl3L N113_s_0(.a(N113),.q0(N113_0),.q1(N113_1),.q2(_w_1224));
  bfr _b_1161(.a(_w_1580),.q(_w_1581));
  spl2 g408_s_0(.a(n408),.q0(n408_0),.q1(n408_1));
  spl2 N113_s_2(.a(N113_5),.q0(N113_6),.q1(N113_7));
  bfr _b_992(.a(_w_1411),.q(_w_1412));
  bfr _b_1052(.a(_w_1471),.q(_w_1472));
  spl2 g79_s_0(.a(n79),.q0(n79_0),.q1(n79_1));
  spl3L N109_s_0(.a(N109),.q0(N109_0),.q1(N109_1),.q2(N109_2));
  spl3L N109_s_1(.a(N109_2),.q0(N109_3),.q1(N109_4),.q2(_w_1201));
  bfr _b_1494(.a(_w_1913),.q(_w_1914));
  bfr _b_1238(.a(_w_1657),.q(_w_1658));
  bfr _b_727(.a(_w_1146),.q(_w_1147));
  bfr _b_883(.a(_w_1302),.q(_w_1303));
  spl3L N1_s_1(.a(N1_2),.q0(N1_3),.q1(N1_4),.q2(_w_1177));
  spl3L N69_s_0(.a(N69),.q0(N69_0),.q1(N69_1),.q2(N69_2));
  bfr _b_851(.a(_w_1270),.q(_w_1271));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(_w_1174));
  bfr _b_845(.a(_w_1264),.q(_w_1265));
  spl3L N105_s_0(.a(N105),.q0(N105_0),.q1(N105_1),.q2(N105_2));
  or_bb g148(.a(n137_1),.b(n146_1),.q(n148));
  bfr _b_720(.a(_w_1139),.q(_w_1140));
  spl2 N105_s_2(.a(N105_5),.q0(N105_6),.q1(N105_7));
  bfr _b_1126(.a(_w_1545),.q(_w_1546));
  spl3L N101_s_0(.a(N101),.q0(N101_0),.q1(N101_1),.q2(_w_1171));
  spl2 N21_s_2(.a(N21_5),.q0(N21_6),.q1(N21_7));
  spl2 g259_s_1(.a(n259_2),.q0(n259_3),.q1(_w_1702));
  bfr _b_715(.a(_w_1134),.q(_w_1135));
  bfr _b_919(.a(_w_1338),.q(n278_4));
  bfr _b_842(.a(_w_1261),.q(_w_1262));
  spl2 g97_s_0(.a(n97),.q0(n97_0),.q1(n97_1));
  spl2 g82_s_0(.a(n82),.q0(n82_0),.q1(n82_1));
  spl2 g106_s_0(.a(n106),.q0(n106_0),.q1(n106_1));
  spl4L g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1),.q2(n109_2),.q3(n109_3));
  bfr _b_703(.a(_w_1122),.q(_w_1123));
  bfr _b_744(.a(_w_1163),.q(_w_1164));
  spl2 g197_s_0(.a(n197),.q0(n197_0),.q1(n197_1));
  spl2 g211_s_0(.a(n211),.q0(n211_0),.q1(_w_1146));
  spl2 N109_s_2(.a(N109_5),.q0(N109_6),.q1(N109_7));
  spl4L g175_s_0(.a(n175),.q0(n175_0),.q1(n175_1),.q2(n175_2),.q3(n175_3));
  spl2 N53_s_2(.a(N53_5),.q0(N53_6),.q1(N53_7));
  and_bb g348(.a(n233_11),.b(n335_3),.q(n348));
  bfr _b_876(.a(_w_1295),.q(_w_1296));
  and_bi g153(.a(n115_0),.b(n152_0),.q(n153));
  spl2 g224_s_0(.a(n224),.q0(n224_0),.q1(n224_1));
  bfr _b_1485(.a(_w_1904),.q(_w_1905));
  spl2 g184_s_0(.a(n184),.q0(n184_0),.q1(n184_1));
  spl2 g134_s_0(.a(n134),.q0(n134_0),.q1(n134_1));
  bfr _b_1368(.a(_w_1787),.q(_w_1788));
  spl3L N13_s_0(.a(N13),.q0(N13_0),.q1(N13_1),.q2(N13_2));
  bfr _b_658(.a(_w_1077),.q(_w_1078));
  spl2 N25_s_2(.a(N25_5),.q0(N25_6),.q1(N25_7));
  bfr _b_1437(.a(_w_1856),.q(_w_1857));
  spl3L g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1),.q2(_w_1145));
  spl2 g152_s_1(.a(n152_2),.q0(n152_3),.q1(_w_1138));
  and_bb g388(.a(N89_6),.b(n387_0),.q(n388));
  spl4L g152_s_2(.a(n152_4),.q0(n152_5),.q1(n152_6),.q2(n152_7),.q3(n152_8));
  spl2 g154_s_0(.a(n154),.q0(n154_0),.q1(n154_1));
  spl3L N65_s_1(.a(N65_2),.q0(N65_3),.q1(N65_4),.q2(_w_1115));
  and_bi g71(.a(n66_1),.b(n69_1),.q(n71));
  spl2 g396_s_0(.a(n396),.q0(n396_0),.q1(n396_1));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  bfr _b_1075(.a(_w_1494),.q(_w_1495));
  spl2 g160_s_0(.a(n160),.q0(n160_0),.q1(n160_1));
  spl3L N125_s_1(.a(N125_2),.q0(N125_3),.q1(N125_4),.q2(_w_1092));
  bfr _b_933(.a(_w_1352),.q(_w_1353));
  and_bi g94(.a(n92),.b(n93),.q(n94));
  bfr _b_848(.a(_w_1267),.q(_w_1268));
  bfr _b_1006(.a(_w_1425),.q(_w_1426));
  and_bi g96(.a(N5_4),.b(N1_4),.q(n96));
  spl2 N125_s_2(.a(N125_5),.q0(N125_6),.q1(N125_7));
  spl2 g178_s_0(.a(n178),.q0(n178_0),.q1(n178_1));
  bfr _b_1223(.a(_w_1642),.q(_w_1643));
  bfr _b_1062(.a(_w_1481),.q(_w_1482));
  spl2 g181_s_1(.a(n181_3),.q0(n181_4),.q1(_w_1084));
  spl4L g181_s_2(.a(n181_5),.q0(n181_6),.q1(n181_7),.q2(n181_8),.q3(n181_9));
  spl2 g290_s_0(.a(n290),.q0(n290_0),.q1(n290_1));
  spl2 g200_s_0(.a(n200),.q0(n200_0),.q1(n200_1));
  spl2 g44_s_0(.a(n44),.q0(n44_0),.q1(n44_1));
  spl4L g203_s_0(.a(n203),.q0(n203_0),.q1(n203_1),.q2(n203_2),.q3(n203_3));
  spl3L N89_s_0(.a(N89),.q0(N89_0),.q1(N89_1),.q2(N89_2));
  spl4L g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1),.q2(n63_2),.q3(n63_3));
  spl2 g115_s_1(.a(n115_2),.q0(n115_3),.q1(_w_1077));
  and_bi g386(.a(n384),.b(n385),.q(_w_1437));
  bfr _b_798(.a(_w_1217),.q(_w_1218));
  spl3L g209_s_0(.a(n209),.q0(n209_0),.q1(n209_1),.q2(_w_1074));
  bfr _b_1284(.a(_w_1703),.q(_w_1704));
  bfr _b_1252(.a(_w_1671),.q(N37_5));
  bfr _b_974(.a(_w_1393),.q(N53_2));
  spl2 g209_s_1(.a(n209_2),.q0(n209_3),.q1(_w_1067));
  spl4L g209_s_2(.a(n209_4),.q0(n209_5),.q1(n209_6),.q2(n209_7),.q3(n209_8));
  spl2 g212_s_0(.a(n212),.q0(n212_0),.q1(_w_1060));
  bfr _b_642(.a(_w_1061),.q(_w_1062));
  spl2 g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1));
  bfr _b_644(.a(_w_1063),.q(_w_1064));
  bfr _b_1066(.a(_w_1485),.q(_w_1486));
  bfr _b_648(.a(_w_1067),.q(_w_1068));
  and_bb g79(.a(_w_1971),.b(N137_4),.q(_w_1515));
  bfr _b_768(.a(_w_1187),.q(_w_1188));
  and_bi g257(.a(n256_0),.b(n253_0),.q(n257));
  bfr _b_650(.a(_w_1069),.q(_w_1070));
  bfr _b_651(.a(_w_1070),.q(_w_1071));
  bfr _b_653(.a(_w_1072),.q(_w_1073));
  bfr _b_654(.a(_w_1073),.q(n209_4));
  bfr _b_1044(.a(_w_1463),.q(_w_1464));
  bfr _b_662(.a(_w_1081),.q(_w_1082));
  bfr _b_663(.a(_w_1082),.q(_w_1083));
  bfr _b_1446(.a(_w_1865),.q(_w_1866));
  bfr _b_664(.a(_w_1083),.q(n115_4));
  bfr _b_686(.a(_w_1105),.q(_w_1106));
  bfr _b_979(.a(_w_1398),.q(_w_1399));
  bfr _b_665(.a(_w_1084),.q(_w_1085));
  spl3L N17_s_1(.a(N17_2),.q0(N17_3),.q1(N17_4),.q2(_w_1820));
  or_bb g401(.a(N101_6),.b(n400_0),.q(n401));
  bfr _b_786(.a(_w_1205),.q(_w_1206));
  bfr _b_886(.a(_w_1305),.q(_w_1306));
  bfr _b_1225(.a(_w_1644),.q(_w_1645));
  bfr _b_669(.a(_w_1088),.q(_w_1089));
  bfr _b_1096(.a(_w_1515),.q(_w_1516));
  bfr _b_670(.a(_w_1089),.q(_w_1090));
  bfr _b_1400(.a(_w_1819),.q(N41_5));
  bfr _b_891(.a(_w_1310),.q(N744));
  bfr _b_671(.a(_w_1090),.q(_w_1091));
  bfr _b_729(.a(_w_1148),.q(_w_1149));
  bfr _b_1202(.a(_w_1621),.q(_w_1622));
  and_bi g124(.a(n119_1),.b(n122_1),.q(n124));
  bfr _b_672(.a(_w_1091),.q(n181_5));
  bfr _b_675(.a(_w_1094),.q(_w_1095));
  bfr _b_661(.a(_w_1080),.q(_w_1081));
  bfr _b_676(.a(_w_1095),.q(_w_1096));
  bfr _b_678(.a(_w_1097),.q(_w_1098));
  spl3L N21_s_1(.a(N21_2),.q0(N21_3),.q1(N21_4),.q2(_w_1770));
  bfr _b_679(.a(_w_1098),.q(_w_1099));
  bfr _b_1019(.a(_w_1438),.q(_w_1439));
  or_bb g172(.a(n170),.b(n171),.q(n172));
  or_bb g48(.a(n46),.b(n47),.q(n48));
  bfr _b_938(.a(_w_1357),.q(_w_1358));
  bfr _b_682(.a(_w_1101),.q(_w_1102));
  bfr _b_683(.a(_w_1102),.q(_w_1103));
  bfr _b_1365(.a(_w_1784),.q(_w_1785));
  bfr _b_685(.a(_w_1104),.q(_w_1105));
  bfr _b_1448(.a(_w_1867),.q(N9_5));
  spl2 g66_s_0(.a(n66),.q0(n66_0),.q1(n66_1));
  bfr _b_766(.a(_w_1185),.q(_w_1186));
  bfr _b_896(.a(_w_1315),.q(_w_1316));
  bfr _b_1285(.a(_w_1704),.q(_w_1705));
  bfr _b_1038(.a(_w_1457),.q(_w_1458));
  bfr _b_687(.a(_w_1106),.q(_w_1107));
  bfr _b_689(.a(_w_1108),.q(_w_1109));
  bfr _b_694(.a(_w_1113),.q(_w_1114));
  bfr _b_699(.a(_w_1118),.q(_w_1119));
  bfr _b_1367(.a(_w_1786),.q(_w_1787));
  spl3L N1_s_0(.a(N1),.q0(N1_0),.q1(N1_1),.q2(N1_2));
  bfr _b_704(.a(_w_1123),.q(_w_1124));
  bfr _b_1326(.a(_w_1745),.q(_w_1746));
  bfr _b_1005(.a(_w_1424),.q(_w_1425));
  and_bi g230(.a(n229),.b(n228),.q(n230));
  bfr _b_707(.a(_w_1126),.q(_w_1127));
  spl2 g103_s_0(.a(n103),.q0(n103_0),.q1(n103_1));
  bfr _b_996(.a(_w_1415),.q(_w_1416));
  bfr _b_708(.a(_w_1127),.q(_w_1128));
  bfr _b_893(.a(_w_1312),.q(_w_1313));
  and_bi g303(.a(n301),.b(n302),.q(N728));
  spl2 g358_s_0(.a(n358),.q0(n358_0),.q1(n358_1));
  bfr _b_709(.a(_w_1128),.q(_w_1129));
  bfr _b_710(.a(_w_1129),.q(_w_1130));
  bfr _b_711(.a(_w_1130),.q(_w_1131));
  bfr _b_1488(.a(_w_1907),.q(_w_1908));
  bfr _b_1333(.a(_w_1752),.q(_w_1753));
  bfr _b_712(.a(_w_1131),.q(_w_1132));
  bfr _b_716(.a(_w_1135),.q(_w_1136));
  bfr _b_930(.a(_w_1349),.q(_w_1350));
  bfr _b_717(.a(_w_1136),.q(_w_1137));
  spl2 g336_s_0(.a(n336),.q0(n336_0),.q1(n336_1));
  bfr _b_721(.a(_w_1140),.q(_w_1141));
  bfr _b_1049(.a(_w_1468),.q(_w_1469));
  spl3L N45_s_0(.a(N45),.q0(N45_0),.q1(N45_1),.q2(N45_2));
  bfr _b_722(.a(_w_1141),.q(_w_1142));
  bfr _b_831(.a(_w_1250),.q(_w_1251));
  bfr _b_1008(.a(_w_1427),.q(_w_1428));
  bfr _b_723(.a(_w_1142),.q(_w_1143));
  bfr _b_724(.a(_w_1143),.q(_w_1144));
  bfr _b_1054(.a(_w_1473),.q(_w_1474));
  and_bi g159(.a(N25_1),.b(N9_1),.q(n159));
  spl2 N101_s_2(.a(N101_5),.q0(N101_6),.q1(N101_7));
  bfr _b_1022(.a(_w_1441),.q(n115_2));
  bfr _b_725(.a(_w_1144),.q(n152_4));
  bfr _b_1390(.a(_w_1809),.q(_w_1810));
  bfr _b_728(.a(_w_1147),.q(_w_1148));
  bfr _b_734(.a(_w_1153),.q(_w_1154));
  bfr _b_677(.a(_w_1096),.q(_w_1097));
  bfr _b_884(.a(_w_1303),.q(_w_1304));
  and_bi g189(.a(n185_0),.b(n188_0),.q(n189));
  bfr _b_735(.a(_w_1154),.q(_w_1155));
  and_bi g235(.a(n181_2),.b(n233_0),.q(n235));
  and_bi g149(.a(n148),.b(n147),.q(n149));
  bfr _b_738(.a(_w_1157),.q(_w_1158));
  spl3L N81_s_0(.a(N81),.q0(N81_0),.q1(N81_1),.q2(N81_2));
  bfr _b_739(.a(_w_1158),.q(_w_1159));
  bfr _b_1097(.a(_w_1516),.q(_w_1517));
  bfr _b_783(.a(_w_1202),.q(_w_1203));
  bfr _b_732(.a(_w_1151),.q(_w_1152));
  bfr _b_743(.a(_w_1162),.q(_w_1163));
  and_bi g136(.a(n131_1),.b(n134_1),.q(n136));
  bfr _b_808(.a(_w_1227),.q(_w_1228));
  bfr _b_745(.a(_w_1164),.q(_w_1165));
  bfr _b_748(.a(_w_1167),.q(_w_1168));
  bfr _b_749(.a(_w_1168),.q(_w_1169));
  bfr _b_939(.a(_w_1358),.q(_w_1359));
  or_bb g146(.a(n144),.b(n145),.q(n146));
  bfr _b_751(.a(_w_1170),.q(N101_5));
  bfr _b_785(.a(_w_1204),.q(_w_1205));
  spl4L g100_s_0(.a(n100),.q0(n100_0),.q1(n100_1),.q2(n100_2),.q3(n100_3));
  bfr _b_815(.a(_w_1234),.q(_w_1235));
  bfr _b_1055(.a(_w_1474),.q(_w_1475));
  bfr _b_752(.a(_w_1171),.q(_w_1172));
  bfr _b_753(.a(_w_1172),.q(_w_1173));
  bfr _b_779(.a(_w_1198),.q(_w_1199));
  bfr _b_755(.a(_w_1174),.q(_w_1175));
  bfr _b_756(.a(_w_1175),.q(_w_1176));
  bfr _b_757(.a(_w_1176),.q(n235_1));
  bfr _b_927(.a(_w_1346),.q(_w_1347));
  bfr _b_758(.a(_w_1177),.q(_w_1178));
  and_bi g357(.a(n355),.b(n356),.q(n357));
  bfr _b_759(.a(_w_1178),.q(_w_1179));
  spl2 g54_s_0(.a(n54),.q0(n54_0),.q1(n54_1));
  bfr _b_762(.a(_w_1181),.q(_w_1182));
  bfr _b_763(.a(_w_1182),.q(_w_1183));
  and_bi g142(.a(N53_1),.b(N49_1),.q(n142));
  bfr _b_764(.a(_w_1183),.q(_w_1184));
  bfr _b_1102(.a(_w_1521),.q(_w_1522));
  bfr _b_773(.a(_w_1192),.q(_w_1193));
  bfr _b_817(.a(_w_1236),.q(_w_1237));
  bfr _b_1009(.a(_w_1428),.q(_w_1429));
  and_bi g145(.a(n140_1),.b(n143_1),.q(n145));
  bfr _b_774(.a(_w_1193),.q(_w_1194));
  bfr _b_775(.a(_w_1194),.q(_w_1195));
  bfr _b_852(.a(_w_1271),.q(_w_1272));
  bfr _b_776(.a(_w_1195),.q(_w_1196));
  bfr _b_1016(.a(_w_1435),.q(_w_1436));
  bfr _b_1547(.a(N132),.q(_w_1967));
  bfr _b_778(.a(_w_1197),.q(_w_1198));
  bfr _b_788(.a(_w_1207),.q(_w_1208));
  and_bi g403(.a(n401),.b(n402),.q(_w_1680));
  bfr _b_789(.a(_w_1208),.q(_w_1209));
  spl3L N113_s_1(.a(N113_2),.q0(N113_3),.q1(N113_4),.q2(_w_1290));
  bfr _b_791(.a(_w_1210),.q(_w_1211));
  bfr _b_771(.a(_w_1190),.q(_w_1191));
  bfr _b_792(.a(_w_1211),.q(_w_1212));
  bfr _b_793(.a(_w_1212),.q(_w_1213));
  bfr _b_796(.a(_w_1215),.q(_w_1216));
  bfr _b_799(.a(_w_1218),.q(_w_1219));
  bfr _b_1505(.a(_w_1924),.q(_w_1925));
  bfr _b_947(.a(_w_1366),.q(_w_1367));
  bfr _b_977(.a(_w_1396),.q(_w_1397));
  bfr _b_1026(.a(_w_1445),.q(_w_1446));
  bfr _b_800(.a(_w_1219),.q(_w_1220));
  bfr _b_801(.a(_w_1220),.q(_w_1221));
  bfr _b_802(.a(_w_1221),.q(_w_1222));
  bfr _b_952(.a(_w_1371),.q(_w_1372));
  bfr _b_803(.a(_w_1222),.q(_w_1223));
  bfr _b_804(.a(_w_1223),.q(N109_5));
  bfr _b_806(.a(_w_1225),.q(_w_1226));
  bfr _b_809(.a(_w_1228),.q(_w_1229));
  bfr _b_1308(.a(_w_1727),.q(_w_1728));
  spl4L g181_s_0(.a(n181),.q0(n181_0),.q1(n181_1),.q2(n181_2),.q3(n181_3));
  bfr _b_810(.a(_w_1229),.q(_w_1230));
  bfr _b_811(.a(_w_1230),.q(_w_1231));
  bfr _b_826(.a(_w_1245),.q(_w_1246));
  bfr _b_812(.a(_w_1231),.q(_w_1232));
  bfr _b_1511(.a(_w_1930),.q(_w_1931));
  bfr _b_816(.a(_w_1235),.q(_w_1236));
  bfr _b_821(.a(_w_1240),.q(_w_1241));
  bfr _b_823(.a(_w_1242),.q(_w_1243));
  and_bi g411(.a(n410),.b(n409),.q(_w_1681));
  bfr _b_825(.a(_w_1244),.q(_w_1245));
  bfr _b_827(.a(_w_1246),.q(_w_1247));
  bfr _b_649(.a(_w_1068),.q(_w_1069));
  and_bi g98(.a(n97_0),.b(n94_0),.q(n98));
  bfr _b_828(.a(_w_1247),.q(_w_1248));
  bfr _b_953(.a(_w_1372),.q(_w_1373));
  bfr _b_830(.a(_w_1249),.q(N121_5));
  bfr _b_742(.a(_w_1161),.q(_w_1162));
  bfr _b_935(.a(_w_1354),.q(_w_1355));
  spl2 N49_s_2(.a(N49_5),.q0(N49_6),.q1(N49_7));
  bfr _b_833(.a(_w_1252),.q(_w_1253));
  bfr _b_674(.a(_w_1093),.q(_w_1094));
  bfr _b_834(.a(_w_1253),.q(_w_1254));
  bfr _b_1208(.a(_w_1627),.q(_w_1628));
  and_bi g351(.a(n350),.b(n349),.q(N739));
  bfr _b_835(.a(_w_1254),.q(_w_1255));
  bfr _b_837(.a(_w_1256),.q(_w_1257));
  spl3L N97_s_1(.a(N97_2),.q0(N97_3),.q1(N97_4),.q2(_w_1311));
  bfr _b_846(.a(_w_1265),.q(_w_1266));
  bfr _b_968(.a(_w_1387),.q(_w_1388));
  bfr _b_991(.a(_w_1410),.q(_w_1411));
  spl3L N25_s_1(.a(N25_2),.q0(N25_3),.q1(N25_4),.q2(_w_1340));
  bfr _b_840(.a(_w_1259),.q(_w_1260));
  bfr _b_841(.a(_w_1260),.q(_w_1261));
  bfr _b_1411(.a(_w_1830),.q(_w_1831));
  bfr _b_843(.a(_w_1262),.q(_w_1263));
  or_bb g181(.a(n179),.b(n180),.q(_w_1794));
  bfr _b_645(.a(_w_1064),.q(_w_1065));
  bfr _b_667(.a(_w_1086),.q(_w_1087));
  bfr _b_847(.a(_w_1266),.q(_w_1267));
  bfr _b_1041(.a(_w_1460),.q(_w_1461));
  spl3L N17_s_0(.a(N17),.q0(N17_0),.q1(N17_1),.q2(N17_2));
  bfr _b_854(.a(_w_1273),.q(_w_1274));
  and_bi g68(.a(N85_1),.b(N81_1),.q(n68));
  bfr _b_855(.a(_w_1274),.q(n263));
  bfr _b_857(.a(_w_1276),.q(n233));
  bfr _b_860(.a(_w_1279),.q(_w_1280));
  bfr _b_862(.a(_w_1281),.q(n116));
  bfr _b_864(.a(_w_1283),.q(_w_1284));
  bfr _b_693(.a(_w_1112),.q(_w_1113));
  bfr _b_1069(.a(_w_1488),.q(N33_5));
  bfr _b_865(.a(_w_1284),.q(n215));
  bfr _b_866(.a(_w_1285),.q(_w_1286));
  bfr _b_1538(.a(_w_1957),.q(_w_1958));
  bfr _b_868(.a(_w_1287),.q(_w_1288));
  and_bi g293(.a(n292),.b(n291),.q(N726));
  or_bb g51(.a(n49),.b(n50),.q(n51));
  bfr _b_869(.a(_w_1288),.q(_w_1289));
  bfr _b_870(.a(_w_1289),.q(n213_1));
  bfr _b_1261(.a(_w_1680),.q(N749));
  bfr _b_872(.a(_w_1291),.q(_w_1292));
  bfr _b_1478(.a(_w_1897),.q(_w_1898));
  bfr _b_877(.a(_w_1296),.q(_w_1297));
  bfr _b_719(.a(_w_1138),.q(_w_1139));
  bfr _b_878(.a(_w_1297),.q(_w_1298));
  bfr _b_879(.a(_w_1298),.q(_w_1299));
  bfr _b_885(.a(_w_1304),.q(_w_1305));
  bfr _b_887(.a(_w_1306),.q(_w_1307));
  bfr _b_888(.a(_w_1307),.q(_w_1308));
  bfr _b_1031(.a(_w_1450),.q(_w_1451));
  bfr _b_1383(.a(_w_1802),.q(_w_1803));
  and_bi g416(.a(n414),.b(n415),.q(_w_1682));
  and_bi g87(.a(n82_1),.b(n85_1),.q(n87));
  bfr _b_892(.a(_w_1311),.q(_w_1312));
  bfr _b_925(.a(_w_1344),.q(_w_1345));
  bfr _b_1003(.a(_w_1422),.q(_w_1423));
  bfr _b_894(.a(_w_1313),.q(_w_1314));
  bfr _b_1469(.a(_w_1888),.q(_w_1889));
  bfr _b_705(.a(_w_1124),.q(_w_1125));
  bfr _b_895(.a(_w_1314),.q(_w_1315));
  bfr _b_897(.a(_w_1316),.q(_w_1317));
  bfr _b_901(.a(_w_1320),.q(_w_1321));
  bfr _b_1315(.a(_w_1734),.q(_w_1735));
  bfr _b_902(.a(_w_1321),.q(_w_1322));
  and_bi g81(.a(N121_4),.b(N105_4),.q(n81));
  bfr _b_903(.a(_w_1322),.q(_w_1323));
  bfr _b_904(.a(_w_1323),.q(_w_1324));
  bfr _b_905(.a(_w_1324),.q(_w_1325));
  bfr _b_1346(.a(_w_1765),.q(_w_1766));
  bfr _b_906(.a(_w_1325),.q(_w_1326));
  spl2 g60_s_0(.a(n60),.q0(n60_0),.q1(n60_1));
  bfr _b_907(.a(_w_1326),.q(_w_1327));
  bfr _b_889(.a(_w_1308),.q(_w_1309));
  bfr _b_909(.a(_w_1328),.q(_w_1329));
  bfr _b_1105(.a(_w_1524),.q(_w_1525));
  bfr _b_972(.a(_w_1391),.q(_w_1392));
  spl4L g281_s_0(.a(n281),.q0(n281_0),.q1(n281_1),.q2(n281_2),.q3(n281_3));
  bfr _b_741(.a(_w_1160),.q(_w_1161));
  bfr _b_910(.a(_w_1329),.q(_w_1330));
  bfr _b_911(.a(_w_1330),.q(N97_5));
  or_bb g266(.a(n264),.b(n265),.q(n266));
  bfr _b_913(.a(_w_1332),.q(_w_1333));
  spl2 N1_s_2(.a(N1_5),.q0(N1_6),.q1(N1_7));
  bfr _b_916(.a(_w_1335),.q(_w_1336));
  bfr _b_917(.a(_w_1336),.q(_w_1337));
  bfr _b_918(.a(_w_1337),.q(_w_1338));
  bfr _b_920(.a(_w_1339),.q(n244));
  and_bi g279(.a(n259_0),.b(n278_0),.q(n279));
  spl2 g319_s_0(.a(n319),.q0(n319_0),.q1(n319_1));
  bfr _b_921(.a(_w_1340),.q(_w_1341));
  bfr _b_923(.a(_w_1342),.q(_w_1343));
  bfr _b_1182(.a(_w_1601),.q(_w_1602));
  bfr _b_929(.a(_w_1348),.q(_w_1349));
  bfr _b_1492(.a(_w_1911),.q(_w_1912));
  bfr _b_1392(.a(_w_1811),.q(_w_1812));
  and_bb g323(.a(n209_7),.b(n318_1),.q(n323));
  bfr _b_931(.a(_w_1350),.q(_w_1351));
  bfr _b_937(.a(_w_1356),.q(_w_1357));
  bfr _b_941(.a(_w_1360),.q(_w_1361));
  bfr _b_945(.a(_w_1364),.q(_w_1365));
  bfr _b_1382(.a(_w_1801),.q(_w_1802));
  bfr _b_948(.a(_w_1367),.q(_w_1368));
  bfr _b_949(.a(_w_1368),.q(_w_1369));
  bfr _b_950(.a(_w_1369),.q(_w_1370));
  bfr _b_973(.a(_w_1392),.q(n153_1));
  bfr _b_951(.a(_w_1370),.q(_w_1371));
  bfr _b_955(.a(_w_1374),.q(_w_1375));
  bfr _b_761(.a(_w_1180),.q(_w_1181));
  bfr _b_975(.a(_w_1394),.q(_w_1395));
  bfr _b_1015(.a(_w_1434),.q(_w_1435));
  bfr _b_956(.a(_w_1375),.q(_w_1376));
  bfr _b_958(.a(_w_1377),.q(_w_1378));
  bfr _b_1209(.a(_w_1628),.q(_w_1629));
  bfr _b_960(.a(_w_1379),.q(_w_1380));
  bfr _b_961(.a(_w_1380),.q(_w_1381));
  bfr _b_1353(.a(_w_1772),.q(_w_1773));
  bfr _b_962(.a(_w_1381),.q(_w_1382));
  bfr _b_963(.a(_w_1382),.q(_w_1383));
  and_bi g54(.a(n52),.b(n53),.q(n54));
  bfr _b_965(.a(_w_1384),.q(_w_1385));
  bfr _b_971(.a(_w_1390),.q(_w_1391));
  or_bb g205(.a(n175_3),.b(n203_1),.q(n205));
  bfr _b_966(.a(_w_1385),.q(_w_1386));
  bfr _b_969(.a(_w_1388),.q(_w_1389));
  bfr _b_980(.a(_w_1399),.q(_w_1400));
  bfr _b_982(.a(_w_1401),.q(_w_1402));
  bfr _b_983(.a(_w_1402),.q(_w_1403));
  bfr _b_1197(.a(_w_1616),.q(_w_1617));
  or_bb g362(.a(N65_6),.b(n361_0),.q(n362));
  bfr _b_985(.a(_w_1404),.q(_w_1405));
  bfr _b_736(.a(_w_1155),.q(_w_1156));
  bfr _b_987(.a(_w_1406),.q(_w_1407));
  spl3L N101_s_1(.a(N101_2),.q0(N101_3),.q1(N101_4),.q2(_w_1151));
  bfr _b_989(.a(_w_1408),.q(_w_1409));
  spl3L N61_s_0(.a(N61),.q0(N61_0),.q1(N61_1),.q2(N61_2));
  bfr _b_993(.a(_w_1412),.q(_w_1413));
  bfr _b_1001(.a(_w_1420),.q(_w_1421));
  bfr _b_994(.a(_w_1413),.q(N117_5));
  bfr _b_995(.a(_w_1414),.q(_w_1415));
  spl3L N61_s_1(.a(N61_2),.q0(N61_3),.q1(N61_4),.q2(_w_1626));
  bfr _b_997(.a(_w_1416),.q(_w_1417));
  or_bb g44(.a(n42),.b(n43),.q(n44));
  bfr _b_998(.a(_w_1417),.q(_w_1418));
  bfr _b_1002(.a(_w_1421),.q(_w_1422));
  bfr _b_1004(.a(_w_1423),.q(_w_1424));
  bfr _b_1007(.a(_w_1426),.q(_w_1427));
  bfr _b_1010(.a(_w_1429),.q(_w_1430));
  bfr _b_986(.a(_w_1405),.q(_w_1406));
  bfr _b_1011(.a(_w_1430),.q(_w_1431));
  bfr _b_1487(.a(_w_1906),.q(_w_1907));
  bfr _b_1012(.a(_w_1431),.q(_w_1432));
  bfr _b_1013(.a(_w_1432),.q(_w_1433));
  bfr _b_1486(.a(_w_1905),.q(_w_1906));
  bfr _b_1014(.a(_w_1433),.q(_w_1434));
  bfr _b_1331(.a(_w_1750),.q(_w_1751));
  and_bi g239(.a(n237),.b(n238),.q(n239));
  bfr _b_946(.a(_w_1365),.q(_w_1366));
  bfr _b_1017(.a(_w_1436),.q(N93_5));
  bfr _b_1020(.a(_w_1439),.q(_w_1440));
  bfr _b_1021(.a(_w_1440),.q(n78_2));
  bfr _b_1030(.a(_w_1449),.q(_w_1450));
  and_bb g284(.a(N1_7),.b(n282_1),.q(n284));
  bfr _b_1032(.a(_w_1451),.q(_w_1452));
  bfr _b_1034(.a(_w_1453),.q(_w_1454));
  bfr _b_1036(.a(_w_1455),.q(_w_1456));
  bfr _b_1037(.a(_w_1456),.q(_w_1457));
  bfr _b_680(.a(_w_1099),.q(_w_1100));
  spl3L N33_s_0(.a(_w_1975),.q0(N33_0),.q1(N33_1),.q2(_w_1679));
  bfr _b_1046(.a(_w_1465),.q(N13_5));
  bfr _b_1476(.a(_w_1895),.q(_w_1896));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(n280_1));
  bfr _b_1048(.a(_w_1467),.q(_w_1468));
  bfr _b_822(.a(_w_1241),.q(_w_1242));
  bfr _b_1050(.a(_w_1469),.q(_w_1470));
  bfr _b_1452(.a(_w_1871),.q(_w_1872));
  bfr _b_1051(.a(_w_1470),.q(_w_1471));
  spl2 N17_s_2(.a(N17_5),.q0(N17_6),.q1(N17_7));
  and_bb g139(.a(N57_4),.b(N61_4),.q(n139));
  bfr _b_954(.a(_w_1373),.q(_w_1374));
  bfr _b_936(.a(_w_1355),.q(_w_1356));
  bfr _b_1053(.a(_w_1472),.q(_w_1473));
  bfr _b_1435(.a(_w_1854),.q(_w_1855));
  and_bi g133(.a(N21_4),.b(N17_4),.q(n133));
  bfr _b_1057(.a(_w_1476),.q(_w_1477));
  bfr _b_1296(.a(_w_1715),.q(n78_4));
  spl4L g378_s_0(.a(n378),.q0(n378_0),.q1(n378_1),.q2(n378_2),.q3(n378_3));
  bfr _b_1058(.a(_w_1477),.q(_w_1478));
  bfr _b_1185(.a(_w_1604),.q(_w_1605));
  bfr _b_1059(.a(_w_1478),.q(_w_1479));
  bfr _b_1060(.a(_w_1479),.q(_w_1480));
  bfr _b_1064(.a(_w_1483),.q(_w_1484));
  bfr _b_1065(.a(_w_1484),.q(_w_1485));
  bfr _b_978(.a(_w_1397),.q(_w_1398));
  bfr _b_1107(.a(_w_1526),.q(_w_1527));
  bfr _b_1070(.a(_w_1489),.q(n45));
  bfr _b_1072(.a(_w_1491),.q(_w_1492));
  bfr _b_1184(.a(_w_1603),.q(n210_1));
  bfr _b_1074(.a(_w_1493),.q(_w_1494));
  bfr _b_1076(.a(_w_1495),.q(_w_1496));
  bfr _b_1438(.a(_w_1857),.q(_w_1858));
  bfr _b_1078(.a(_w_1497),.q(_w_1498));
  bfr _b_881(.a(_w_1300),.q(_w_1301));
  bfr _b_1080(.a(_w_1499),.q(_w_1500));
  bfr _b_1081(.a(_w_1500),.q(_w_1501));
  bfr _b_1084(.a(_w_1503),.q(_w_1504));
  bfr _b_1088(.a(_w_1507),.q(_w_1508));
  bfr _b_805(.a(_w_1224),.q(_w_1225));
  bfr _b_1089(.a(_w_1508),.q(_w_1509));
  bfr _b_1090(.a(_w_1509),.q(_w_1510));
  bfr _b_1093(.a(_w_1512),.q(_w_1513));
  bfr _b_1094(.a(_w_1513),.q(_w_1514));
  bfr _b_900(.a(_w_1319),.q(_w_1320));
  bfr _b_819(.a(_w_1238),.q(_w_1239));
  bfr _b_1095(.a(_w_1514),.q(N45_5));
  bfr _b_1099(.a(_w_1518),.q(n79));
  bfr _b_1101(.a(_w_1520),.q(_w_1521));
  bfr _b_1104(.a(_w_1523),.q(_w_1524));
  bfr _b_1558(.a(N49),.q(_w_1977));
  bfr _b_1108(.a(_w_1527),.q(_w_1528));
endmodule
