module c432 (N1,N102,N105,N108,N11,N112,N115,N14,N17,N21,N24,N27,N30,N34,N37,N4,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N8,N82,N86,N89,N92,N95,N99,N223,N329,N370,N421,N430,N431,N432);
  input N1,N102,N105,N108,N11,N112,N115,N14,N17,N21,N24,N27,N30,N34,N37,N4,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N8,N82,N86,N89,N92,N95,N99;
  output N223,N329,N370,N421,N430,N431,N432;
  wire _w_1236,_w_1235,_w_1234,_w_1233,_w_1229,_w_1228,_w_1226,_w_1224,_w_1223,_w_1222,_w_1221,_w_1220,_w_1217,_w_1215,_w_1214,_w_1213,_w_1211,_w_1210,_w_1208,_w_1206,_w_1204,_w_1203,_w_1202,_w_1201,_w_1200,_w_1197,_w_1196,_w_1194,_w_1193,_w_1191,_w_1190,_w_1186,_w_1184,_w_1219,_w_1183,_w_1182,_w_1179,_w_1177,_w_1176,_w_1175,_w_1174,_w_1173,_w_1171,_w_1166,_w_1164,_w_1163,_w_1162,_w_1161,_w_1159,_w_1158,_w_1156,_w_1155,_w_1154,_w_1153,_w_1151,_w_1150,_w_1148,_w_1146,_w_1145,_w_1144,_w_1141,_w_1139,_w_1134,_w_1133,_w_1131,_w_1130,_w_1129,_w_1127,_w_1126,_w_1122,_w_1120,_w_1119,_w_1114,_w_1113,_w_1112,_w_1111,N21_3,N34_0,N69_2,N69_1,N27_1,n62_0,_w_855,_w_943,N30_2,N37_1,n38_3,n55_8,_w_1185,_w_1057,N43_0,N47_3,_w_622,_w_921,N47_1,_w_769,N56_3,N56_1,N60_0,N8_2,_w_638,_w_722,N73_3,N73_0,_w_1232,_w_660,_w_1216,_w_1115,N76_0,n168_0,n173,_w_1181,_w_828,n120_0,N112_2,N21_0,_w_793,N82_0,_w_623,N86_3,N86_1,N430_1,N92_0,N95_0,n77_3,_w_1096,N50_0,_w_732,_w_1100,N99_0,N329_11,N329_10,N99_2,n112_0,_w_659,N329_9,n68,N66_1,N329_2,N370_11,_w_700,N370_6,n176,_w_813,n77_4,n39_0,n100_1,_w_583,N370_7,n40_3,n151_0,n40_0,n50_3,n50_0,n51_3,_w_1081,n51_2,n41,n51_1,_w_780,_w_992,_w_1105,n51_0,n95_1,n41_0,n164_3,n130_0,n45_2,_w_571,n46_1,_w_723,n49_6,n41_3,_w_691,n52_4,n46_3,n52_1,n117_3,_w_632,n68_0,_w_1063,n55_11,n55_5,n55_2,_w_670,n55_0,n56_1,_w_953,n57_1,n57_0,_w_833,N56_0,n58_6,n82_4,n58_2,_w_697,n72_0,_w_1070,n192_1,N4_0,n192_0,N4_3,n174_0,n96_1,_w_1058,n156_1,n82_6,n37_0,n146,N43_1,_w_586,N115_0,N105_1,n144,N99_1,N50_1,n82_1,_w_616,n82_0,_w_942,n50_1,n103,n87_0,_w_867,n89_4,N43_3,n80,_w_820,n104_0,n132_1,n194,n108_4,n108_3,n184,_w_669,_w_885,n108_1,n82_3,n142,n186_1,N4_1,_w_763,n186_0,n109_0,n112_1,n55,N21_1,_w_738,n170_0,n49_3,N4_5,_w_680,_w_1073,N95_3,_w_854,n117_0,n174_1,n197_1,n58_9,n120_1,n56_0,_w_847,n138_0,_w_619,n49_1,n198,_w_653,_w_818,_w_1045,n195_1,n126_0,_w_852,_w_600,_w_860,n164_2,n197,n124,_w_948,n93_2,n55_4,n174,n55_1,n111,_w_628,_w_772,_w_634,n40_1,n208,n164,_w_936,n159,N34_1,_w_1199,_w_666,n46_2,_w_578,n89_3,_w_880,_w_816,n49_5,_w_916,N27_0,n135,n55_6,N56_2,_w_814,n172,n40_2,_w_1091,n168,n204,_w_719,N370_1,n153,_w_737,N329_8,n207,n155_3,n42_1,_w_838,n140_0,n61,_w_884,n95_0,_w_597,n108_2,n82_5,_w_654,n117_2,n165,N105_0,n77,N30_0,_w_996,_w_753,_w_1121,_w_767,_w_889,n210,n58_5,_w_1180,N99_3,_w_857,N24_0,n183,n93_3,n187,n44_0,n37,n58_4,n117,n94,_w_1128,_w_841,_w_1032,N47_0,_w_756,n178_0,n96_0,_w_913,n40,n37_2,n47_0,_w_730,n50,n67,_w_1118,n45_1,_w_810,n51,n59,n171_0,n42,n191_1,_w_598,_w_1048,n43,n87_5,n37_1,n118,n46,n47,N4_4,_w_1067,_w_1137,N34_2,_w_1076,n144_1,n49,n52,n83,n54,_w_897,n195,_w_726,n189_0,_w_792,n56,N370_5,n87_4,N79_0,n57,n72_1,_w_733,n132,n196,n58,n60,n64,n87_1,_w_1087,_w_1147,n44_1,n65,N82_2,_w_589,n69,n143,_w_1061,n191_0,_w_1037,_w_1010,_w_1110,n71,N92_1,n72,N60_3,_w_807,n38_1,n52_3,n108_5,n48,_w_808,_w_1079,_w_752,_w_1195,n79,n73_1,n96,n156,n156_0,n181_1,n87_6,n82,N95_2,n174_2,n170,n85,N73_2,n155_4,_w_773,_w_802,N69_3,_w_1011,N76_1,_w_648,n86,n76,N115_1,n87,n88,n89,n109_1,n58_8,n90,_w_1192,n113,n169,_w_576,n91,N329_6,N37_0,_w_626,n99,n195_0,_w_1005,_w_971,_w_1093,n102,N60_1,_w_1089,_w_720,n101,_w_630,_w_1140,_w_764,N21_2,_w_1012,_w_1025,_w_805,_w_1054,n68_1,n105,_w_636,n163,_w_825,_w_862,n180_3,_w_1075,_w_599,n138_1,n77_0,n89_0,_w_804,_w_688,_w_1062,n108,n109,n110,_w_1001,N370_8,n186,_w_871,n112,N370_9,n58_7,n52_6,_w_735,n114,N1_0,n116,N329_1,n55_7,n84,n144_0,n52_5,n136,_w_642,_w_950,_w_1143,n52_0,n87_2,n122,_w_715,n105_1,n123,n149,n49_4,N43_2,n130_1,n168_1,n55_3,_w_827,n41_2,n74,n49_0,n78,N30_1,_w_849,N60_2,_w_944,n181_3,_w_878,_w_675,_w_1123,n58_11,_w_912,_w_1142,n103_1,_w_1078,_w_1077,_w_1099,_w_1205,_w_1198,n47_1,n128,n50_2,n125,_w_1085,n130,_w_591,N47_2,n121_1,N329_7,_w_822,n121,_w_1097,n131,n75,_w_1047,N4_2,n133,N370_3,n105_0,n134,_w_922,_w_711,n138,n52_2,n126_1,_w_1027,_w_1135,n41_1,n139,_w_1136,n63_1,_w_993,N53_0,n140,_w_679,n104,_w_624,n141,_w_928,n104_1,_w_1064,n189_1,n147,_w_977,n63,n148,n202,_w_896,_w_682,_w_899,_w_1152,_w_667,n37_3,_w_698,n58_1,n151,_w_678,n42_0,n98,_w_746,_w_761,n154,n178,N329_3,N329_5,n157,n170_1,n193,n160,N66_0,_w_635,_w_927,n162,_w_1095,N95_1,n166,N370_2,n117_1,n171,n46_0,n177,_w_1167,n188_1,n167_0,n155,n180,n137_1,_w_749,N329_4,n152,N329_0,n99_0,n100_0,n87_3,N82_3,n73,_w_904,n108_0,n188,n200,n49_2,_w_972,n77_2,N8_1,N8_3,_w_681,_w_1084,_w_907,n70,_w_935,n190,N73_1,n140_1,n191,N370_0,n129,n44,n192,n201,_w_982,n39_1,n181_2,_w_798,n115,_w_610,_w_973,_w_980,n151_1,_w_1157,N69_0,N34_4,n209,_w_1023,N30_4,N430_0,n180_0,_w_674,n181_0,n100,n180_1,N82_1,_w_594,n99_1,_w_895,n38_2,n164_0,n155_1,n155_5,n45_0,n89_1,n164_1,_w_1189,_w_1042,n185,n188_0,n137_0,n175_1,_w_868,n146_1,n62,_w_811,n132_0,N17_0,n146_0,_w_713,N17_2,n55_10,_w_1052,n93_0,N17_3,_w_1172,_w_1071,N14_0,_w_748,n175,_w_740,_w_1138,N34_5,N112_1,N11_0,_w_1124,_w_924,n120,N11_1,N108_0,_w_1065,N108_2,_w_585,N108_3,N102_0,N102_1,_w_762,_w_861,N1_1,N1_3,_w_790,_w_568,N108_1,_w_613,_w_570,N86_0,_w_572,_w_573,_w_796,_w_1169,_w_574,_w_1116,_w_1050,_w_575,_w_580,n69_1,n103_0,_w_900,n81,_w_582,_w_584,_w_937,n127,_w_587,_w_588,_w_590,n58_3,N17_1,_w_592,_w_593,_w_887,_w_596,_w_1039,_w_1178,n181,_w_602,_w_1168,_w_835,N14_1,_w_850,_w_604,n137,_w_607,n175_0,_w_608,n93_1,_w_611,_w_891,_w_612,_w_614,_w_615,_w_617,_w_1117,_w_618,_w_620,_w_625,_w_629,_w_966,_w_631,n45_3,_w_633,n197_0,_w_725,_w_846,_w_637,_w_983,_w_640,_w_851,_w_643,n178_1,_w_989,_w_751,_w_645,_w_882,n158,_w_646,_w_803,N112_0,_w_647,_w_834,_w_649,_w_1187,_w_651,_w_741,_w_952,_w_1101,_w_655,_w_843,_w_829,_w_656,N112_3,_w_997,_w_657,_w_658,_w_661,_w_662,_w_663,_w_664,_w_754,_w_665,_w_799,_w_668,_w_603,_w_671,_w_673,N24_1,_w_1102,_w_676,_w_677,_w_683,n73_0,_w_684,_w_1149,_w_750,_w_1021,n63_0,_w_685,_w_689,_w_696,_w_692,n58_10,_w_693,_w_601,_w_859,_w_694,_w_695,_w_699,_w_701,_w_702,_w_704,_w_939,_w_705,n167,_w_1060,_w_902,_w_706,_w_707,n155_0,_w_708,_w_1002,_w_709,_w_710,_w_712,_w_714,_w_1033,n189,_w_716,_w_718,_w_863,_w_721,_w_1104,_w_842,_w_1000,_w_724,n179,_w_1036,_w_569,_w_839,_w_728,_w_729,n145,_w_731,_w_734,_w_639,n93,_w_736,_w_1038,n89_2,_w_742,_w_743,n121_0,_w_845,_w_745,_w_747,_w_1046,_w_757,_w_758,_w_765,_w_1008,_w_1098,_w_766,_w_768,_w_844,n92,_w_770,_w_771,_w_774,_w_775,_w_776,_w_777,_w_778,_w_941,N79_1,_w_781,N34_3,_w_903,_w_1230,_w_782,n199,_w_783,_w_1231,n39,n167_1,_w_785,_w_786,_w_788,_w_791,_w_1034,_w_794,_w_956,_w_760,_w_1056,_w_795,_w_652,_w_934,N370_10,_w_797,N8_0,_w_806,_w_801,_w_809,_w_1132,_w_755,_w_812,_w_779,_w_962,_w_815,_w_817,_w_821,n119,_w_932,n97,n66,_w_831,_w_836,_w_837,_w_840,_w_848,N86_2,_w_853,_w_856,_w_605,_w_858,_w_864,_w_1019,_w_865,_w_869,_w_1209,_w_717,_w_872,_w_870,_w_873,_w_1006,_w_874,_w_875,_w_876,_w_931,_w_1170,_w_1044,_w_866,_w_877,_w_879,_w_881,_w_883,_w_886,_w_888,_w_577,_w_890,n55_9,_w_832,_w_892,_w_581,_w_893,_w_579,_w_894,_w_898,n150,_w_901,_w_990,_w_905,n58_0,_w_906,_w_1109,_w_595,_w_739,_w_908,_w_976,n82_2,_w_909,_w_910,_w_1082,_w_823,_w_672,_w_911,n38,_w_914,_w_915,n82_7,_w_819,_w_917,_w_918,_w_789,_w_919,_w_826,_w_920,_w_1009,_w_923,_w_925,_w_926,_w_929,_w_930,_w_787,_w_824,_w_933,_w_938,n206,_w_621,_w_1094,n126,_w_940,_w_951,_w_627,_w_945,_w_644,_w_946,_w_947,_w_609,_w_949,_w_954,_w_641,_w_800,_w_955,_w_957,n45,_w_958,_w_1212,_w_690,_w_959,_w_960,n107,_w_961,_w_963,_w_994,N30_3,_w_964,_w_965,_w_967,n62_1,_w_968,_w_1225,_w_969,_w_970,_w_1207,_w_974,_w_975,_w_978,_w_1227,_w_998,_w_1125,_w_979,_w_981,_w_984,_w_985,_w_1160,_w_1024,N53_1,_w_986,_w_650,_w_987,_w_988,n38_0,_w_991,_w_995,_w_999,_w_784,_w_1003,_w_1090,_w_1004,_w_1007,_w_1013,_w_1014,_w_1015,_w_1165,_w_1016,N370_4,_w_1017,n77_1,_w_687,_w_1018,n171_1,_w_1020,_w_1022,_w_1026,n155_2,_w_1028,_w_1029,_w_1030,_w_1031,_w_1040,_w_1035,_w_1041,_w_1043,_w_1049,_w_686,_w_1051,_w_1053,_w_1055,_w_1059,_w_1066,_w_606,_w_1068,_w_703,_w_744,_w_727,_w_1069,_w_1072,N1_2,n69_0,_w_1074,_w_1080,_w_1218,_w_759,_w_830,_w_1083,n95,_w_1086,_w_1088,_w_1188,_w_1092,_w_1103,n180_2,_w_1106,_w_1107,_w_1108;

  bfr _b_1004(.a(_w_1236),.q(_w_1228));
  bfr _b_1002(.a(_w_1234),.q(_w_1235));
  bfr _b_1001(.a(_w_1233),.q(_w_1234));
  bfr _b_997(.a(_w_1229),.q(_w_1230));
  bfr _b_995(.a(_w_1227),.q(_w_1214));
  bfr _b_993(.a(_w_1225),.q(_w_1226));
  bfr _b_992(.a(_w_1224),.q(_w_1225));
  bfr _b_989(.a(_w_1221),.q(_w_1222));
  bfr _b_987(.a(_w_1219),.q(_w_1220));
  bfr _b_985(.a(_w_1217),.q(_w_1218));
  bfr _b_983(.a(_w_1215),.q(_w_1216));
  bfr _b_980(.a(_w_1212),.q(_w_1210));
  bfr _b_978(.a(N86),.q(_w_1211));
  bfr _b_976(.a(_w_1208),.q(_w_1209));
  bfr _b_974(.a(_w_1206),.q(_w_1207));
  bfr _b_972(.a(_w_1204),.q(_w_1205));
  bfr _b_969(.a(N8),.q(_w_1202));
  bfr _b_966(.a(_w_1198),.q(_w_1199));
  bfr _b_964(.a(_w_1196),.q(_w_1197));
  bfr _b_963(.a(_w_1195),.q(_w_1196));
  bfr _b_962(.a(_w_1194),.q(_w_1195));
  bfr _b_961(.a(_w_1193),.q(_w_1194));
  bfr _b_960(.a(_w_1192),.q(_w_1193));
  bfr _b_958(.a(_w_1190),.q(_w_1191));
  bfr _b_956(.a(_w_1188),.q(_w_1189));
  bfr _b_975(.a(_w_1207),.q(_w_1208));
  bfr _b_955(.a(N79),.q(_w_1188));
  bfr _b_951(.a(_w_1183),.q(_w_1184));
  bfr _b_973(.a(_w_1205),.q(_w_1206));
  bfr _b_950(.a(_w_1182),.q(_w_1183));
  bfr _b_949(.a(_w_1181),.q(_w_1182));
  bfr _b_948(.a(_w_1180),.q(_w_1181));
  bfr _b_946(.a(N73),.q(_w_1179));
  bfr _b_945(.a(_w_1177),.q(_w_1163));
  bfr _b_970(.a(_w_1202),.q(_w_1203));
  bfr _b_944(.a(_w_1176),.q(_w_1177));
  bfr _b_942(.a(_w_1174),.q(_w_1175));
  bfr _b_941(.a(_w_1173),.q(_w_1174));
  bfr _b_937(.a(_w_1169),.q(_w_1170));
  bfr _b_936(.a(_w_1168),.q(_w_1169));
  bfr _b_934(.a(_w_1166),.q(_w_1167));
  bfr _b_933(.a(_w_1165),.q(_w_1166));
  bfr _b_931(.a(N66),.q(_w_1164));
  bfr _b_930(.a(N63),.q(_w_1162));
  bfr _b_929(.a(_w_1161),.q(_w_1160));
  bfr _b_923(.a(_w_1155),.q(_w_1156));
  bfr _b_920(.a(_w_1152),.q(_w_1153));
  bfr _b_918(.a(_w_1150),.q(_w_1151));
  bfr _b_916(.a(_w_1148),.q(_w_1149));
  bfr _b_915(.a(_w_1147),.q(_w_1148));
  bfr _b_914(.a(_w_1146),.q(_w_1147));
  bfr _b_912(.a(_w_1144),.q(_w_1143));
  bfr _b_913(.a(N53),.q(_w_1146));
  bfr _b_911(.a(N47),.q(_w_1144));
  bfr _b_909(.a(_w_1141),.q(_w_1142));
  bfr _b_906(.a(_w_1138),.q(_w_1139));
  bfr _b_905(.a(_w_1137),.q(_w_1138));
  bfr _b_903(.a(_w_1135),.q(_w_1136));
  bfr _b_901(.a(_w_1133),.q(_w_1134));
  bfr _b_898(.a(_w_1130),.q(_w_1131));
  bfr _b_897(.a(_w_1129),.q(_w_1130));
  bfr _b_895(.a(_w_1127),.q(_w_1128));
  bfr _b_894(.a(_w_1126),.q(_w_1127));
  bfr _b_1003(.a(_w_1235),.q(_w_1236));
  bfr _b_925(.a(_w_1157),.q(_w_1158));
  bfr _b_892(.a(N40),.q(_w_1125));
  bfr _b_887(.a(_w_1119),.q(_w_1120));
  bfr _b_885(.a(_w_1117),.q(_w_1118));
  bfr _b_883(.a(_w_1115),.q(_w_1116));
  bfr _b_881(.a(_w_1113),.q(_w_1114));
  bfr _b_890(.a(N4),.q(_w_1123));
  bfr _b_880(.a(_w_1112),.q(_w_1113));
  bfr _b_879(.a(_w_1111),.q(_w_1112));
  bfr _b_878(.a(_w_1110),.q(_w_1111));
  bfr _b_877(.a(_w_1109),.q(_w_1110));
  bfr _b_872(.a(N21),.q(_w_1105));
  bfr _b_869(.a(_w_1101),.q(_w_1102));
  bfr _b_866(.a(_w_1098),.q(_w_1099));
  bfr _b_865(.a(_w_1097),.q(_w_1098));
  bfr _b_860(.a(_w_1092),.q(_w_1093));
  bfr _b_859(.a(_w_1091),.q(_w_1092));
  bfr _b_858(.a(N14),.q(_w_1091));
  bfr _b_857(.a(_w_1089),.q(_w_1075));
  bfr _b_854(.a(_w_1086),.q(_w_1087));
  bfr _b_853(.a(_w_1085),.q(_w_1086));
  bfr _b_850(.a(_w_1082),.q(_w_1083));
  bfr _b_849(.a(_w_1081),.q(_w_1082));
  bfr _b_847(.a(_w_1079),.q(_w_1080));
  bfr _b_840(.a(N112),.q(_w_1073));
  bfr _b_838(.a(_w_1070),.q(_w_1071));
  bfr _b_968(.a(_w_1200),.q(_w_1187));
  bfr _b_846(.a(_w_1078),.q(_w_1079));
  bfr _b_837(.a(_w_1069),.q(_w_1070));
  bfr _b_836(.a(_w_1068),.q(_w_1069));
  bfr _b_835(.a(_w_1067),.q(_w_1068));
  bfr _b_834(.a(_w_1066),.q(_w_1067));
  bfr _b_935(.a(_w_1167),.q(_w_1168));
  bfr _b_830(.a(_w_1062),.q(_w_1063));
  bfr _b_829(.a(_w_1061),.q(_w_1062));
  bfr _b_828(.a(_w_1060),.q(_w_1061));
  bfr _b_827(.a(_w_1059),.q(_w_1060));
  bfr _b_825(.a(_w_1057),.q(_w_1058));
  bfr _b_824(.a(N105),.q(_w_1057));
  bfr _b_823(.a(_w_1055),.q(_w_1054));
  bfr _b_821(.a(_w_1053),.q(n41_1));
  bfr _b_816(.a(_w_1048),.q(_w_1049));
  bfr _b_813(.a(_w_1045),.q(n72_1));
  bfr _b_812(.a(_w_1044),.q(_w_1045));
  bfr _b_953(.a(_w_1185),.q(_w_1186));
  bfr _b_826(.a(_w_1058),.q(_w_1059));
  bfr _b_811(.a(_w_1043),.q(n121_1));
  bfr _b_809(.a(_w_1041),.q(_w_1042));
  bfr _b_807(.a(_w_1039),.q(n64));
  bfr _b_806(.a(n174_1),.q(n174_2));
  bfr _b_805(.a(_w_1037),.q(n163));
  bfr _b_952(.a(_w_1184),.q(_w_1185));
  bfr _b_802(.a(_w_1034),.q(_w_1035));
  bfr _b_801(.a(_w_1033),.q(_w_1034));
  bfr _b_977(.a(_w_1209),.q(_w_1201));
  bfr _b_947(.a(_w_1179),.q(_w_1180));
  bfr _b_799(.a(_w_1031),.q(_w_1032));
  bfr _b_798(.a(_w_1030),.q(n194));
  bfr _b_900(.a(_w_1132),.q(_w_1133));
  bfr _b_794(.a(_w_1026),.q(_w_1027));
  bfr _b_793(.a(_w_1025),.q(_w_1026));
  bfr _b_792(.a(_w_1024),.q(_w_1025));
  bfr _b_789(.a(_w_1021),.q(n195_1));
  bfr _b_787(.a(_w_1019),.q(_w_1020));
  bfr _b_778(.a(_w_1010),.q(n178_1));
  bfr _b_776(.a(_w_1008),.q(_w_1009));
  bfr _b_774(.a(_w_1006),.q(n112_1));
  bfr _b_771(.a(_w_1003),.q(_w_1004));
  bfr _b_940(.a(_w_1172),.q(_w_1173));
  bfr _b_770(.a(_w_1002),.q(_w_1003));
  bfr _b_764(.a(_w_996),.q(_w_997));
  bfr _b_763(.a(_w_995),.q(n175_1));
  bfr _b_762(.a(_w_994),.q(_w_995));
  bfr _b_761(.a(_w_993),.q(_w_994));
  bfr _b_924(.a(_w_1156),.q(_w_1157));
  bfr _b_760(.a(_w_992),.q(n151_1));
  bfr _b_759(.a(_w_991),.q(n155_5));
  bfr _b_758(.a(_w_990),.q(N370));
  bfr _b_756(.a(_w_988),.q(_w_989));
  bfr _b_755(.a(_w_987),.q(_w_988));
  bfr _b_817(.a(_w_1049),.q(n46_1));
  bfr _b_754(.a(_w_986),.q(_w_987));
  bfr _b_779(.a(_w_1011),.q(_w_1012));
  bfr _b_753(.a(N370_9),.q(_w_986));
  bfr _b_752(.a(_w_984),.q(n113));
  bfr _b_750(.a(_w_982),.q(_w_983));
  bfr _b_939(.a(_w_1171),.q(_w_1172));
  bfr _b_749(.a(_w_981),.q(n156_1));
  bfr _b_748(.a(_w_980),.q(n168_1));
  bfr _b_808(.a(n121_0),.q(_w_1041));
  bfr _b_743(.a(_w_975),.q(_w_976));
  bfr _b_741(.a(n38_2),.q(n131));
  bfr _b_991(.a(_w_1223),.q(_w_1224));
  bfr _b_740(.a(_w_972),.q(n93_3));
  bfr _b_739(.a(_w_971),.q(n171_1));
  bfr _b_735(.a(_w_967),.q(_w_968));
  bfr _b_733(.a(_w_965),.q(_w_966));
  bfr _b_731(.a(_w_963),.q(n140_1));
  bfr _b_728(.a(n180_0),.q(_w_961));
  bfr _b_725(.a(_w_957),.q(_w_958));
  bfr _b_723(.a(_w_955),.q(N86_1));
  bfr _b_831(.a(_w_1063),.q(_w_1064));
  bfr _b_722(.a(_w_954),.q(_w_955));
  bfr _b_718(.a(_w_950),.q(_w_951));
  bfr _b_717(.a(_w_949),.q(_w_950));
  bfr _b_919(.a(_w_1151),.q(_w_1152));
  bfr _b_715(.a(_w_947),.q(_w_948));
  bfr _b_714(.a(_w_946),.q(_w_947));
  bfr _b_711(.a(_w_943),.q(N431));
  bfr _b_710(.a(_w_942),.q(n201));
  bfr _b_893(.a(_w_1125),.q(_w_1126));
  bfr _b_708(.a(_w_940),.q(_w_941));
  bfr _b_705(.a(_w_937),.q(n189_1));
  bfr _b_702(.a(_w_934),.q(_w_935));
  bfr _b_784(.a(_w_1016),.q(n186_1));
  bfr _b_701(.a(_w_933),.q(_w_934));
  bfr _b_783(.a(_w_1015),.q(_w_1016));
  bfr _b_698(.a(_w_930),.q(_w_931));
  bfr _b_781(.a(_w_1013),.q(_w_1014));
  bfr _b_697(.a(_w_929),.q(_w_930));
  bfr _b_695(.a(_w_927),.q(N73_1));
  bfr _b_692(.a(_w_924),.q(_w_925));
  bfr _b_691(.a(_w_923),.q(_w_924));
  bfr _b_690(.a(_w_922),.q(_w_923));
  bfr _b_736(.a(_w_968),.q(_w_969));
  bfr _b_689(.a(_w_921),.q(_w_922));
  bfr _b_682(.a(n52_5),.q(_w_915));
  bfr _b_679(.a(_w_911),.q(_w_912));
  bfr _b_678(.a(_w_910),.q(_w_911));
  bfr _b_674(.a(_w_906),.q(_w_907));
  bfr _b_839(.a(_w_1071),.q(_w_1056));
  bfr _b_673(.a(_w_905),.q(n170_1));
  bfr _b_729(.a(_w_961),.q(n180_1));
  bfr _b_671(.a(_w_903),.q(n198));
  bfr _b_670(.a(_w_902),.q(_w_903));
  bfr _b_669(.a(_w_901),.q(_w_902));
  bfr _b_663(.a(_w_895),.q(_w_896));
  bfr _b_662(.a(_w_894),.q(_w_895));
  bfr _b_661(.a(_w_893),.q(n169));
  bfr _b_658(.a(_w_890),.q(_w_891));
  bfr _b_984(.a(_w_1216),.q(_w_1217));
  bfr _b_657(.a(_w_889),.q(_w_890));
  bfr _b_981(.a(N89),.q(_w_1213));
  bfr _b_818(.a(n45_2),.q(n139));
  bfr _b_655(.a(_w_887),.q(_w_888));
  bfr _b_654(.a(_w_886),.q(N56_1));
  bfr _b_650(.a(_w_882),.q(_w_883));
  bfr _b_649(.a(_w_881),.q(_w_882));
  bfr _b_938(.a(_w_1170),.q(_w_1171));
  bfr _b_768(.a(_w_1000),.q(n146_1));
  bfr _b_648(.a(n96_0),.q(n96_1));
  bfr _b_642(.a(_w_874),.q(n46_3));
  bfr _b_638(.a(_w_870),.q(N223));
  bfr _b_637(.a(_w_869),.q(_w_870));
  bfr _b_636(.a(_w_868),.q(_w_869));
  bfr _b_635(.a(_w_867),.q(_w_868));
  bfr _b_633(.a(_w_865),.q(_w_866));
  bfr _b_630(.a(_w_862),.q(_w_863));
  bfr _b_629(.a(_w_861),.q(_w_862));
  bfr _b_876(.a(_w_1108),.q(_w_1109));
  bfr _b_747(.a(_w_979),.q(_w_980));
  bfr _b_628(.a(_w_860),.q(_w_861));
  bfr _b_627(.a(_w_859),.q(_w_860));
  bfr _b_875(.a(N27),.q(_w_1108));
  bfr _b_632(.a(_w_864),.q(_w_865));
  bfr _b_626(.a(_w_858),.q(_w_859));
  bfr _b_625(.a(_w_857),.q(_w_858));
  bfr _b_624(.a(_w_856),.q(_w_857));
  bfr _b_623(.a(_w_855),.q(_w_856));
  bfr _b_796(.a(_w_1028),.q(_w_1029));
  bfr _b_622(.a(_w_854),.q(_w_855));
  bfr _b_620(.a(_w_852),.q(_w_853));
  bfr _b_619(.a(_w_851),.q(_w_852));
  bfr _b_618(.a(_w_850),.q(_w_851));
  bfr _b_616(.a(_w_848),.q(_w_849));
  bfr _b_965(.a(_w_1197),.q(_w_1198));
  bfr _b_614(.a(_w_846),.q(_w_847));
  bfr _b_612(.a(_w_844),.q(_w_845));
  bfr _b_639(.a(_w_871),.q(n109_1));
  bfr _b_611(.a(_w_843),.q(_w_844));
  bfr _b_773(.a(_w_1005),.q(N102_1));
  bfr _b_610(.a(_w_842),.q(n68_1));
  bfr _b_609(.a(_w_841),.q(_w_842));
  bfr _b_608(.a(_w_840),.q(n38_1));
  bfr _b_602(.a(_w_834),.q(_w_835));
  bfr _b_601(.a(_w_833),.q(n62));
  bfr _b_598(.a(_w_830),.q(n93_1));
  bfr _b_596(.a(_w_828),.q(_w_829));
  bfr _b_592(.a(_w_824),.q(n111));
  bfr _b_641(.a(_w_873),.q(n62_1));
  bfr _b_591(.a(_w_823),.q(_w_824));
  bfr _b_932(.a(_w_1164),.q(_w_1165));
  bfr _b_589(.a(_w_821),.q(_w_822));
  bfr _b_588(.a(_w_820),.q(n82_1));
  bfr _b_587(.a(_w_819),.q(_w_820));
  bfr _b_584(.a(n188_0),.q(n188_1));
  bfr _b_582(.a(_w_814),.q(_w_815));
  bfr _b_886(.a(_w_1118),.q(_w_1119));
  bfr _b_667(.a(_w_899),.q(_w_900));
  bfr _b_581(.a(_w_813),.q(_w_814));
  bfr _b_578(.a(_w_810),.q(_w_811));
  bfr _b_577(.a(_w_809),.q(_w_810));
  bfr _b_709(.a(_w_941),.q(n196));
  bfr _b_576(.a(n117_0),.q(_w_809));
  bfr _b_574(.a(_w_806),.q(n128));
  bfr _b_659(.a(_w_891),.q(_w_892));
  bfr _b_573(.a(_w_805),.q(n187));
  bfr _b_572(.a(_w_804),.q(_w_805));
  bfr _b_988(.a(_w_1220),.q(_w_1221));
  bfr _b_570(.a(_w_802),.q(_w_803));
  bfr _b_569(.a(_w_801),.q(_w_802));
  bfr _b_568(.a(_w_800),.q(N73_3));
  bfr _b_590(.a(_w_822),.q(N82_1));
  bfr _b_567(.a(_w_799),.q(n51_1));
  bfr _b_868(.a(_w_1100),.q(_w_1101));
  bfr _b_621(.a(_w_853),.q(_w_854));
  bfr _b_599(.a(_w_831),.q(_w_832));
  bfr _b_566(.a(_w_798),.q(_w_799));
  bfr _b_564(.a(n51_0),.q(_w_797));
  bfr _b_563(.a(_w_795),.q(N79_1));
  bfr _b_896(.a(_w_1128),.q(_w_1129));
  bfr _b_766(.a(_w_998),.q(_w_999));
  bfr _b_685(.a(_w_917),.q(_w_918));
  bfr _b_561(.a(N79_0),.q(_w_794));
  bfr _b_560(.a(_w_792),.q(N34_5));
  bfr _b_559(.a(_w_791),.q(_w_792));
  bfr _b_557(.a(_w_789),.q(n132));
  bfr _b_556(.a(_w_788),.q(_w_789));
  bfr _b_555(.a(_w_787),.q(_w_788));
  bfr _b_917(.a(_w_1149),.q(_w_1150));
  bfr _b_549(.a(_w_781),.q(_w_782));
  bfr _b_833(.a(_w_1065),.q(_w_1066));
  bfr _b_548(.a(N76_0),.q(_w_781));
  bfr _b_786(.a(_w_1018),.q(_w_1019));
  bfr _b_665(.a(_w_897),.q(_w_898));
  bfr _b_544(.a(_w_776),.q(_w_777));
  bfr _b_543(.a(N53_0),.q(_w_776));
  bfr _b_541(.a(_w_773),.q(_w_774));
  spl2 g41_s_0(.a(n41),.q0(n41_0),.q1(_w_1051));
  spl2 g42_s_0(.a(n42),.q0(n42_0),.q1(n42_1));
  spl2 g44_s_0(.a(n44),.q0(n44_0),.q1(n44_1));
  bfr _b_486(.a(N329_9),.q(_w_719));
  bfr _b_742(.a(n167_0),.q(n183));
  maj_bbi g87(.a(n41_3),.b(n86),.c(n49_2),.q(n87));
  spl2 g46_s_0(.a(n46),.q0(n46_0),.q1(_w_1047));
  bfr _b_863(.a(_w_1095),.q(_w_1096));
  bfr _b_463(.a(_w_695),.q(_w_696));
  spl4L g55_s_1(.a(n55_0),.q0(n59),.q1(n55_5),.q2(n55_6),.q3(n55_7));
  spl4L g55_s_0(.a(n55),.q0(n55_0),.q1(n55_1),.q2(n55_2),.q3(n55_3));
  bfr _b_571(.a(_w_803),.q(_w_804));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(_w_1046));
  spl2 g72_s_0(.a(n72),.q0(n72_0),.q1(_w_1044));
  bfr _b_652(.a(_w_884),.q(_w_885));
  or_bb g89(.a(n83),.b(n88),.q(n89));
  bfr _b_458(.a(N66_0),.q(_w_691));
  spl2 g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1));
  spl2 g87_s_2(.a(n87_3),.q0(n87_5),.q1(_w_1030));
  and_bb g91(.a(N69_3),.b(n90),.q(n91));
  spl2 g87_s_0(.a(n87),.q0(n87_0),.q1(_w_1024));
  bfr _b_790(.a(_w_1022),.q(n108_5));
  bfr _b_553(.a(_w_785),.q(_w_786));
  or_bb g116(.a(n115),.b(n51_2),.q(n51_3));
  spl3L g89_s_0(.a(n89),.q0(n89_0),.q1(n89_1),.q2(n89_2));
  bfr _b_575(.a(_w_807),.q(n41_3));
  spl2 g100_s_0(.a(n100),.q0(n100_0),.q1(_w_1023));
  spl2 g108_s_2(.a(n108_2),.q0(n108_4),.q1(_w_1022));
  spl2 g108_s_1(.a(n108_1),.q0(n108_2),.q1(n108_3));
  bfr _b_797(.a(_w_1029),.q(n87_1));
  bfr _b_580(.a(_w_812),.q(_w_813));
  spl2 g121_s_0(.a(n121),.q0(n121_0),.q1(_w_1040));
  maj_bbi g158(.a(n156_1),.b(n157),.c(N86_3),.q(n158));
  bfr _b_438(.a(_w_670),.q(_w_671));
  spl3L g49_s_1(.a(n49_1),.q0(n49_4),.q1(n49_5),.q2(n49_6));
  bfr _b_800(.a(_w_1032),.q(_w_1033));
  bfr _b_499(.a(_w_731),.q(N329));
  bfr _b_510(.a(_w_742),.q(n40_1));
  bfr _b_732(.a(n73_0),.q(n73_1));
  spl2 g108_s_0(.a(n108),.q0(n108_0),.q1(n108_1));
  and_bb g85(.a(N95_3),.b(n84),.q(n85));
  spl2 g186_s_0(.a(n186),.q0(n186_0),.q1(_w_1011));
  spl2 N102_s_0(.a(N102),.q0(N102_0),.q1(_w_1001));
  spl2 g47_s_0(.a(n47),.q0(n47_0),.q1(n47_1));
  bfr _b_676(.a(_w_908),.q(_w_909));
  bfr _b_342(.a(_w_574),.q(_w_575));
  spl2 g126_s_0(.a(n126),.q0(n127),.q1(n126_1));
  bfr _b_867(.a(_w_1099),.q(_w_1100));
  or_bb g92(.a(n46_2),.b(n91),.q(n92));
  spl2 g45_s_0(.a(n45),.q0(n45_0),.q1(_w_996));
  bfr _b_429(.a(_w_661),.q(_w_662));
  spl2 g175_s_0(.a(n175),.q0(n175_0),.q1(_w_993));
  spl2 N4_s_2(.a(N4_2),.q0(N4_4),.q1(N4_5));
  bfr _b_352(.a(_w_584),.q(_w_585));
  spl4L g161_s_2(.a(N370_5),.q0(N370_9),.q1(N370_10),.q2(N370_11),.q3(_w_985));
  spl4L g106_s_0(.a(N329_0),.q0(N329_1),.q1(N329_2),.q2(N329_3),.q3(N329_4));
  bfr _b_526(.a(_w_758),.q(n56_1));
  spl2 g155_s_1(.a(n155_1),.q0(n155_2),.q1(n155_3));
  spl2 N99_s_1(.a(N99_1),.q0(N99_2),.q1(_w_982));
  bfr _b_683(.a(_w_915),.q(_w_916));
  spl3L g174_s_0(.a(n174),.q0(n174_0),.q1(n174_1),.q2(_w_1038));
  spl2 g156_s_0(.a(n156),.q0(n156_0),.q1(_w_981));
  spl2 g146_s_0(.a(n146),.q0(n146_0),.q1(_w_1000));
  spl2 g168_s_0(.a(n168),.q0(n168_0),.q1(_w_975));
  spl2 g167_s_0(.a(n167),.q0(n167_0),.q1(_w_974));
  spl2 g38_s_1(.a(n38_1),.q0(n38_2),.q1(n58_8));
  spl2 g164_s_0(.a(n164),.q0(n164_0),.q1(n164_1));
  bfr _b_910(.a(_w_1142),.q(_w_1124));
  bfr _b_603(.a(_w_835),.q(N4_1));
  spl2 g93_s_1(.a(n93_1),.q0(n93_2),.q1(_w_972));
  bfr _b_848(.a(_w_1080),.q(_w_1081));
  spl2 g171_s_0(.a(n171),.q0(n171_0),.q1(_w_965));
  and_bi g189(.a(n93_3),.b(n126_1),.q(n189));
  spl2 g180_s_1(.a(n180_1),.q0(n180_2),.q1(_w_962));
  bfr _b_470(.a(_w_702),.q(n157));
  spl2 g181_s_1(.a(n181_0),.q0(n181_2),.q1(_w_959));
  spl2 g181_s_0(.a(n181),.q0(n181_0),.q1(n181_1));
  and_bi g204(.a(n174_2),.b(_w_959),.q(n204));
  spl2 N86_s_0(.a(_w_1210),.q0(N86_0),.q1(_w_945));
  bfr _b_706(.a(_w_938),.q(_w_939));
  maj_bbi g211(.a(n180_3),.b(n209),.c(n210),.q(_w_944));
  or_bb g159(.a(n153),.b(n158),.q(n159));
  bfr _b_437(.a(_w_669),.q(_w_670));
  maj_bbi g71(.a(n69_1),.b(n70),.c(n55_5),.q(n71));
  bfr _b_443(.a(_w_675),.q(_w_676));
  bfr _b_466(.a(_w_698),.q(N82_3));
  bfr _b_382(.a(N21_0),.q(_w_615));
  bfr _b_407(.a(_w_639),.q(_w_640));
  or_bb g192(.a(n188_1),.b(n191_1),.q(n192));
  spl2 g155_s_0(.a(n155),.q0(n155_0),.q1(n155_1));
  bfr _b_819(.a(n41_0),.q(_w_1052));
  bfr _b_363(.a(_w_595),.q(_w_596));
  and_bi g185(.a(n155_4),.b(n184),.q(n185));
  bfr _b_653(.a(_w_885),.q(n166));
  spl4L g52_s_0(.a(n52),.q0(n52_0),.q1(n52_1),.q2(n52_2),.q3(n52_3));
  bfr _b_452(.a(_w_684),.q(_w_685));
  spl3L g87_s_1(.a(n87_1),.q0(n87_2),.q1(n87_3),.q2(n87_4));
  and_bb g199(.a(N115_1),.b(_w_985),.q(n199));
  spl2 N73_s_0(.a(_w_1178),.q0(N73_0),.q1(_w_926));
  and_bi g194(.a(n87_5),.b(n193),.q(n87_6));
  bfr _b_640(.a(_w_872),.q(n117_3));
  and_bi g179(.a(n178_0),.b(N27_1),.q(_w_917));
  bfr _b_841(.a(_w_1073),.q(_w_1074));
  bfr _b_521(.a(_w_753),.q(_w_754));
  and_bi g177(.a(n108_4),.b(n176),.q(n177));
  bfr _b_546(.a(_w_778),.q(_w_779));
  bfr _b_456(.a(_w_688),.q(_w_689));
  spl2 g195_s_0(.a(n195),.q0(n195_0),.q1(_w_1017));
  maj_bbi g173(.a(n171_1),.b(n172),.c(N370_6),.q(n173));
  bfr _b_403(.a(_w_635),.q(N69_1));
  bfr _b_441(.a(_w_673),.q(_w_674));
  spl2 g99_s_0(.a(n99),.q0(n99_0),.q1(_w_906));
  spl2 g170_s_0(.a(n170),.q0(n170_0),.q1(_w_904));
  and_bi g168(.a(n140_1),.b(n138_1),.q(n168));
  spl2 g73_s_0(.a(n73),.q0(n73_0),.q1(_w_964));
  maj_bbi g102(.a(n100_1),.b(n101),.c(n55_3),.q(n102));
  bfr _b_645(.a(_w_877),.q(_w_878));
  bfr _b_386(.a(_w_618),.q(_w_619));
  bfr _b_908(.a(_w_1140),.q(_w_1141));
  or_bb g58(.a(n42_0),.b(n44_1),.q(n58));
  bfr _b_675(.a(_w_907),.q(n99_1));
  bfr _b_634(.a(_w_866),.q(_w_867));
  bfr _b_489(.a(_w_721),.q(_w_722));
  spl2 g45_s_1(.a(n45_1),.q0(n45_2),.q1(_w_1050));
  maj_bbi g167(.a(n164_3),.b(n166),.c(N370_10),.q(_w_887));
  spl2 N56_s_0(.a(N56),.q0(N56_0),.q1(_w_886));
  bfr _b_959(.a(_w_1191),.q(_w_1192));
  and_bi g166(.a(n164_2),.b(n165),.q(_w_881));
  bfr _b_487(.a(_w_719),.q(_w_720));
  or_bb g209(.a(n206),.b(n208),.q(n209));
  bfr _b_861(.a(_w_1093),.q(_w_1094));
  or_bb g174(.a(n170_0),.b(n173),.q(n174));
  and_bi g163(.a(n82_6),.b(n162),.q(n82_7));
  or_bb g122(.a(n114),.b(_w_1040),.q(n122));
  bfr _b_891(.a(_w_1123),.q(_w_1122));
  and_bi g37(.a(N17_0),.b(_w_578),.q(n37));
  bfr _b_922(.a(_w_1154),.q(_w_1155));
  and_bi g38(.a(N56_0),.b(_w_668),.q(n38));
  spl2 g96_s_0(.a(n96),.q0(n96_0),.q1(_w_880));
  bfr _b_694(.a(N73_0),.q(_w_927));
  spl2 g180_s_0(.a(n180),.q0(n180_0),.q1(_w_960));
  bfr _b_376(.a(_w_608),.q(_w_609));
  bfr _b_473(.a(_w_705),.q(_w_706));
  maj_bbi g60(.a(n57_1),.b(n59),.c(n55_4),.q(n60));
  bfr _b_719(.a(_w_951),.q(_w_952));
  bfr _b_476(.a(_w_708),.q(N95_3));
  and_bi g171(.a(n132_1),.b(n130_1),.q(n171));
  bfr _b_527(.a(N14_0),.q(_w_760));
  bfr _b_769(.a(N102_0),.q(_w_1002));
  and_bi g207(.a(n197_0),.b(_w_816),.q(n207));
  and_bi g44(.a(N4_0),.b(_w_768),.q(n44));
  bfr _b_646(.a(_w_878),.q(_w_879));
  or_bb g104(.a(n103_0),.b(n94),.q(n104));
  bfr _b_874(.a(_w_1106),.q(_w_1104));
  bfr _b_814(.a(n69_0),.q(n69_1));
  bfr _b_413(.a(_w_645),.q(_w_646));
  bfr _b_734(.a(_w_966),.q(_w_967));
  bfr _b_344(.a(_w_576),.q(_w_577));
  or_bb g47(.a(n45_0),.b(_w_1047),.q(n47));
  bfr _b_391(.a(_w_623),.q(_w_624));
  maj_bbi g64(.a(n62_0),.b(n63_0),.c(N34_3),.q(_w_1039));
  spl2 g46_s_1(.a(n46_1),.q0(n46_2),.q1(_w_874));
  bfr _b_795(.a(_w_1027),.q(_w_1028));
  bfr _b_680(.a(_w_912),.q(_w_913));
  maj_bbi g195(.a(n194),.b(n87_6),.c(_w_718),.q(n195));
  bfr _b_999(.a(_w_1231),.q(_w_1232));
  or_bb g49(.a(n43),.b(n48),.q(n49));
  spl2 g117_s_1(.a(n117_1),.q0(n117_2),.q1(_w_872));
  and_bi g50(.a(N108_0),.b(_w_1001),.q(n50));
  and_bi g65(.a(n62_1),.b(_w_790),.q(n65));
  bfr _b_744(.a(_w_976),.q(_w_977));
  bfr _b_703(.a(_w_935),.q(_w_936));
  spl2 g109_s_0(.a(n109),.q0(n109_0),.q1(_w_871));
  and_bi g51(.a(N30_0),.b(_w_626),.q(n51));
  and_bb g165(.a(N14_1),.b(n164_1),.q(n165));
  bfr _b_928(.a(N60),.q(_w_1161));
  maj_bbi g205(.a(n181_3),.b(n192_1),.c(n204),.q(_w_943));
  and_bi g68(.a(N108_2),.b(_w_583),.q(n68));
  and_bb g80(.a(N1_3),.b(_w_914),.q(n80));
  and_bb g162(.a(N8_2),.b(n82_5),.q(n162));
  bfr _b_558(.a(N34_4),.q(_w_791));
  spl2 g89_s_1(.a(n89_0),.q0(n89_3),.q1(n89_4));
  bfr _b_449(.a(_w_681),.q(_w_682));
  and_bb g129(.a(N60_2),.b(_w_732),.q(n129));
  or_bb g53(.a(n49_4),.b(n52_6),.q(_w_848));
  bfr _b_979(.a(_w_1211),.q(_w_1212));
  bfr _b_686(.a(_w_918),.q(_w_919));
  bfr _b_664(.a(_w_896),.q(_w_897));
  bfr _b_349(.a(_w_581),.q(_w_582));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  maj_bbi g108(.a(n107),.b(n37_3),.c(n55_7),.q(_w_843));
  or_bb g55(.a(n52_4),.b(n54),.q(n55));
  and_bi g141(.a(n140_0),.b(_w_775),.q(n138_0));
  spl2 g57_s_0(.a(n57),.q0(n57_0),.q1(n58_4));
  and_bi g56(.a(N17_2),.b(_w_614),.q(n56));
  bfr _b_472(.a(_w_704),.q(_w_705));
  and_bi g72(.a(N82_2),.b(_w_945),.q(n72));
  bfr _b_788(.a(_w_1020),.q(_w_1021));
  bfr _b_431(.a(_w_663),.q(_w_664));
  or_bb g208(.a(n170_1),.b(n207),.q(n208));
  and_bi g99(.a(N56_2),.b(_w_680),.q(n99));
  bfr _b_496(.a(_w_728),.q(_w_729));
  bfr _b_684(.a(_w_916),.q(n52_6));
  and_bi g57(.a(n56_0),.b(N11_1),.q(n57));
  bfr _b_843(.a(N115),.q(_w_1076));
  spl2 g68_s_0(.a(n68),.q0(n68_0),.q1(_w_841));
  spl2 g82_s_2(.a(n82_3),.q0(n82_4),.q1(n82_5));
  bfr _b_506(.a(n40_2),.q(n154));
  spl2 g38_s_0(.a(n38),.q0(n38_0),.q1(_w_837));
  bfr _b_562(.a(_w_794),.q(_w_795));
  maj_bbi g93(.a(n46_3),.b(n92),.c(n49_3),.q(n93));
  bfr _b_508(.a(_w_740),.q(_w_741));
  maj_bbi g59(.a(n56_1),.b(_w_928),.c(n58_4),.q(n55_4));
  bfr _b_820(.a(_w_1052),.q(_w_1053));
  bfr _b_713(.a(N86_0),.q(_w_946));
  maj_bbi g197(.a(n195_1),.b(n196),.c(N370_8),.q(n197));
  bfr _b_791(.a(_w_1023),.q(n100_1));
  bfr _b_406(.a(_w_638),.q(_w_639));
  spl2 g132_s_0(.a(n132),.q0(n132_0),.q1(_w_836));
  bfr _b_986(.a(_w_1218),.q(_w_1219));
  spl2 N4_s_0(.a(_w_1122),.q0(N4_0),.q1(_w_834));
  or_bb g67(.a(n60),.b(n66),.q(n67));
  maj_bbi g120(.a(n117_3),.b(n119),.c(N329_2),.q(n120));
  and_bi g62(.a(n61),.b(N24_1),.q(_w_831));
  bfr _b_615(.a(_w_847),.q(n108));
  spl2 g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1));
  spl2 g82_s_1(.a(n82_1),.q0(n82_2),.q1(n82_3));
  bfr _b_726(.a(_w_958),.q(N17_1));
  maj_bbi g186(.a(n155_5),.b(n185),.c(N329_8),.q(n186));
  maj_bbi g178(.a(n108_5),.b(n177),.c(N329_11),.q(n178));
  spl2 g93_s_0(.a(n93),.q0(n93_0),.q1(_w_827));
  and_bi g69(.a(n68_0),.b(N102_1),.q(n69));
  bfr _b_547(.a(_w_779),.q(n123));
  and_bi g198(.a(n146_1),.b(n144_1),.q(_w_894));
  maj_bbi g175(.a(n120_1),.b(n121_1),.c(N370_3),.q(n175));
  maj_bbi g70(.a(n68_1),.b(_w_1046),.c(n58_5),.q(n70));
  bfr _b_660(.a(_w_892),.q(_w_893));
  or_bb g202(.a(n192_0),.b(n201),.q(n167_1));
  bfr _b_350(.a(_w_582),.q(N11_1));
  bfr _b_492(.a(_w_724),.q(_w_725));
  bfr _b_533(.a(_w_765),.q(_w_766));
  spl2 g164_s_1(.a(n164_0),.q0(n164_2),.q1(_w_1031));
  spl3L g52_s_1(.a(n52_0),.q0(n52_4),.q1(n52_5),.q2(_w_914));
  maj_bbi g66(.a(n64),.b(n65),.c(n49_5),.q(n66));
  maj_bbi g74(.a(n72_1),.b(_w_964),.c(n58_6),.q(n74));
  or_bb g42(.a(n40_0),.b(_w_1051),.q(n42));
  spl2 g182_s_0(.a(N430_0),.q0(N430_1),.q1(_w_825));
  bfr _b_851(.a(_w_1083),.q(_w_1084));
  spl2 N1_s_1(.a(N1_1),.q0(N1_2),.q1(N1_3));
  maj_bbi g75(.a(n73_1),.b(n74),.c(n55_6),.q(n75));
  bfr _b_810(.a(_w_1042),.q(_w_1043));
  spl2 g130_s_0(.a(n130),.q0(n133),.q1(n130_1));
  bfr _b_430(.a(_w_662),.q(_w_663));
  and_bi g81(.a(N4_5),.b(n80),.q(n49_0));
  bfr _b_943(.a(_w_1175),.q(_w_1176));
  spl4L g58_s_0(.a(n58),.q0(n58_0),.q1(n58_1),.q2(n58_2),.q3(n58_3));
  maj_bbi g82(.a(n79),.b(n81),.c(n49_0),.q(n82));
  and_bb g184(.a(N86_2),.b(n155_3),.q(n184));
  bfr _b_643(.a(_w_875),.q(_w_876));
  bfr _b_341(.a(_w_573),.q(_w_574));
  and_bi g83(.a(n82_0),.b(_w_607),.q(n83));
  or_bb g86(.a(n41_2),.b(n85),.q(n86));
  and_bi g134(.a(n133),.b(n130_0),.q(n134));
  and_bi g94(.a(n93_0),.b(_w_926),.q(n94));
  bfr _b_777(.a(_w_1009),.q(_w_1010));
  and_bi g73(.a(n72_0),.b(N76_1),.q(n73));
  and_bi g96(.a(n95_0),.b(N37_1),.q(n96));
  bfr _b_425(.a(_w_657),.q(N47_3));
  maj_bbi g180(.a(n178_1),.b(n179),.c(N370_4),.q(n180));
  maj_bbi g101(.a(n100_0),.b(n99_1),.c(n58_3),.q(n101));
  bfr _b_772(.a(_w_1004),.q(_w_1005));
  and_bi g157(.a(n156_0),.b(N329_4),.q(N86_3));
  bfr _b_356(.a(_w_588),.q(_w_589));
  or_bb g201(.a(n197_1),.b(n200),.q(_w_942));
  and_bi g113(.a(n112_0),.b(N329_10),.q(N99_3));
  and_bi g79(.a(N4_4),.b(n78),.q(n81));
  maj_bbi g164(.a(n163),.b(n82_7),.c(N329_7),.q(n164));
  bfr _b_359(.a(_w_591),.q(N112_1));
  and_bi g63(.a(N30_3),.b(n52_1),.q(n63));
  or_bb g150(.a(n135),.b(n149),.q(n150));
  or_bb g106(.a(n105_0),.b(n77_4),.q(N329_0));
  and_bi g109(.a(n108_0),.b(_w_636),.q(n109));
  bfr _b_605(.a(n38_0),.q(_w_838));
  and_bi g110(.a(n109_0),.b(N329_6),.q(N21_3));
  bfr _b_550(.a(_w_782),.q(_w_783));
  bfr _b_375(.a(N8_0),.q(_w_608));
  bfr _b_529(.a(_w_761),.q(_w_762));
  bfr _b_451(.a(_w_683),.q(_w_684));
  maj_bbi g111(.a(n109_1),.b(n110),.c(N21_3),.q(_w_823));
  spl4L g49_s_0(.a(n49),.q0(n79),.q1(n49_1),.q2(n49_2),.q3(n49_3));
  bfr _b_882(.a(_w_1114),.q(_w_1115));
  bfr _b_597(.a(_w_829),.q(_w_830));
  bfr _b_435(.a(_w_667),.q(N47_1));
  bfr _b_842(.a(_w_1074),.q(_w_1072));
  and_bi g112(.a(n87_2),.b(_w_568),.q(n112));
  spl2 N82_s_0(.a(N82),.q0(N82_0),.q1(_w_821));
  bfr _b_368(.a(_w_600),.q(_w_601));
  bfr _b_600(.a(_w_832),.q(_w_833));
  spl2 g82_s_0(.a(n82),.q0(n82_0),.q1(_w_817));
  or_bb g54(.a(n39_1),.b(n47_1),.q(n54));
  bfr _b_994(.a(_w_1226),.q(_w_1227));
  bfr _b_408(.a(_w_640),.q(N27_1));
  bfr _b_585(.a(_w_817),.q(_w_818));
  and_bb g118(.a(N34_5),.b(_w_808),.q(_w_812));
  and_bi g183(.a(N430_1),.b(_w_974),.q(n202));
  bfr _b_844(.a(_w_1076),.q(_w_1077));
  and_bi g119(.a(n117_2),.b(n118),.q(n119));
  and_bi g121(.a(n120_0),.b(_w_1124),.q(n121));
  or_bb g123(.a(n111),.b(n122),.q(n160));
  bfr _b_696(.a(n57_0),.q(n57_1));
  bfr _b_554(.a(_w_786),.q(_w_787));
  or_bb g125(.a(n103_1),.b(n77_1),.q(n125));
  bfr _b_822(.a(N1),.q(_w_1055));
  bfr _b_651(.a(_w_883),.q(_w_884));
  bfr _b_583(.a(_w_815),.q(n118));
  bfr _b_427(.a(_w_659),.q(_w_660));
  bfr _b_864(.a(_w_1096),.q(_w_1097));
  bfr _b_475(.a(_w_707),.q(N92_1));
  bfr _b_971(.a(_w_1203),.q(_w_1204));
  bfr _b_688(.a(_w_920),.q(_w_921));
  or_bb g48(.a(n44_0),.b(n47_0),.q(n48));
  spl2 g117_s_0(.a(n117),.q0(n117_0),.q1(_w_808));
  bfr _b_681(.a(_w_913),.q(n172));
  bfr _b_502(.a(_w_734),.q(_w_735));
  and_bb g78(.a(N1_2),.b(N4_3),.q(n78));
  maj_bbb g126(.a(N73_3),.b(n124),.c(n125),.q(n126));
  bfr _b_926(.a(_w_1158),.q(_w_1159));
  and_bb g193(.a(N99_2),.b(n87_4),.q(n193));
  and_bi g128(.a(n127),.b(n126_0),.q(_w_806));
  and_bi g187(.a(n186_0),.b(N92_1),.q(_w_801));
  spl2 N73_s_1(.a(N73_1),.q0(N73_2),.q1(_w_800));
  spl2 g41_s_1(.a(n41_1),.q0(n41_2),.q1(_w_807));
  spl2 N4_s_1(.a(N4_1),.q0(N4_2),.q1(N4_3));
  bfr _b_957(.a(_w_1189),.q(_w_1190));
  and_bi g61(.a(N30_1),.b(_w_644),.q(N24_1));
  bfr _b_870(.a(_w_1102),.q(_w_1103));
  bfr _b_355(.a(_w_587),.q(_w_588));
  bfr _b_540(.a(_w_772),.q(_w_773));
  bfr _b_967(.a(_w_1199),.q(_w_1200));
  bfr _b_631(.a(_w_863),.q(_w_864));
  maj_bbb g130(.a(N60_3),.b(n105_1),.c(n129),.q(n130));
  bfr _b_737(.a(_w_969),.q(_w_970));
  spl2 g51_s_0(.a(n51),.q0(n51_0),.q1(_w_796));
  bfr _b_927(.a(_w_1159),.q(_w_1145));
  bfr _b_757(.a(_w_989),.q(_w_990));
  spl2 N79_s_0(.a(_w_1187),.q0(N79_0),.q1(_w_793));
  and_bi g152(.a(n151_0),.b(N329_3),.q(N8_3));
  spl2 N34_s_2(.a(N34_2),.q0(N34_4),.q1(_w_790));
  bfr _b_595(.a(_w_827),.q(_w_828));
  bfr _b_593(.a(_w_825),.q(_w_826));
  maj_bbi g98(.a(n96_1),.b(n97),.c(n55_2),.q(n98));
  bfr _b_405(.a(_w_637),.q(_w_638));
  and_bb g176(.a(N21_2),.b(n108_3),.q(n176));
  spl4L g55_s_2(.a(n55_1),.q0(n38_3),.q1(n55_9),.q2(n55_10),.q3(n55_11));
  or_bb g103(.a(n102),.b(n98),.q(n103));
  bfr _b_716(.a(_w_948),.q(_w_949));
  spl2 N76_s_0(.a(N76),.q0(N76_0),.q1(_w_780));
  bfr _b_491(.a(_w_723),.q(_w_724));
  or_bb g160(.a(n150),.b(n159),.q(_w_778));
  bfr _b_416(.a(_w_648),.q(_w_649));
  and_bi g95(.a(N43_2),.b(_w_658),.q(n95));
  bfr _b_384(.a(_w_616),.q(_w_617));
  bfr _b_370(.a(_w_602),.q(N115_1));
  and_bi g90(.a(N69_2),.b(n52_3),.q(n90));
  and_bi g133(.a(n132_0),.b(_w_690),.q(n130_0));
  and_bi g200(.a(n198),.b(n199),.q(n200));
  bfr _b_1000(.a(_w_1232),.q(_w_1233));
  spl2 g138_s_0(.a(n138),.q0(n141),.q1(n138_1));
  and_bi g172(.a(n171_0),.b(N66_1),.q(_w_908));
  spl2 N53_s_0(.a(_w_1145),.q0(N53_0),.q1(_w_775));
  maj_bbi g154(.a(N82_3),.b(_w_738),.c(n58_11),.q(n40_3));
  or_bb g137(.a(n104_1),.b(n77_2),.q(n137));
  spl2 g151_s_0(.a(n151),.q0(n151_0),.q1(_w_992));
  and_bi g88(.a(n87_0),.b(_w_712),.q(n88));
  spl2 g104_s_0(.a(n104),.q0(n104_0),.q1(n104_1));
  maj_bbi g140(.a(n139),.b(n45_3),.c(n55_9),.q(_w_770));
  bfr _b_474(.a(_w_706),.q(_w_707));
  bfr _b_693(.a(_w_925),.q(n120_1));
  and_bi g142(.a(n141),.b(n138_0),.q(n142));
  and_bb g136(.a(N47_2),.b(n89_3),.q(n136));
  and_bi g151(.a(n82_2),.b(_w_759),.q(n151));
  bfr _b_498(.a(_w_730),.q(_w_731));
  spl4L g58_s_2(.a(n58_1),.q0(_w_973),.q1(n58_9),.q2(n58_10),.q3(n58_11));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(_w_1006));
  or_bb g39(.a(n37_0),.b(_w_837),.q(n39));
  maj_bbi g139(.a(N43_3),.b(_w_1050),.c(n58_9),.q(n45_3));
  bfr _b_369(.a(_w_601),.q(_w_602));
  and_bi g147(.a(n146_0),.b(_w_592),.q(n144_0));
  bfr _b_420(.a(_w_652),.q(_w_653));
  bfr _b_411(.a(_w_643),.q(N112_3));
  maj_bbi g117(.a(n116),.b(n51_3),.c(n49_6),.q(n117));
  and_bi g148(.a(n147),.b(n144_0),.q(n148));
  bfr _b_343(.a(_w_575),.q(N108_3));
  and_bi g210(.a(n175_1),.b(_w_962),.q(n210));
  bfr _b_503(.a(_w_735),.q(_w_736));
  and_bb g115(.a(N30_4),.b(n63_1),.q(n51_2));
  maj_bbi g153(.a(n151_1),.b(n152),.c(N8_3),.q(n153));
  spl2 N1_s_0(.a(_w_1054),.q0(N1_0),.q1(_w_768));
  maj_bbi g155(.a(n154),.b(n40_3),.c(n55_11),.q(_w_764));
  spl2 g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1));
  maj_bbi g203(.a(n183),.b(n202),.c(n167_1),.q(N421));
  or_bb g105(.a(n104_0),.b(n89_1),.q(n105));
  maj_bbi g170(.a(n168_1),.b(n169),.c(N370_2),.q(n170));
  spl2 N14_s_0(.a(_w_1090),.q0(N14_0),.q1(_w_759));
  bfr _b_721(.a(_w_953),.q(_w_954));
  spl2 g56_s_0(.a(n56),.q0(n56_0),.q1(_w_757));
  bfr _b_954(.a(_w_1186),.q(_w_1178));
  and_bb g143(.a(N112_2),.b(n89_4),.q(n143));
  spl4L g106_s_1(.a(N329_1),.q0(N329_5),.q1(N329_6),.q2(N329_7),.q3(N329_8));
  bfr _b_873(.a(_w_1105),.q(_w_1106));
  bfr _b_700(.a(_w_932),.q(_w_933));
  bfr _b_440(.a(_w_672),.q(_w_673));
  and_bi g190(.a(n189_0),.b(N79_1),.q(_w_749));
  and_bi g196(.a(n195_0),.b(N105_1),.q(_w_938));
  spl2 g51_s_1(.a(n51_1),.q0(n115),.q1(_w_748));
  bfr _b_724(.a(_w_956),.q(n197_1));
  bfr _b_354(.a(_w_586),.q(_w_587));
  spl2 g105_s_0(.a(n105),.q0(n105_0),.q1(n105_1));
  spl2 N17_s_0(.a(N17),.q0(N17_0),.q1(_w_957));
  bfr _b_374(.a(_w_606),.q(N17_3));
  bfr _b_419(.a(_w_651),.q(_w_652));
  spl2 g50_s_0(.a(n50),.q0(n50_0),.q1(_w_744));
  bfr _b_990(.a(_w_1222),.q(_w_1223));
  spl2 g50_s_1(.a(n50_1),.q0(n50_2),.q1(_w_743));
  bfr _b_738(.a(_w_970),.q(_w_971));
  bfr _b_462(.a(_w_694),.q(n103_1));
  spl2 g82_s_3(.a(n82_4),.q0(n82_6),.q1(_w_1037));
  bfr _b_442(.a(_w_674),.q(_w_675));
  spl2 g40_s_0(.a(n40),.q0(n40_0),.q1(_w_739));
  or_bb g77(.a(n67),.b(n76),.q(n77));
  spl2 g40_s_1(.a(n40_1),.q0(n40_2),.q1(_w_738));
  bfr _b_884(.a(_w_1116),.q(_w_1117));
  bfr _b_515(.a(_w_747),.q(n50_1));
  spl2 g189_s_0(.a(n189),.q0(n189_0),.q1(_w_929));
  bfr _b_436(.a(N50_0),.q(_w_669));
  bfr _b_871(.a(_w_1103),.q(_w_1090));
  spl2 g37_s_1(.a(n37_1),.q0(n37_2),.q1(_w_733));
  bfr _b_606(.a(_w_838),.q(_w_839));
  bfr _b_530(.a(_w_762),.q(_w_763));
  bfr _b_668(.a(_w_900),.q(_w_901));
  and_bi g84(.a(N95_2),.b(n52_2),.q(n84));
  spl3L g77_s_0(.a(n77),.q0(n77_0),.q1(n77_1),.q2(n77_2));
  bfr _b_699(.a(_w_931),.q(_w_932));
  spl2 g77_s_1(.a(n77_0),.q0(n77_3),.q1(_w_732));
  spl4L g161_s_0(.a(N370_0),.q0(N370_1),.q1(N370_2),.q2(N370_3),.q3(N370_4));
  spl4L g161_s_1(.a(N370_1),.q0(N370_5),.q1(N370_6),.q2(N370_7),.q3(N370_8));
  bfr _b_482(.a(_w_714),.q(_w_715));
  bfr _b_392(.a(_w_624),.q(_w_625));
  spl4L g106_s_2(.a(N329_5),.q0(N329_9),.q1(N329_10),.q2(N329_11),.q3(_w_718));
  spl2 N99_s_0(.a(_w_1228),.q0(N99_0),.q1(_w_712));
  and_bb g124(.a(N73_2),.b(n89_2),.q(n124));
  spl2 N95_s_0(.a(N95),.q0(N95_0),.q1(_w_709));
  bfr _b_607(.a(_w_839),.q(_w_840));
  spl2 N95_s_1(.a(N95_1),.q0(N95_2),.q1(_w_708));
  and_bi g127(.a(n93_2),.b(_w_793),.q(n126_0));
  spl2 N92_s_0(.a(_w_1214),.q0(N92_0),.q1(_w_703));
  spl2 N86_s_1(.a(N86_1),.q0(N86_2),.q1(_w_701));
  spl2 g95_s_0(.a(n95),.q0(n95_0),.q1(_w_699));
  bfr _b_765(.a(_w_997),.q(_w_998));
  bfr _b_730(.a(n180_2),.q(n180_3));
  and_bi g100(.a(n99_0),.b(N50_1),.q(n100));
  bfr _b_512(.a(_w_744),.q(_w_745));
  maj_bbi g131(.a(N56_3),.b(_w_973),.c(n58_8),.q(n55_8));
  bfr _b_358(.a(_w_590),.q(_w_591));
  spl2 N82_s_1(.a(N82_1),.q0(N82_2),.q1(_w_695));
  and_bi g40(.a(N82_0),.b(_w_780),.q(n40));
  spl2 g103_s_0(.a(n103),.q0(n103_0),.q1(_w_693));
  bfr _b_647(.a(_w_879),.q(n146));
  maj_bbi g146(.a(n145),.b(n50_3),.c(n55_10),.q(_w_875));
  spl2 N60_s_0(.a(_w_1160),.q0(N60_0),.q1(_w_680));
  bfr _b_545(.a(_w_777),.q(N53_1));
  spl2 g178_s_0(.a(n178),.q0(n178_0),.q1(_w_1007));
  spl2 N8_s_1(.a(N8_1),.q0(N8_2),.q1(_w_678));
  bfr _b_845(.a(_w_1077),.q(_w_1078));
  spl2 N60_s_1(.a(N60_1),.q0(N60_2),.q1(_w_677));
  bfr _b_996(.a(N99),.q(_w_1229));
  bfr _b_707(.a(_w_939),.q(_w_940));
  spl2 N56_s_1(.a(N56_1),.q0(N56_2),.q1(_w_672));
  bfr _b_565(.a(_w_797),.q(_w_798));
  bfr _b_481(.a(_w_713),.q(_w_714));
  bfr _b_644(.a(_w_876),.q(_w_877));
  spl2 N50_s_0(.a(N50),.q0(N50_0),.q1(_w_668));
  spl2 N47_s_0(.a(_w_1143),.q0(N47_0),.q1(_w_658));
  bfr _b_448(.a(N60_0),.q(_w_681));
  spl2 N47_s_1(.a(N47_1),.q0(N47_2),.q1(_w_657));
  spl2 N43_s_0(.a(N43),.q0(N43_0),.q1(_w_656));
  bfr _b_998(.a(_w_1230),.q(_w_1231));
  bfr _b_444(.a(_w_676),.q(N56_3));
  spl2 N37_s_0(.a(N37),.q0(N37_0),.q1(_w_647));
  bfr _b_804(.a(_w_1036),.q(n164_3));
  spl3L N30_s_0(.a(N30),.q0(N30_0),.q1(N34_0),.q2(_w_644));
  or_bb g161(.a(n123),.b(n160),.q(N370_0));
  spl2 N112_s_1(.a(N112_1),.q0(N112_2),.q1(_w_643));
  bfr _b_852(.a(_w_1084),.q(_w_1085));
  bfr _b_775(.a(_w_1007),.q(_w_1008));
  bfr _b_337(.a(_w_569),.q(_w_570));
  bfr _b_531(.a(_w_763),.q(N14_1));
  spl2 g120_s_0(.a(n120),.q0(n120_0),.q1(_w_920));
  spl2 N30_s_1(.a(N30_2),.q0(N30_3),.q1(_w_641));
  spl2 N27_s_0(.a(_w_1107),.q0(N27_0),.q1(_w_636));
  bfr _b_746(.a(_w_978),.q(_w_979));
  spl2 N69_s_0(.a(N69),.q0(N69_0),.q1(_w_633));
  bfr _b_379(.a(_w_611),.q(N8_1));
  bfr _b_677(.a(_w_909),.q(_w_910));
  spl2 N69_s_1(.a(N69_1),.q0(N69_2),.q1(_w_632));
  spl2 N34_s_0(.a(N34),.q0(N30_1),.q1(_w_627));
  spl2 N34_s_1(.a(N34_1),.q0(N34_2),.q1(N34_3));
  spl2 N24_s_0(.a(N24),.q0(N24_0),.q1(_w_626));
  bfr _b_594(.a(_w_826),.q(N430));
  and_bi g206(.a(n191_0),.b(_w_1038),.q(n206));
  spl2 N21_s_0(.a(_w_1104),.q0(N21_0),.q1(_w_614));
  spl2 N21_s_1(.a(N21_1),.q0(N21_2),.q1(_w_612));
  bfr _b_745(.a(_w_977),.q(_w_978));
  spl2 N8_s_0(.a(_w_1201),.q0(N8_0),.q1(_w_607));
  spl2 N17_s_1(.a(N17_1),.q0(N17_2),.q1(_w_603));
  bfr _b_727(.a(n181_2),.q(n181_3));
  spl2 N115_s_0(.a(_w_1075),.q0(N115_0),.q1(_w_592));
  bfr _b_409(.a(_w_641),.q(_w_642));
  spl2 N112_s_0(.a(_w_1072),.q0(N112_0),.q1(_w_583));
  and_bi g46(.a(N69_0),.b(_w_1162),.q(n46));
  bfr _b_377(.a(_w_609),.q(_w_610));
  bfr _b_907(.a(_w_1139),.q(_w_1140));
  spl2 g39_s_0(.a(n39),.q0(n39_0),.q1(n39_1));
  spl2 N11_s_0(.a(N11),.q0(N11_0),.q1(_w_578));
  bfr _b_524(.a(_w_756),.q(n190));
  spl2 N108_s_0(.a(N108),.q0(N108_0),.q1(_w_576));
  spl2 N108_s_1(.a(N108_1),.q0(N108_2),.q1(_w_572));
  bfr _b_720(.a(_w_952),.q(_w_953));
  spl2 N105_s_0(.a(_w_1056),.q0(N105_0),.q1(_w_568));
  bfr _b_336(.a(N105_0),.q(_w_569));
  bfr _b_338(.a(_w_570),.q(_w_571));
  bfr _b_339(.a(_w_571),.q(N105_1));
  bfr _b_507(.a(_w_739),.q(_w_740));
  bfr _b_340(.a(_w_572),.q(_w_573));
  bfr _b_367(.a(_w_599),.q(_w_600));
  bfr _b_421(.a(_w_653),.q(_w_654));
  spl2 g144_s_0(.a(n144),.q0(n147),.q1(n144_1));
  maj_bbi g145(.a(N108_3),.b(_w_743),.c(n58_10),.q(n50_3));
  bfr _b_497(.a(_w_729),.q(_w_730));
  bfr _b_345(.a(_w_577),.q(N108_1));
  bfr _b_346(.a(N11_0),.q(_w_579));
  bfr _b_347(.a(_w_579),.q(_w_580));
  bfr _b_501(.a(n37_2),.q(n107));
  bfr _b_348(.a(_w_580),.q(_w_581));
  bfr _b_902(.a(_w_1134),.q(_w_1135));
  bfr _b_351(.a(N112_0),.q(_w_584));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(_w_963));
  bfr _b_483(.a(_w_715),.q(_w_716));
  bfr _b_353(.a(_w_585),.q(_w_586));
  bfr _b_357(.a(_w_589),.q(_w_590));
  bfr _b_815(.a(n46_0),.q(_w_1048));
  bfr _b_785(.a(_w_1017),.q(_w_1018));
  bfr _b_751(.a(_w_983),.q(_w_984));
  bfr _b_509(.a(_w_741),.q(_w_742));
  bfr _b_479(.a(_w_711),.q(N95_1));
  spl4L g58_s_1(.a(n58_0),.q0(_w_928),.q1(n58_5),.q2(n58_6),.q3(n58_7));
  and_bi g41(.a(N95_0),.b(_w_1213),.q(n41));
  bfr _b_360(.a(N115_0),.q(_w_593));
  maj_bbb g144(.a(N112_3),.b(n137_0),.c(n143),.q(n144));
  bfr _b_361(.a(_w_593),.q(_w_594));
  bfr _b_362(.a(_w_594),.q(_w_595));
  bfr _b_364(.a(_w_596),.q(_w_597));
  bfr _b_500(.a(n77_3),.q(n77_4));
  bfr _b_365(.a(_w_597),.q(_w_598));
  bfr _b_371(.a(_w_603),.q(_w_604));
  bfr _b_398(.a(_w_630),.q(_w_631));
  bfr _b_982(.a(N92),.q(_w_1215));
  bfr _b_372(.a(_w_604),.q(_w_605));
  bfr _b_373(.a(_w_605),.q(_w_606));
  bfr _b_380(.a(_w_612),.q(_w_613));
  bfr _b_782(.a(_w_1014),.q(_w_1015));
  bfr _b_586(.a(_w_818),.q(_w_819));
  bfr _b_381(.a(_w_613),.q(n110));
  bfr _b_383(.a(_w_615),.q(_w_616));
  maj_bbb g138(.a(N47_3),.b(n136),.c(n137_1),.q(n138));
  bfr _b_518(.a(_w_750),.q(_w_751));
  bfr _b_704(.a(_w_936),.q(_w_937));
  bfr _b_385(.a(_w_617),.q(_w_618));
  bfr _b_832(.a(_w_1064),.q(_w_1065));
  bfr _b_666(.a(_w_898),.q(_w_899));
  or_bb g76(.a(n71),.b(n75),.q(n76));
  maj_bbi g107(.a(N17_3),.b(_w_733),.c(n58_7),.q(n37_3));
  bfr _b_387(.a(_w_619),.q(_w_620));
  bfr _b_388(.a(_w_620),.q(_w_621));
  bfr _b_389(.a(_w_621),.q(_w_622));
  bfr _b_579(.a(_w_811),.q(n117_1));
  spl2 g37_s_0(.a(n37),.q0(n37_0),.q1(_w_734));
  bfr _b_390(.a(_w_622),.q(_w_623));
  bfr _b_604(.a(_w_836),.q(n132_1));
  bfr _b_393(.a(_w_625),.q(N21_1));
  bfr _b_395(.a(_w_627),.q(_w_628));
  bfr _b_495(.a(_w_727),.q(_w_728));
  spl2 N66_s_0(.a(_w_1163),.q0(N66_0),.q1(_w_690));
  bfr _b_402(.a(_w_634),.q(_w_635));
  bfr _b_493(.a(_w_725),.q(_w_726));
  bfr _b_396(.a(_w_628),.q(_w_629));
  maj_bbi g188(.a(n186_1),.b(n187),.c(N370_7),.q(n188));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(_w_816));
  bfr _b_397(.a(_w_629),.q(_w_630));
  bfr _b_399(.a(_w_631),.q(N34_1));
  spl2 g197_s_0(.a(n197),.q0(n197_0),.q1(_w_956));
  bfr _b_516(.a(_w_748),.q(n116));
  bfr _b_400(.a(_w_632),.q(N69_3));
  bfr _b_528(.a(_w_760),.q(_w_761));
  bfr _b_401(.a(_w_633),.q(_w_634));
  bfr _b_542(.a(_w_774),.q(n140));
  bfr _b_410(.a(_w_642),.q(N30_4));
  bfr _b_412(.a(N34_0),.q(_w_645));
  bfr _b_378(.a(_w_610),.q(_w_611));
  bfr _b_505(.a(_w_737),.q(n37_1));
  bfr _b_415(.a(N37_0),.q(_w_648));
  bfr _b_417(.a(_w_649),.q(_w_650));
  bfr _b_687(.a(_w_919),.q(n179));
  bfr _b_418(.a(_w_650),.q(N37_1));
  bfr _b_422(.a(_w_654),.q(_w_655));
  bfr _b_423(.a(_w_655),.q(N43_3));
  bfr _b_888(.a(_w_1120),.q(_w_1121));
  spl2 g155_s_2(.a(n155_2),.q0(n155_4),.q1(_w_991));
  bfr _b_424(.a(_w_656),.q(N43_1));
  bfr _b_539(.a(_w_771),.q(_w_772));
  or_bb g135(.a(n128),.b(n134),.q(n135));
  bfr _b_426(.a(N47_0),.q(_w_659));
  or_bb g181(.a(n175_0),.b(_w_960),.q(n181));
  bfr _b_428(.a(_w_660),.q(_w_661));
  bfr _b_551(.a(_w_783),.q(_w_784));
  maj_bbi g114(.a(n112_1),.b(n113),.c(N99_3),.q(n114));
  bfr _b_432(.a(_w_664),.q(_w_665));
  maj_bbi g132(.a(n131),.b(n38_3),.c(n55_8),.q(_w_785));
  bfr _b_394(.a(N24_0),.q(n61));
  bfr _b_478(.a(_w_710),.q(_w_711));
  bfr _b_434(.a(_w_666),.q(_w_667));
  bfr _b_613(.a(_w_845),.q(_w_846));
  bfr _b_439(.a(_w_671),.q(N50_1));
  spl2 g62_s_0(.a(n62),.q0(n62_0),.q1(_w_873));
  and_bi g156(.a(n155_0),.b(_w_703),.q(n156));
  bfr _b_446(.a(_w_678),.q(_w_679));
  bfr _b_617(.a(_w_849),.q(_w_850));
  bfr _b_447(.a(_w_679),.q(n152));
  bfr _b_450(.a(_w_682),.q(_w_683));
  bfr _b_453(.a(_w_685),.q(_w_686));
  bfr _b_780(.a(_w_1012),.q(_w_1013));
  bfr _b_454(.a(_w_686),.q(_w_687));
  bfr _b_455(.a(_w_687),.q(_w_688));
  bfr _b_889(.a(_w_1121),.q(_w_1107));
  bfr _b_464(.a(_w_696),.q(_w_697));
  bfr _b_457(.a(_w_689),.q(N60_1));
  bfr _b_921(.a(_w_1153),.q(_w_1154));
  bfr _b_459(.a(_w_691),.q(_w_692));
  bfr _b_460(.a(_w_692),.q(N66_1));
  bfr _b_803(.a(_w_1035),.q(_w_1036));
  bfr _b_461(.a(_w_693),.q(_w_694));
  bfr _b_465(.a(_w_697),.q(_w_698));
  and_bi g45(.a(N43_0),.b(_w_647),.q(n45));
  bfr _b_467(.a(_w_699),.q(_w_700));
  bfr _b_504(.a(_w_736),.q(_w_737));
  bfr _b_468(.a(_w_700),.q(n95_1));
  bfr _b_404(.a(N27_0),.q(_w_637));
  bfr _b_469(.a(_w_701),.q(_w_702));
  bfr _b_471(.a(N92_0),.q(_w_704));
  bfr _b_856(.a(_w_1088),.q(_w_1089));
  bfr _b_477(.a(_w_709),.q(_w_710));
  bfr _b_767(.a(_w_999),.q(n45_1));
  bfr _b_445(.a(_w_677),.q(N60_3));
  or_bb g149(.a(n142),.b(n148),.q(n149));
  bfr _b_480(.a(N99_0),.q(_w_713));
  bfr _b_513(.a(_w_745),.q(_w_746));
  bfr _b_484(.a(_w_716),.q(_w_717));
  bfr _b_485(.a(_w_717),.q(N99_1));
  bfr _b_899(.a(_w_1131),.q(_w_1132));
  bfr _b_552(.a(_w_784),.q(N76_1));
  or_bb g52(.a(n50_0),.b(_w_796),.q(n52));
  bfr _b_366(.a(_w_598),.q(_w_599));
  spl2 N43_s_1(.a(N43_1),.q0(N43_2),.q1(_w_651));
  bfr _b_488(.a(_w_720),.q(_w_721));
  bfr _b_514(.a(_w_746),.q(_w_747));
  bfr _b_862(.a(_w_1094),.q(_w_1095));
  bfr _b_490(.a(_w_722),.q(_w_723));
  bfr _b_904(.a(_w_1136),.q(_w_1137));
  bfr _b_494(.a(_w_726),.q(_w_727));
  bfr _b_414(.a(_w_646),.q(N30_2));
  bfr _b_511(.a(n50_2),.q(n145));
  bfr _b_517(.a(_w_749),.q(_w_750));
  bfr _b_519(.a(_w_751),.q(_w_752));
  bfr _b_855(.a(_w_1087),.q(_w_1088));
  bfr _b_520(.a(_w_752),.q(_w_753));
  bfr _b_433(.a(_w_665),.q(_w_666));
  bfr _b_522(.a(_w_754),.q(_w_755));
  bfr _b_672(.a(_w_904),.q(_w_905));
  bfr _b_523(.a(_w_755),.q(_w_756));
  and_bi g169(.a(n168_0),.b(N53_1),.q(_w_889));
  bfr _b_525(.a(_w_757),.q(_w_758));
  bfr _b_532(.a(_w_764),.q(_w_765));
  bfr _b_712(.a(_w_944),.q(N432));
  bfr _b_534(.a(_w_766),.q(_w_767));
  maj_bbi g191(.a(n189_1),.b(n190),.c(N370_11),.q(n191));
  or_bb g182(.a(n174_0),.b(n181_1),.q(N430_0));
  or_bb g43(.a(n39_0),.b(n42_1),.q(n43));
  bfr _b_535(.a(_w_767),.q(n155));
  bfr _b_656(.a(_w_888),.q(n167));
  maj_bbi g97(.a(n95_1),.b(_w_880),.c(n58_2),.q(n97));
  bfr _b_536(.a(N1_0),.q(_w_769));
  bfr _b_537(.a(_w_769),.q(N1_1));
  bfr _b_538(.a(_w_770),.q(_w_771));
endmodule
