module c3540 ( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 , G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G6 , G7 , G8 , G9 ;
  output G3519 , G3520 , G3521 , G3522 , G3523 , G3524 , G3525 , G3526 , G3527 , G3528 , G3529 , G3530 , G3531 , G3532 , G3533 , G3534 , G3535 , G3536 , G3537 , G3538 , G3539 , G3540 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 ;
  assign n51 = G8 | G9 ;
  assign n52 = G10 | G7 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = G12 | G13 ;
  assign n55 = ~G11 | ~n54 ;
  assign n56 = G1 | G3 ;
  assign n57 = G32 & ~G9 ;
  assign n58 = G31 & ~G8 ;
  assign n59 = n57 | n58 ;
  assign n60 = ~G13 & G36 ;
  assign n61 = ~G14 & G37 ;
  assign n62 = n60 | n61 ;
  assign n63 = n59 | n62 ;
  assign n64 = ~G11 & G34 ;
  assign n65 = ~G12 & G35 ;
  assign n66 = n64 | n65 ;
  assign n67 = ~G10 & G33 ;
  assign n68 = G30 & ~G7 ;
  assign n69 = n67 | n68 ;
  assign n70 = n66 | n69 ;
  assign n71 = n63 | n70 ;
  assign n72 = n56 & n71 ;
  assign n73 = ~G1 & G2 ;
  assign n74 = ~G3 & n73 ;
  assign n75 = ~G7 & n51 ;
  assign n76 = n74 & n75 ;
  assign n77 = G2 | n56 ;
  assign n78 = G35 | G36 ;
  assign n79 = G34 & n78 ;
  assign n80 = ~n77 & n79 ;
  assign n81 = n76 | n80 ;
  assign n82 = ~n72 & ~n81 ;
  assign n83 = G36 | G37 ;
  assign n84 = G36 & G37 ;
  assign n85 = n83 & ~n84 ;
  assign n86 = G34 & ~G35 ;
  assign n87 = ~G34 & G35 ;
  assign n88 = n86 | n87 ;
  assign n89 = n85 | n88 ;
  assign n90 = n85 & n88 ;
  assign n91 = n89 & ~n90 ;
  assign n92 = G30 & ~G31 ;
  assign n93 = ~G30 & G31 ;
  assign n94 = n92 | n93 ;
  assign n95 = G32 | G33 ;
  assign n96 = G32 & G33 ;
  assign n97 = n95 & ~n96 ;
  assign n98 = n94 | n97 ;
  assign n99 = n94 & n97 ;
  assign n100 = n98 & ~n99 ;
  assign n101 = n91 | n100 ;
  assign n102 = n91 & n100 ;
  assign n103 = n101 & ~n102 ;
  assign n104 = G8 & G9 ;
  assign n105 = n51 & ~n104 ;
  assign n106 = G10 & G7 ;
  assign n107 = n52 & ~n106 ;
  assign n108 = ~n105 & n107 ;
  assign n109 = n105 & ~n107 ;
  assign n110 = n108 | n109 ;
  assign n111 = ~G11 & G13 ;
  assign n112 = G11 & ~G13 ;
  assign n113 = n111 | n112 ;
  assign n114 = G12 | G14 ;
  assign n115 = G12 & G14 ;
  assign n116 = n114 & ~n115 ;
  assign n117 = n113 & ~n116 ;
  assign n118 = ~n113 & n116 ;
  assign n119 = n117 | n118 ;
  assign n120 = n110 & n119 ;
  assign n121 = n110 | n119 ;
  assign n122 = ~n120 & n121 ;
  assign n123 = G3 & n73 ;
  assign n124 = G7 | n123 ;
  assign n125 = ~G1 & G3 ;
  assign n126 = G1 & G2 ;
  assign n127 = G1 & G3 ;
  assign n128 = G4 & n127 ;
  assign n129 = n126 | n128 ;
  assign n130 = n125 | n129 ;
  assign n131 = G7 & n130 ;
  assign n132 = n124 & ~n131 ;
  assign n133 = G7 | n51 ;
  assign n134 = G3 & n133 ;
  assign n135 = G3 | G4 ;
  assign n136 = G21 & ~n135 ;
  assign n137 = ~G3 & G4 ;
  assign n138 = ~G8 & n137 ;
  assign n139 = n136 | n138 ;
  assign n140 = n134 | n139 ;
  assign n141 = n129 & n140 ;
  assign n142 = n132 | n141 ;
  assign n143 = G25 | G26 ;
  assign n144 = G5 | G6 ;
  assign n145 = ~G1 & n144 ;
  assign n146 = G4 & G5 ;
  assign n147 = n126 & ~n146 ;
  assign n148 = G38 & ~n147 ;
  assign n149 = n145 & n148 ;
  assign n150 = G30 & ~n145 ;
  assign n151 = G4 | G49 ;
  assign n152 = G28 & ~n151 ;
  assign n153 = G10 & ~G4 ;
  assign n154 = G29 & G4 ;
  assign n155 = n153 | n154 ;
  assign n156 = n152 | n155 ;
  assign n157 = n150 | n156 ;
  assign n158 = ~n147 & n157 ;
  assign n159 = n149 | n158 ;
  assign n160 = n143 & ~n159 ;
  assign n161 = n142 | n160 ;
  assign n162 = G23 | G24 ;
  assign n163 = ~n159 & n162 ;
  assign n164 = n142 & n163 ;
  assign n165 = n161 & ~n164 ;
  assign n166 = G8 & n130 ;
  assign n167 = G8 | n123 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = G3 & n105 ;
  assign n170 = ~G9 & n137 ;
  assign n171 = G22 & ~G3 ;
  assign n172 = ~G4 & n171 ;
  assign n173 = n170 | n172 ;
  assign n174 = n169 | n173 ;
  assign n175 = n129 & n174 ;
  assign n176 = n168 | n175 ;
  assign n177 = G31 & ~n145 ;
  assign n178 = G29 & ~n151 ;
  assign n179 = G11 | G4 ;
  assign n180 = ~G30 & G4 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n178 | n181 ;
  assign n183 = n177 | n182 ;
  assign n184 = ~n147 & n183 ;
  assign n185 = n149 | n184 ;
  assign n186 = n143 & ~n185 ;
  assign n187 = n176 | n186 ;
  assign n188 = n162 & ~n185 ;
  assign n189 = n176 & n188 ;
  assign n190 = n187 & ~n189 ;
  assign n191 = n165 & n190 ;
  assign n192 = G3 & n129 ;
  assign n193 = n130 & ~n192 ;
  assign n194 = G10 & ~n193 ;
  assign n195 = ~G10 & n123 ;
  assign n196 = G8 | n135 ;
  assign n197 = ~G11 & n137 ;
  assign n198 = n196 & ~n197 ;
  assign n199 = n129 & ~n198 ;
  assign n200 = n195 | n199 ;
  assign n201 = n194 | n200 ;
  assign n202 = G33 & ~n145 ;
  assign n203 = G31 & ~n151 ;
  assign n204 = G13 | G4 ;
  assign n205 = ~G32 & G4 ;
  assign n206 = n204 & ~n205 ;
  assign n207 = n203 | n206 ;
  assign n208 = n202 | n207 ;
  assign n209 = ~n147 & n208 ;
  assign n210 = n149 | n209 ;
  assign n211 = n143 & ~n210 ;
  assign n212 = n201 | n211 ;
  assign n213 = n162 & ~n210 ;
  assign n214 = n201 & n213 ;
  assign n215 = n212 & ~n214 ;
  assign n216 = n123 | n192 ;
  assign n217 = ~G9 & n216 ;
  assign n218 = G7 & ~n135 ;
  assign n219 = G10 & n137 ;
  assign n220 = n218 | n219 ;
  assign n221 = n129 & n220 ;
  assign n222 = G9 & ~n130 ;
  assign n223 = n221 | n222 ;
  assign n224 = n217 | n223 ;
  assign n225 = G32 & ~n145 ;
  assign n226 = G30 & ~n151 ;
  assign n227 = G12 | G4 ;
  assign n228 = ~G31 & G4 ;
  assign n229 = n227 & ~n228 ;
  assign n230 = n226 | n229 ;
  assign n231 = n225 | n230 ;
  assign n232 = ~n147 & n231 ;
  assign n233 = n149 | n232 ;
  assign n234 = n143 & ~n233 ;
  assign n235 = n224 | n234 ;
  assign n236 = n162 & ~n233 ;
  assign n237 = n224 & n236 ;
  assign n238 = n235 & ~n237 ;
  assign n239 = n215 & n238 ;
  assign n240 = n191 & n239 ;
  assign n241 = G11 | n54 ;
  assign n242 = G3 & n241 ;
  assign n243 = G9 | n135 ;
  assign n244 = ~G12 & n137 ;
  assign n245 = n243 & ~n244 ;
  assign n246 = ~n242 & n245 ;
  assign n247 = n129 & ~n246 ;
  assign n248 = ~G1 & G4 ;
  assign n249 = n123 | n248 ;
  assign n250 = n129 | n249 ;
  assign n251 = G11 & ~n250 ;
  assign n252 = ~G11 & n123 ;
  assign n253 = n251 | n252 ;
  assign n254 = n247 | n253 ;
  assign n255 = G32 & ~n151 ;
  assign n256 = G14 | G4 ;
  assign n257 = ~G33 & G4 ;
  assign n258 = n256 & ~n257 ;
  assign n259 = n255 | n258 ;
  assign n260 = G1 | G6 ;
  assign n261 = G38 | n260 ;
  assign n262 = ~G34 & n260 ;
  assign n263 = n261 & ~n262 ;
  assign n264 = n259 | n263 ;
  assign n265 = ~n147 & n264 ;
  assign n266 = n162 & ~n265 ;
  assign n267 = n254 & n266 ;
  assign n268 = n143 & ~n265 ;
  assign n269 = n254 | n268 ;
  assign n270 = ~n267 & n269 ;
  assign n271 = G12 | n123 ;
  assign n272 = G12 & n250 ;
  assign n273 = n271 & ~n272 ;
  assign n274 = G12 & G13 ;
  assign n275 = n54 & ~n274 ;
  assign n276 = n192 & n275 ;
  assign n277 = ~G3 & n126 ;
  assign n278 = G13 & G4 ;
  assign n279 = n153 | n278 ;
  assign n280 = n277 & n279 ;
  assign n281 = n276 | n280 ;
  assign n282 = n273 | n281 ;
  assign n283 = G5 | n260 ;
  assign n284 = n148 & ~n283 ;
  assign n285 = G35 & n283 ;
  assign n286 = G33 & ~n151 ;
  assign n287 = G39 | G4 ;
  assign n288 = ~G34 & G4 ;
  assign n289 = n287 & ~n288 ;
  assign n290 = n286 | n289 ;
  assign n291 = n285 | n290 ;
  assign n292 = ~n147 & n291 ;
  assign n293 = n284 | n292 ;
  assign n294 = n162 & ~n293 ;
  assign n295 = n282 & n294 ;
  assign n296 = n143 & ~n293 ;
  assign n297 = n282 | n296 ;
  assign n298 = ~n295 & n297 ;
  assign n299 = n270 & n298 ;
  assign n300 = ~G13 & n216 ;
  assign n301 = G13 & ~n250 ;
  assign n302 = G14 & G4 ;
  assign n303 = n179 & ~n302 ;
  assign n304 = n277 & ~n303 ;
  assign n305 = n301 | n304 ;
  assign n306 = n300 | n305 ;
  assign n307 = G36 & n283 ;
  assign n308 = G35 & G4 ;
  assign n309 = ~G4 & G40 ;
  assign n310 = n308 | n309 ;
  assign n311 = G34 & ~n151 ;
  assign n312 = n310 | n311 ;
  assign n313 = n307 | n312 ;
  assign n314 = ~n147 & n313 ;
  assign n315 = n284 | n314 ;
  assign n316 = n162 & ~n315 ;
  assign n317 = n306 & n316 ;
  assign n318 = n143 & ~n315 ;
  assign n319 = n306 | n318 ;
  assign n320 = ~n317 & n319 ;
  assign n321 = n299 & n320 ;
  assign n322 = ~n192 & n250 ;
  assign n323 = G14 & ~n322 ;
  assign n324 = ~G14 & n123 ;
  assign n325 = G39 & G4 ;
  assign n326 = n227 & ~n325 ;
  assign n327 = n277 & ~n326 ;
  assign n328 = n324 | n327 ;
  assign n329 = n323 | n328 ;
  assign n330 = G37 & n283 ;
  assign n331 = G36 & G4 ;
  assign n332 = ~G4 & G41 ;
  assign n333 = n331 | n332 ;
  assign n334 = G35 & ~n151 ;
  assign n335 = n333 | n334 ;
  assign n336 = n330 | n335 ;
  assign n337 = ~n147 & n336 ;
  assign n338 = n284 | n337 ;
  assign n339 = n162 & ~n338 ;
  assign n340 = n329 & n339 ;
  assign n341 = n143 & ~n338 ;
  assign n342 = n329 | n341 ;
  assign n343 = ~n340 & n342 ;
  assign n344 = n321 & n343 ;
  assign n345 = n240 & n344 ;
  assign n346 = n321 & n340 ;
  assign n347 = n299 & n317 ;
  assign n348 = n269 & n295 ;
  assign n349 = n267 | n348 ;
  assign n350 = n347 | n349 ;
  assign n351 = n346 | n350 ;
  assign n352 = n240 & n351 ;
  assign n353 = n214 & n235 ;
  assign n354 = n237 | n353 ;
  assign n355 = n191 & n354 ;
  assign n356 = n161 & n189 ;
  assign n357 = n164 | n356 ;
  assign n358 = n355 | n357 ;
  assign n359 = n352 | n358 ;
  assign n360 = G27 & G48 ;
  assign n361 = ~n77 & n360 ;
  assign n362 = n306 & n361 ;
  assign n363 = n320 | n362 ;
  assign n364 = n320 & n362 ;
  assign n365 = n363 & ~n364 ;
  assign n366 = n329 & n361 ;
  assign n367 = n343 | n366 ;
  assign n368 = n343 & n366 ;
  assign n369 = n367 & ~n368 ;
  assign n370 = G47 & n369 ;
  assign n371 = ~n365 & n370 ;
  assign n372 = G5 & ~n77 ;
  assign n373 = n75 & ~n372 ;
  assign n374 = n351 & ~n361 ;
  assign n375 = ~G1 & n374 ;
  assign n376 = n373 | n375 ;
  assign n377 = ~G2 & n137 ;
  assign n378 = n369 & n377 ;
  assign n379 = ~G6 & n372 ;
  assign n380 = ~G23 & G3 ;
  assign n381 = n73 & ~n380 ;
  assign n382 = G25 & G3 ;
  assign n383 = G24 & G3 ;
  assign n384 = G26 & ~n383 ;
  assign n385 = n382 & n384 ;
  assign n386 = G39 | G43 ;
  assign n387 = ~n385 & n386 ;
  assign n388 = ~G3 & G41 ;
  assign n389 = G4 & ~n388 ;
  assign n390 = ~n387 & n389 ;
  assign n391 = G24 | n143 ;
  assign n392 = G3 & n391 ;
  assign n393 = G40 & n392 ;
  assign n394 = G26 | n383 ;
  assign n395 = n382 | n394 ;
  assign n396 = G44 & n395 ;
  assign n397 = n393 | n396 ;
  assign n398 = ~n382 & n384 ;
  assign n399 = G41 | G45 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = n382 & ~n394 ;
  assign n402 = G42 | G46 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = n400 | n403 ;
  assign n405 = n397 | n404 ;
  assign n406 = n390 & ~n405 ;
  assign n407 = G3 & n398 ;
  assign n408 = G11 | n407 ;
  assign n409 = G13 | n385 ;
  assign n410 = n408 & n409 ;
  assign n411 = G9 | n385 ;
  assign n412 = G7 | n398 ;
  assign n413 = n411 & n412 ;
  assign n414 = G10 | n401 ;
  assign n415 = ~G8 & n395 ;
  assign n416 = n414 & ~n415 ;
  assign n417 = n413 & n416 ;
  assign n418 = G22 & ~n401 ;
  assign n419 = G4 | n418 ;
  assign n420 = ~G12 & n392 ;
  assign n421 = n419 | n420 ;
  assign n422 = n417 & ~n421 ;
  assign n423 = n410 & n422 ;
  assign n424 = n406 | n423 ;
  assign n425 = ~n381 & n424 ;
  assign n426 = n379 & ~n425 ;
  assign n427 = ~n378 & n426 ;
  assign n428 = G47 & ~n369 ;
  assign n429 = ~G47 & n369 ;
  assign n430 = n379 | n429 ;
  assign n431 = n428 | n430 ;
  assign n432 = n427 | ~n431 ;
  assign n433 = n201 & n361 ;
  assign n434 = n215 | n433 ;
  assign n435 = n215 & n433 ;
  assign n436 = n434 & ~n435 ;
  assign n437 = ~G2 & G4 ;
  assign n438 = n436 & n437 ;
  assign n439 = G20 & n395 ;
  assign n440 = ~G8 & n392 ;
  assign n441 = G19 & ~n398 ;
  assign n442 = n440 | n441 ;
  assign n443 = n439 | n442 ;
  assign n444 = G7 | n407 ;
  assign n445 = G18 & ~n401 ;
  assign n446 = ~G21 & G9 ;
  assign n447 = n385 | n446 ;
  assign n448 = ~n445 & n447 ;
  assign n449 = ~n419 & n448 ;
  assign n450 = n444 & n449 ;
  assign n451 = ~n443 & n450 ;
  assign n452 = G40 & n395 ;
  assign n453 = n420 | n452 ;
  assign n454 = G41 & ~n398 ;
  assign n455 = G11 & ~G39 ;
  assign n456 = n385 | n455 ;
  assign n457 = ~n454 & n456 ;
  assign n458 = ~n453 & n457 ;
  assign n459 = G13 | n407 ;
  assign n460 = G14 & ~G42 ;
  assign n461 = n401 | n460 ;
  assign n462 = G4 & n461 ;
  assign n463 = n459 & n462 ;
  assign n464 = n458 & n463 ;
  assign n465 = n451 | n464 ;
  assign n466 = ~n381 & n465 ;
  assign n467 = n379 & ~n466 ;
  assign n468 = ~n438 & n467 ;
  assign n469 = n314 | n337 ;
  assign n470 = G24 | n265 ;
  assign n471 = n469 | n470 ;
  assign n472 = n293 | n471 ;
  assign n473 = n315 & n338 ;
  assign n474 = G24 & n265 ;
  assign n475 = n293 & n474 ;
  assign n476 = n473 & n475 ;
  assign n477 = n472 & ~n476 ;
  assign n478 = n361 | n477 ;
  assign n479 = n344 & n361 ;
  assign n480 = n478 & ~n479 ;
  assign n481 = G47 & ~n480 ;
  assign n482 = ~n374 & n436 ;
  assign n483 = ~n215 & n374 ;
  assign n484 = n482 | n483 ;
  assign n485 = n481 | n484 ;
  assign n486 = n481 & n484 ;
  assign n487 = n379 | n486 ;
  assign n488 = n485 & ~n487 ;
  assign n489 = n468 | n488 ;
  assign n490 = G47 & n480 ;
  assign n491 = n224 & n361 ;
  assign n492 = n238 & ~n491 ;
  assign n493 = ~n238 & n491 ;
  assign n494 = n492 | n493 ;
  assign n495 = n436 & n494 ;
  assign n496 = G27 & ~n77 ;
  assign n497 = n176 & n496 ;
  assign n498 = n190 | n497 ;
  assign n499 = n190 & n497 ;
  assign n500 = n498 & ~n499 ;
  assign n501 = n495 & n500 ;
  assign n502 = n240 & n501 ;
  assign n503 = n240 | n501 ;
  assign n504 = ~n502 & n503 ;
  assign n505 = n490 & ~n504 ;
  assign n506 = n240 | n374 ;
  assign n507 = ~n358 & n506 ;
  assign n508 = n237 & ~n361 ;
  assign n509 = n214 & ~n361 ;
  assign n510 = n494 & ~n509 ;
  assign n511 = n508 | n510 ;
  assign n512 = n500 & n511 ;
  assign n513 = n189 & ~n496 ;
  assign n514 = n512 | n513 ;
  assign n515 = n507 & n514 ;
  assign n516 = n507 | n514 ;
  assign n517 = ~n515 & n516 ;
  assign n518 = n505 & n517 ;
  assign n519 = n505 | n517 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = G1 | G2 ;
  assign n522 = n56 & n521 ;
  assign n523 = ~n520 & n522 ;
  assign n524 = G7 & ~G9 ;
  assign n525 = n52 | n105 ;
  assign n526 = ~n524 & n525 ;
  assign n527 = n521 | n526 ;
  assign n528 = ~G14 & n74 ;
  assign n529 = ~n275 & n528 ;
  assign n530 = n527 & ~n529 ;
  assign n531 = n523 | ~n530 ;
  assign n532 = ~n125 & n260 ;
  assign n533 = ~n73 & n532 ;
  assign n534 = n340 & ~n361 ;
  assign n535 = n365 | n534 ;
  assign n536 = n320 & n534 ;
  assign n537 = n535 & ~n536 ;
  assign n538 = n428 | n537 ;
  assign n539 = n428 & n537 ;
  assign n540 = n538 & ~n539 ;
  assign n541 = n374 & n540 ;
  assign n542 = n372 | n541 ;
  assign n543 = n282 & n361 ;
  assign n544 = n298 | n543 ;
  assign n545 = n298 & n543 ;
  assign n546 = n544 & ~n545 ;
  assign n547 = n317 & ~n361 ;
  assign n548 = n535 & ~n547 ;
  assign n549 = n546 | n548 ;
  assign n550 = n546 & n548 ;
  assign n551 = n549 & ~n550 ;
  assign n552 = ~n371 & n551 ;
  assign n553 = n371 & ~n551 ;
  assign n554 = n552 | n553 ;
  assign n555 = n374 & ~n554 ;
  assign n556 = n542 | n555 ;
  assign n557 = ~n533 & n556 ;
  assign n558 = n295 & ~n361 ;
  assign n559 = n549 & ~n558 ;
  assign n560 = n254 & n361 ;
  assign n561 = n270 | n560 ;
  assign n562 = n270 & n560 ;
  assign n563 = n561 & ~n562 ;
  assign n564 = n559 & ~n563 ;
  assign n565 = ~n559 & n563 ;
  assign n566 = n564 | n565 ;
  assign n567 = n553 & ~n566 ;
  assign n568 = ~n553 & n566 ;
  assign n569 = n567 | n568 ;
  assign n570 = ~n557 & n569 ;
  assign n571 = n377 & n563 ;
  assign n572 = ~G19 & G7 ;
  assign n573 = n401 | n572 ;
  assign n574 = G21 & n395 ;
  assign n575 = G20 & ~n398 ;
  assign n576 = n574 | n575 ;
  assign n577 = n573 & ~n576 ;
  assign n578 = G10 & ~G22 ;
  assign n579 = n385 | n578 ;
  assign n580 = n577 & n579 ;
  assign n581 = ~G9 & n392 ;
  assign n582 = G8 | n407 ;
  assign n583 = ~n581 & n582 ;
  assign n584 = ~G4 & n583 ;
  assign n585 = n580 & n584 ;
  assign n586 = n386 & ~n401 ;
  assign n587 = G12 & ~G40 ;
  assign n588 = n385 | n587 ;
  assign n589 = ~n586 & n588 ;
  assign n590 = G42 & ~n398 ;
  assign n591 = G41 & n395 ;
  assign n592 = n590 | n591 ;
  assign n593 = G14 | n407 ;
  assign n594 = ~G13 & n392 ;
  assign n595 = G4 & ~n594 ;
  assign n596 = n593 & n595 ;
  assign n597 = ~n592 & n596 ;
  assign n598 = n589 & n597 ;
  assign n599 = n585 | n598 ;
  assign n600 = ~n381 & n599 ;
  assign n601 = n379 & ~n600 ;
  assign n602 = ~n571 & n601 ;
  assign n603 = n570 | n602 ;
  assign n604 = n374 | n540 ;
  assign n605 = ~n542 & n604 ;
  assign n606 = n533 & ~n540 ;
  assign n607 = n365 & n377 ;
  assign n608 = G39 & n392 ;
  assign n609 = G44 & ~n398 ;
  assign n610 = n608 | n609 ;
  assign n611 = n399 & ~n401 ;
  assign n612 = G43 & n395 ;
  assign n613 = n611 | n612 ;
  assign n614 = n610 | n613 ;
  assign n615 = G40 & ~n407 ;
  assign n616 = n385 | n460 ;
  assign n617 = G4 & n616 ;
  assign n618 = ~n615 & n617 ;
  assign n619 = ~n614 & n618 ;
  assign n620 = ~G7 & n395 ;
  assign n621 = G22 & ~n398 ;
  assign n622 = n620 | n621 ;
  assign n623 = G12 | n385 ;
  assign n624 = G9 | n401 ;
  assign n625 = n623 & n624 ;
  assign n626 = ~n622 & n625 ;
  assign n627 = G10 | n407 ;
  assign n628 = G8 | n385 ;
  assign n629 = ~G4 & n628 ;
  assign n630 = ~G11 & n392 ;
  assign n631 = G21 & ~n401 ;
  assign n632 = n630 | n631 ;
  assign n633 = n629 & ~n632 ;
  assign n634 = n627 & n633 ;
  assign n635 = n626 & n634 ;
  assign n636 = n619 | n635 ;
  assign n637 = ~n381 & n636 ;
  assign n638 = n379 & ~n637 ;
  assign n639 = ~n607 & n638 ;
  assign n640 = n606 | n639 ;
  assign n641 = n605 | n640 ;
  assign n642 = ~n372 & n604 ;
  assign n643 = ~n554 & n642 ;
  assign n644 = n377 & n546 ;
  assign n645 = G21 & ~n398 ;
  assign n646 = G8 | n401 ;
  assign n647 = G11 & G7 ;
  assign n648 = n385 | n647 ;
  assign n649 = n646 & n648 ;
  assign n650 = ~n645 & n649 ;
  assign n651 = G9 | n407 ;
  assign n652 = G20 & ~n401 ;
  assign n653 = G4 | n652 ;
  assign n654 = ~G10 & n392 ;
  assign n655 = G22 & n395 ;
  assign n656 = n654 | n655 ;
  assign n657 = n653 | n656 ;
  assign n658 = n651 & ~n657 ;
  assign n659 = n650 & n658 ;
  assign n660 = G42 & n395 ;
  assign n661 = G40 | G44 ;
  assign n662 = ~n401 & n661 ;
  assign n663 = n660 | n662 ;
  assign n664 = G43 & ~n398 ;
  assign n665 = ~G14 & n392 ;
  assign n666 = n664 | n665 ;
  assign n667 = n663 | n666 ;
  assign n668 = G39 & ~n407 ;
  assign n669 = G13 & ~G41 ;
  assign n670 = n385 | n669 ;
  assign n671 = G4 & n670 ;
  assign n672 = ~n668 & n671 ;
  assign n673 = ~n667 & n672 ;
  assign n674 = n659 | n673 ;
  assign n675 = ~n381 & n674 ;
  assign n676 = n379 & ~n675 ;
  assign n677 = ~n644 & n676 ;
  assign n678 = n372 | n604 ;
  assign n679 = ~n533 & n678 ;
  assign n680 = n554 & ~n679 ;
  assign n681 = n677 | n680 ;
  assign n682 = n643 | n681 ;
  assign n683 = n490 & n501 ;
  assign n684 = n490 & n495 ;
  assign n685 = n500 | n511 ;
  assign n686 = ~n512 & n685 ;
  assign n687 = ~n684 & n686 ;
  assign n688 = n683 | n687 ;
  assign n689 = n482 | n509 ;
  assign n690 = n436 & n490 ;
  assign n691 = n494 | n690 ;
  assign n692 = ~n684 & n691 ;
  assign n693 = n689 | n692 ;
  assign n694 = n689 & n692 ;
  assign n695 = n693 & ~n694 ;
  assign n696 = n490 & ~n507 ;
  assign n697 = n695 | n696 ;
  assign n698 = n372 | n697 ;
  assign n699 = ~n533 & n698 ;
  assign n700 = n688 & ~n699 ;
  assign n701 = ~n372 & n697 ;
  assign n702 = ~n688 & n701 ;
  assign n703 = n437 & n500 ;
  assign n704 = n401 | n587 ;
  assign n705 = n408 & n704 ;
  assign n706 = ~G14 & n395 ;
  assign n707 = n411 & ~n654 ;
  assign n708 = ~n706 & n707 ;
  assign n709 = G39 & ~n398 ;
  assign n710 = G4 & n409 ;
  assign n711 = ~n709 & n710 ;
  assign n712 = n708 & n711 ;
  assign n713 = n705 & n712 ;
  assign n714 = G16 & ~n401 ;
  assign n715 = G17 & ~n398 ;
  assign n716 = G22 & n392 ;
  assign n717 = n715 | n716 ;
  assign n718 = n714 | n717 ;
  assign n719 = G21 & ~n407 ;
  assign n720 = G18 & n395 ;
  assign n721 = n385 | n572 ;
  assign n722 = ~n720 & n721 ;
  assign n723 = ~n719 & n722 ;
  assign n724 = ~n653 & n723 ;
  assign n725 = ~n718 & n724 ;
  assign n726 = n713 | n725 ;
  assign n727 = ~n381 & n726 ;
  assign n728 = n379 & ~n727 ;
  assign n729 = ~n703 & n728 ;
  assign n730 = n702 | n729 ;
  assign n731 = n700 | n730 ;
  assign n732 = n142 & n496 ;
  assign n733 = n165 | n732 ;
  assign n734 = n165 & n732 ;
  assign n735 = n733 & ~n734 ;
  assign n736 = n437 & n735 ;
  assign n737 = G18 | G22 ;
  assign n738 = ~n385 & n737 ;
  assign n739 = G16 & ~n398 ;
  assign n740 = G20 & ~n407 ;
  assign n741 = n739 | n740 ;
  assign n742 = G17 & n395 ;
  assign n743 = G15 | G19 ;
  assign n744 = ~n401 & n743 ;
  assign n745 = n742 | n744 ;
  assign n746 = G21 & n392 ;
  assign n747 = n146 & ~n746 ;
  assign n748 = ~n745 & n747 ;
  assign n749 = ~n741 & n748 ;
  assign n750 = ~n738 & n749 ;
  assign n751 = G5 & n627 ;
  assign n752 = G14 | n398 ;
  assign n753 = ~n581 & n752 ;
  assign n754 = ~G13 & n395 ;
  assign n755 = n623 & ~n754 ;
  assign n756 = n753 & n755 ;
  assign n757 = n401 | n455 ;
  assign n758 = n629 & n757 ;
  assign n759 = n756 & n758 ;
  assign n760 = n751 & n759 ;
  assign n761 = n750 | n760 ;
  assign n762 = ~n381 & n761 ;
  assign n763 = n379 & ~n762 ;
  assign n764 = ~n736 & n763 ;
  assign n765 = n695 & n696 ;
  assign n766 = ~n688 & n696 ;
  assign n767 = n372 | n766 ;
  assign n768 = n765 | n767 ;
  assign n769 = ~n533 & n768 ;
  assign n770 = n514 & ~n735 ;
  assign n771 = ~n514 & n735 ;
  assign n772 = n770 | n771 ;
  assign n773 = n683 & ~n772 ;
  assign n774 = ~n683 & n772 ;
  assign n775 = n773 | n774 ;
  assign n776 = ~n769 & n775 ;
  assign n777 = n764 | n776 ;
  assign n778 = n701 & ~n765 ;
  assign n779 = n437 & n494 ;
  assign n780 = G39 & n395 ;
  assign n781 = G40 & ~n398 ;
  assign n782 = n780 | n781 ;
  assign n783 = G10 & G14 ;
  assign n784 = n385 | n783 ;
  assign n785 = ~n630 & n784 ;
  assign n786 = ~n782 & n785 ;
  assign n787 = G12 | n407 ;
  assign n788 = n401 | n669 ;
  assign n789 = G4 & n788 ;
  assign n790 = n787 & n789 ;
  assign n791 = n786 & n790 ;
  assign n792 = G17 & ~n401 ;
  assign n793 = G19 & n395 ;
  assign n794 = n631 | n793 ;
  assign n795 = n792 | n794 ;
  assign n796 = ~n398 & n737 ;
  assign n797 = n171 | n796 ;
  assign n798 = ~G7 & n392 ;
  assign n799 = G20 & ~n385 ;
  assign n800 = n798 | n799 ;
  assign n801 = n797 | n800 ;
  assign n802 = n629 & ~n801 ;
  assign n803 = ~n795 & n802 ;
  assign n804 = n791 | n803 ;
  assign n805 = ~n381 & n804 ;
  assign n806 = n379 & ~n805 ;
  assign n807 = ~n779 & n806 ;
  assign n808 = n533 & ~n695 ;
  assign n809 = n807 | n808 ;
  assign n810 = n778 | n809 ;
  assign n811 = n731 | n777 ;
  assign n812 = n489 | n810 ;
  assign n813 = n603 | n682 ;
  assign n814 = n432 & ~n641 ;
  assign n815 = ~n813 & n814 ;
  assign n816 = ~n812 & n815 ;
  assign n817 = n811 | ~n816 ;
  assign n818 = G48 & ~n811 ;
  assign n819 = G27 & ~n817 ;
  assign n820 = n818 | ~n819 ;
  assign n821 = n489 & n810 ;
  assign n822 = n812 & ~n821 ;
  assign n823 = ~n432 & n641 ;
  assign n824 = n814 | n823 ;
  assign n825 = n603 & n682 ;
  assign n826 = n813 & ~n825 ;
  assign n827 = n824 | n826 ;
  assign n828 = n824 & n826 ;
  assign n829 = n827 & ~n828 ;
  assign n830 = n822 & n829 ;
  assign n831 = n822 | n829 ;
  assign n832 = ~n830 & n831 ;
  assign n833 = n731 & n777 ;
  assign n834 = n811 & ~n833 ;
  assign n835 = G50 & n834 ;
  assign n836 = G50 | n834 ;
  assign n837 = ~n360 & n836 ;
  assign n838 = ~n835 & n837 ;
  assign n839 = n832 & n838 ;
  assign n840 = n832 | n838 ;
  assign n841 = n839 | ~n840 ;
  assign n842 = n832 | n834 ;
  assign n843 = n832 & n834 ;
  assign n844 = n842 & ~n843 ;
  assign G3519 = n53 ;
  assign G3520 = n55 ;
  assign G3521 = n82 ;
  assign G3522 = n103 ;
  assign G3523 = n122 ;
  assign G3524 = n345 ;
  assign G3525 = n359 ;
  assign G3526 = n371 ;
  assign G3527 = n376 ;
  assign G3528 = n432 ;
  assign G3529 = n489 ;
  assign G3530 = n531 ;
  assign G3531 = n603 ;
  assign G3532 = n641 ;
  assign G3533 = n682 ;
  assign G3534 = n731 ;
  assign G3535 = n777 ;
  assign G3536 = n810 ;
  assign G3537 = n817 ;
  assign G3538 = n820 ;
  assign G3539 = n841 ;
  assign G3540 = n844 ;
endmodule