module counter_128 ( in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ , out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ );
  input in_18_ , in_1_ , in_7_ , in_109_ , in_13_ , in_106_ , in_54_ , in_118_ , in_101_ , in_3_ , in_0_ , in_113_ , in_56_ , in_30_ , in_89_ , in_35_ , in_70_ , in_38_ , in_100_ , in_105_ , in_28_ , in_10_ , in_9_ , in_78_ , in_29_ , in_60_ , in_94_ , in_108_ , in_117_ , in_103_ , in_67_ , in_44_ , in_57_ , in_76_ , in_47_ , in_20_ , in_84_ , in_17_ , in_72_ , in_116_ , in_16_ , in_120_ , in_104_ , in_64_ , in_125_ , in_58_ , in_42_ , in_40_ , in_81_ , in_115_ , in_88_ , in_24_ , in_33_ , in_123_ , in_61_ , in_79_ , in_31_ , in_36_ , in_82_ , in_111_ , in_68_ , in_2_ , in_87_ , in_74_ , in_114_ , in_53_ , in_83_ , in_86_ , in_65_ , in_102_ , in_6_ , in_75_ , in_4_ , in_93_ , in_45_ , in_90_ , in_80_ , in_73_ , in_46_ , in_25_ , in_107_ , in_37_ , in_85_ , in_49_ , in_39_ , in_63_ , in_12_ , in_112_ , in_32_ , in_119_ , in_77_ , in_34_ , in_41_ , in_122_ , in_124_ , in_48_ , in_92_ , in_15_ , in_55_ , in_50_ , in_5_ , in_127_ , in_96_ , in_22_ , in_43_ , in_52_ , in_51_ , in_21_ , in_95_ , in_59_ , in_69_ , in_121_ , in_97_ , in_11_ , in_98_ , in_126_ , in_14_ , in_91_ , in_26_ , in_99_ , in_27_ , in_71_ , in_8_ , in_23_ , in_110_ , in_62_ , in_66_ , in_19_ ;
  output out_3_ , out_2_ , out_5_ , out_1_ , out_0_ , out_7_ , out_4_ , out_6_ ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 ;
  assign n129 = in_127_ & in_126_ ;
  assign n130 = in_125_ | in_124_ ;
  assign n131 = in_117_ | in_116_ ;
  assign n132 = in_113_ | in_112_ ;
  assign n133 = in_115_ & in_114_ ;
  assign n134 = ( n131 & n132 ) | ( n131 & n133 ) | ( n132 & n133 ) ;
  assign n135 = ( ~n131 & n132 ) | ( ~n131 & n133 ) | ( n132 & n133 ) ;
  assign n136 = ( n131 & ~n134 ) | ( n131 & n135 ) | ( ~n134 & n135 ) ;
  assign n137 = in_123_ & in_122_ ;
  assign n138 = in_118_ & in_119_ ;
  assign n139 = in_120_ | in_121_ ;
  assign n140 = ( n137 & n138 ) | ( n137 & n139 ) | ( n138 & n139 ) ;
  assign n141 = ( ~n137 & n138 ) | ( ~n137 & n139 ) | ( n138 & n139 ) ;
  assign n142 = ( n137 & ~n140 ) | ( n137 & n141 ) | ( ~n140 & n141 ) ;
  assign n143 = ( n130 & n136 ) | ( n130 & n142 ) | ( n136 & n142 ) ;
  assign n144 = ( ~n130 & n136 ) | ( ~n130 & n142 ) | ( n136 & n142 ) ;
  assign n145 = ( n130 & ~n143 ) | ( n130 & n144 ) | ( ~n143 & n144 ) ;
  assign n146 = n129 & n145 ;
  assign n147 = n129 | n145 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = in_111_ & in_110_ ;
  assign n150 = in_109_ | in_108_ ;
  assign n151 = in_101_ | in_100_ ;
  assign n152 = in_96_ | in_97_ ;
  assign n153 = in_98_ & in_99_ ;
  assign n154 = ( ~n151 & n152 ) | ( ~n151 & n153 ) | ( n152 & n153 ) ;
  assign n155 = ( n151 & n152 ) | ( n151 & n153 ) | ( n152 & n153 ) ;
  assign n156 = ( n151 & n154 ) | ( n151 & ~n155 ) | ( n154 & ~n155 ) ;
  assign n157 = in_106_ & in_107_ ;
  assign n158 = in_103_ & in_102_ ;
  assign n159 = in_105_ | in_104_ ;
  assign n160 = ( n157 & n158 ) | ( n157 & n159 ) | ( n158 & n159 ) ;
  assign n161 = ( ~n157 & n158 ) | ( ~n157 & n159 ) | ( n158 & n159 ) ;
  assign n162 = ( n157 & ~n160 ) | ( n157 & n161 ) | ( ~n160 & n161 ) ;
  assign n163 = ( n150 & n156 ) | ( n150 & n162 ) | ( n156 & n162 ) ;
  assign n164 = ( ~n150 & n156 ) | ( ~n150 & n162 ) | ( n156 & n162 ) ;
  assign n165 = ( n150 & ~n163 ) | ( n150 & n164 ) | ( ~n163 & n164 ) ;
  assign n166 = n149 & n165 ;
  assign n167 = n149 | n165 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = n148 & n168 ;
  assign n170 = n148 | n168 ;
  assign n171 = ~n169 & n170 ;
  assign n172 = in_94_ & in_95_ ;
  assign n173 = in_93_ | in_92_ ;
  assign n174 = in_84_ | in_85_ ;
  assign n175 = in_81_ | in_80_ ;
  assign n176 = in_82_ & in_83_ ;
  assign n177 = ( n174 & n175 ) | ( n174 & n176 ) | ( n175 & n176 ) ;
  assign n178 = ( ~n174 & n175 ) | ( ~n174 & n176 ) | ( n175 & n176 ) ;
  assign n179 = ( n174 & ~n177 ) | ( n174 & n178 ) | ( ~n177 & n178 ) ;
  assign n180 = in_90_ & in_91_ ;
  assign n181 = in_87_ & in_86_ ;
  assign n182 = in_89_ | in_88_ ;
  assign n183 = ( n180 & n181 ) | ( n180 & n182 ) | ( n181 & n182 ) ;
  assign n184 = ( ~n180 & n181 ) | ( ~n180 & n182 ) | ( n181 & n182 ) ;
  assign n185 = ( n180 & ~n183 ) | ( n180 & n184 ) | ( ~n183 & n184 ) ;
  assign n186 = ( n173 & n179 ) | ( n173 & n185 ) | ( n179 & n185 ) ;
  assign n187 = ( ~n173 & n179 ) | ( ~n173 & n185 ) | ( n179 & n185 ) ;
  assign n188 = ( n173 & ~n186 ) | ( n173 & n187 ) | ( ~n186 & n187 ) ;
  assign n189 = n172 & n188 ;
  assign n190 = n172 | n188 ;
  assign n191 = ~n189 & n190 ;
  assign n192 = in_78_ & in_79_ ;
  assign n193 = in_76_ | in_77_ ;
  assign n194 = in_68_ | in_69_ ;
  assign n195 = in_64_ | in_65_ ;
  assign n196 = in_67_ & in_66_ ;
  assign n197 = ( n194 & n195 ) | ( n194 & n196 ) | ( n195 & n196 ) ;
  assign n198 = ( ~n194 & n195 ) | ( ~n194 & n196 ) | ( n195 & n196 ) ;
  assign n199 = ( n194 & ~n197 ) | ( n194 & n198 ) | ( ~n197 & n198 ) ;
  assign n200 = in_74_ & in_75_ ;
  assign n201 = in_70_ & in_71_ ;
  assign n202 = in_72_ | in_73_ ;
  assign n203 = ( n200 & n201 ) | ( n200 & n202 ) | ( n201 & n202 ) ;
  assign n204 = ( ~n200 & n201 ) | ( ~n200 & n202 ) | ( n201 & n202 ) ;
  assign n205 = ( n200 & ~n203 ) | ( n200 & n204 ) | ( ~n203 & n204 ) ;
  assign n206 = ( n193 & n199 ) | ( n193 & n205 ) | ( n199 & n205 ) ;
  assign n207 = ( ~n193 & n199 ) | ( ~n193 & n205 ) | ( n199 & n205 ) ;
  assign n208 = ( n193 & ~n206 ) | ( n193 & n207 ) | ( ~n206 & n207 ) ;
  assign n209 = n192 & n208 ;
  assign n210 = n192 | n208 ;
  assign n211 = ~n209 & n210 ;
  assign n212 = n191 & n211 ;
  assign n213 = n191 | n211 ;
  assign n214 = ~n212 & n213 ;
  assign n215 = n171 & n214 ;
  assign n216 = ( n134 & n140 ) | ( n134 & n143 ) | ( n140 & n143 ) ;
  assign n217 = ( n134 & n140 ) | ( n134 & ~n143 ) | ( n140 & ~n143 ) ;
  assign n218 = ( n143 & ~n216 ) | ( n143 & n217 ) | ( ~n216 & n217 ) ;
  assign n219 = n146 & n218 ;
  assign n220 = n146 | n218 ;
  assign n221 = ~n219 & n220 ;
  assign n222 = ( n155 & n160 ) | ( n155 & n163 ) | ( n160 & n163 ) ;
  assign n223 = ( n155 & n160 ) | ( n155 & ~n163 ) | ( n160 & ~n163 ) ;
  assign n224 = ( n163 & ~n222 ) | ( n163 & n223 ) | ( ~n222 & n223 ) ;
  assign n225 = n166 & n224 ;
  assign n226 = n166 | n224 ;
  assign n227 = ~n225 & n226 ;
  assign n228 = n221 & n227 ;
  assign n229 = n221 | n227 ;
  assign n230 = ~n228 & n229 ;
  assign n231 = n169 & n230 ;
  assign n232 = n169 | n230 ;
  assign n233 = ~n231 & n232 ;
  assign n234 = ( n177 & n183 ) | ( n177 & n186 ) | ( n183 & n186 ) ;
  assign n235 = ( n177 & n183 ) | ( n177 & ~n186 ) | ( n183 & ~n186 ) ;
  assign n236 = ( n186 & ~n234 ) | ( n186 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = n189 & n236 ;
  assign n238 = n189 | n236 ;
  assign n239 = ~n237 & n238 ;
  assign n240 = ( n197 & n203 ) | ( n197 & n206 ) | ( n203 & n206 ) ;
  assign n241 = ( n197 & n203 ) | ( n197 & ~n206 ) | ( n203 & ~n206 ) ;
  assign n242 = ( n206 & ~n240 ) | ( n206 & n241 ) | ( ~n240 & n241 ) ;
  assign n243 = n209 & n242 ;
  assign n244 = n209 | n242 ;
  assign n245 = ~n243 & n244 ;
  assign n246 = n239 & n245 ;
  assign n247 = n239 | n245 ;
  assign n248 = ~n246 & n247 ;
  assign n249 = n212 & n248 ;
  assign n250 = n212 | n248 ;
  assign n251 = ~n249 & n250 ;
  assign n252 = n233 & n251 ;
  assign n253 = n233 | n251 ;
  assign n254 = ~n252 & n253 ;
  assign n255 = n215 & n254 ;
  assign n256 = n215 | n254 ;
  assign n257 = ~n255 & n256 ;
  assign n258 = n171 | n214 ;
  assign n259 = ~n215 & n258 ;
  assign n260 = in_30_ & in_31_ ;
  assign n261 = in_28_ | in_29_ ;
  assign n262 = in_26_ & in_27_ ;
  assign n263 = in_22_ & in_23_ ;
  assign n264 = in_24_ | in_25_ ;
  assign n265 = ( n262 & n263 ) | ( n262 & n264 ) | ( n263 & n264 ) ;
  assign n266 = ( ~n262 & n263 ) | ( ~n262 & n264 ) | ( n263 & n264 ) ;
  assign n267 = ( n262 & ~n265 ) | ( n262 & n266 ) | ( ~n265 & n266 ) ;
  assign n268 = in_20_ | in_21_ ;
  assign n269 = in_17_ | in_16_ ;
  assign n270 = in_18_ & in_19_ ;
  assign n271 = ( n268 & n269 ) | ( n268 & n270 ) | ( n269 & n270 ) ;
  assign n272 = ( ~n268 & n269 ) | ( ~n268 & n270 ) | ( n269 & n270 ) ;
  assign n273 = ( n268 & ~n271 ) | ( n268 & n272 ) | ( ~n271 & n272 ) ;
  assign n274 = ( n261 & n267 ) | ( n261 & n273 ) | ( n267 & n273 ) ;
  assign n275 = ( ~n261 & n267 ) | ( ~n261 & n273 ) | ( n267 & n273 ) ;
  assign n276 = ( n261 & ~n274 ) | ( n261 & n275 ) | ( ~n274 & n275 ) ;
  assign n277 = n260 & n276 ;
  assign n278 = n260 | n276 ;
  assign n279 = ~n277 & n278 ;
  assign n280 = in_15_ & in_14_ ;
  assign n281 = in_13_ | in_12_ ;
  assign n282 = in_4_ | in_5_ ;
  assign n283 = in_1_ | in_0_ ;
  assign n284 = in_3_ & in_2_ ;
  assign n285 = ( n282 & n283 ) | ( n282 & n284 ) | ( n283 & n284 ) ;
  assign n286 = ( ~n282 & n283 ) | ( ~n282 & n284 ) | ( n283 & n284 ) ;
  assign n287 = ( n282 & ~n285 ) | ( n282 & n286 ) | ( ~n285 & n286 ) ;
  assign n288 = in_10_ & in_11_ ;
  assign n289 = in_7_ & in_6_ ;
  assign n290 = in_9_ | in_8_ ;
  assign n291 = ( n288 & n289 ) | ( n288 & n290 ) | ( n289 & n290 ) ;
  assign n292 = ( ~n288 & n289 ) | ( ~n288 & n290 ) | ( n289 & n290 ) ;
  assign n293 = ( n288 & ~n291 ) | ( n288 & n292 ) | ( ~n291 & n292 ) ;
  assign n294 = ( n281 & n287 ) | ( n281 & n293 ) | ( n287 & n293 ) ;
  assign n295 = ( ~n281 & n287 ) | ( ~n281 & n293 ) | ( n287 & n293 ) ;
  assign n296 = ( n281 & ~n294 ) | ( n281 & n295 ) | ( ~n294 & n295 ) ;
  assign n297 = n280 & n296 ;
  assign n298 = n280 | n296 ;
  assign n299 = ~n297 & n298 ;
  assign n300 = n279 & n299 ;
  assign n301 = n279 | n299 ;
  assign n302 = ~n300 & n301 ;
  assign n303 = in_47_ & in_46_ ;
  assign n304 = in_44_ | in_45_ ;
  assign n305 = in_36_ | in_37_ ;
  assign n306 = in_33_ | in_32_ ;
  assign n307 = in_35_ & in_34_ ;
  assign n308 = ( n305 & n306 ) | ( n305 & n307 ) | ( n306 & n307 ) ;
  assign n309 = ( ~n305 & n306 ) | ( ~n305 & n307 ) | ( n306 & n307 ) ;
  assign n310 = ( n305 & ~n308 ) | ( n305 & n309 ) | ( ~n308 & n309 ) ;
  assign n311 = in_42_ & in_43_ ;
  assign n312 = in_38_ & in_39_ ;
  assign n313 = in_40_ | in_41_ ;
  assign n314 = ( n311 & n312 ) | ( n311 & n313 ) | ( n312 & n313 ) ;
  assign n315 = ( ~n311 & n312 ) | ( ~n311 & n313 ) | ( n312 & n313 ) ;
  assign n316 = ( n311 & ~n314 ) | ( n311 & n315 ) | ( ~n314 & n315 ) ;
  assign n317 = ( n304 & n310 ) | ( n304 & n316 ) | ( n310 & n316 ) ;
  assign n318 = ( ~n304 & n310 ) | ( ~n304 & n316 ) | ( n310 & n316 ) ;
  assign n319 = ( n304 & ~n317 ) | ( n304 & n318 ) | ( ~n317 & n318 ) ;
  assign n320 = n303 & n319 ;
  assign n321 = n303 | n319 ;
  assign n322 = ~n320 & n321 ;
  assign n323 = in_63_ & in_62_ ;
  assign n324 = in_60_ | in_61_ ;
  assign n325 = in_58_ & in_59_ ;
  assign n326 = in_54_ & in_55_ ;
  assign n327 = in_56_ | in_57_ ;
  assign n328 = ( n325 & n326 ) | ( n325 & n327 ) | ( n326 & n327 ) ;
  assign n329 = ( ~n325 & n326 ) | ( ~n325 & n327 ) | ( n326 & n327 ) ;
  assign n330 = ( n325 & ~n328 ) | ( n325 & n329 ) | ( ~n328 & n329 ) ;
  assign n331 = in_53_ | in_52_ ;
  assign n332 = in_49_ | in_48_ ;
  assign n333 = in_50_ & in_51_ ;
  assign n334 = ( n331 & n332 ) | ( n331 & n333 ) | ( n332 & n333 ) ;
  assign n335 = ( ~n331 & n332 ) | ( ~n331 & n333 ) | ( n332 & n333 ) ;
  assign n336 = ( n331 & ~n334 ) | ( n331 & n335 ) | ( ~n334 & n335 ) ;
  assign n337 = ( n324 & n330 ) | ( n324 & n336 ) | ( n330 & n336 ) ;
  assign n338 = ( ~n324 & n330 ) | ( ~n324 & n336 ) | ( n330 & n336 ) ;
  assign n339 = ( n324 & ~n337 ) | ( n324 & n338 ) | ( ~n337 & n338 ) ;
  assign n340 = n323 & n339 ;
  assign n341 = n323 | n339 ;
  assign n342 = ~n340 & n341 ;
  assign n343 = n322 | n342 ;
  assign n344 = n322 & n342 ;
  assign n345 = n343 & ~n344 ;
  assign n346 = n302 & n345 ;
  assign n347 = n302 | n345 ;
  assign n348 = ~n346 & n347 ;
  assign n349 = n259 & n348 ;
  assign n350 = ( n265 & n271 ) | ( n265 & n274 ) | ( n271 & n274 ) ;
  assign n351 = ( n265 & n271 ) | ( n265 & ~n274 ) | ( n271 & ~n274 ) ;
  assign n352 = ( n274 & ~n350 ) | ( n274 & n351 ) | ( ~n350 & n351 ) ;
  assign n353 = n277 | n352 ;
  assign n354 = n277 & n352 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = ( n285 & n291 ) | ( n285 & n294 ) | ( n291 & n294 ) ;
  assign n357 = ( n285 & n291 ) | ( n285 & ~n294 ) | ( n291 & ~n294 ) ;
  assign n358 = ( n294 & ~n356 ) | ( n294 & n357 ) | ( ~n356 & n357 ) ;
  assign n359 = n297 & n358 ;
  assign n360 = n297 | n358 ;
  assign n361 = ~n359 & n360 ;
  assign n362 = n355 & n361 ;
  assign n363 = n355 | n361 ;
  assign n364 = ~n362 & n363 ;
  assign n365 = n300 & n364 ;
  assign n366 = n300 | n364 ;
  assign n367 = ~n365 & n366 ;
  assign n368 = ( n328 & n334 ) | ( n328 & n337 ) | ( n334 & n337 ) ;
  assign n369 = ( n328 & n334 ) | ( n328 & ~n337 ) | ( n334 & ~n337 ) ;
  assign n370 = ( n337 & ~n368 ) | ( n337 & n369 ) | ( ~n368 & n369 ) ;
  assign n371 = n340 & n370 ;
  assign n372 = n340 | n370 ;
  assign n373 = ~n371 & n372 ;
  assign n374 = ( n308 & n314 ) | ( n308 & n317 ) | ( n314 & n317 ) ;
  assign n375 = ( n308 & n314 ) | ( n308 & ~n317 ) | ( n314 & ~n317 ) ;
  assign n376 = ( n317 & ~n374 ) | ( n317 & n375 ) | ( ~n374 & n375 ) ;
  assign n377 = n320 & n376 ;
  assign n378 = n320 | n376 ;
  assign n379 = ~n377 & n378 ;
  assign n380 = n373 & n379 ;
  assign n381 = n373 | n379 ;
  assign n382 = ~n380 & n381 ;
  assign n383 = n344 & n382 ;
  assign n384 = n344 | n382 ;
  assign n385 = ~n383 & n384 ;
  assign n386 = n367 & n385 ;
  assign n387 = n367 | n385 ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n346 & n388 ;
  assign n390 = n346 | n388 ;
  assign n391 = ~n389 & n390 ;
  assign n392 = ( n257 & n349 ) | ( n257 & n391 ) | ( n349 & n391 ) ;
  assign n393 = ( n346 & n367 ) | ( n346 & n385 ) | ( n367 & n385 ) ;
  assign n394 = ( n300 & n355 ) | ( n300 & n361 ) | ( n355 & n361 ) ;
  assign n395 = n350 & n354 ;
  assign n396 = n350 | n354 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = n356 & n359 ;
  assign n399 = n356 | n359 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = n397 & n400 ;
  assign n402 = n397 | n400 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = n394 & n403 ;
  assign n405 = n394 | n403 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = n374 & n377 ;
  assign n408 = n374 | n377 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = n368 & n371 ;
  assign n411 = n368 | n371 ;
  assign n412 = ~n410 & n411 ;
  assign n413 = n409 & n412 ;
  assign n414 = n409 | n412 ;
  assign n415 = ~n413 & n414 ;
  assign n416 = ( n344 & n373 ) | ( n344 & n379 ) | ( n373 & n379 ) ;
  assign n417 = n415 & n416 ;
  assign n418 = n415 | n416 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = n406 & n419 ;
  assign n421 = n406 | n419 ;
  assign n422 = ~n420 & n421 ;
  assign n423 = n393 & n422 ;
  assign n424 = n393 | n422 ;
  assign n425 = ~n423 & n424 ;
  assign n426 = ( n215 & n233 ) | ( n215 & n251 ) | ( n233 & n251 ) ;
  assign n427 = ( n169 & n221 ) | ( n169 & n227 ) | ( n221 & n227 ) ;
  assign n428 = n216 & n219 ;
  assign n429 = n216 | n219 ;
  assign n430 = ~n428 & n429 ;
  assign n431 = n222 & n225 ;
  assign n432 = n222 | n225 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = n430 & n433 ;
  assign n435 = n430 | n433 ;
  assign n436 = ~n434 & n435 ;
  assign n437 = n427 & n436 ;
  assign n438 = n427 | n436 ;
  assign n439 = ~n437 & n438 ;
  assign n440 = ( n212 & n239 ) | ( n212 & n245 ) | ( n239 & n245 ) ;
  assign n441 = n234 & n237 ;
  assign n442 = n234 | n237 ;
  assign n443 = ~n441 & n442 ;
  assign n444 = n240 & n243 ;
  assign n445 = n240 | n243 ;
  assign n446 = ~n444 & n445 ;
  assign n447 = n443 & n446 ;
  assign n448 = n443 | n446 ;
  assign n449 = ~n447 & n448 ;
  assign n450 = n440 & n449 ;
  assign n451 = n440 | n449 ;
  assign n452 = ~n450 & n451 ;
  assign n453 = n439 & n452 ;
  assign n454 = n439 | n452 ;
  assign n455 = ~n453 & n454 ;
  assign n456 = n426 & n455 ;
  assign n457 = n426 | n455 ;
  assign n458 = ~n456 & n457 ;
  assign n459 = n425 & n458 ;
  assign n460 = n425 | n458 ;
  assign n461 = ~n459 & n460 ;
  assign n462 = n392 & n461 ;
  assign n463 = n392 | n461 ;
  assign n464 = ~n462 & n463 ;
  assign n465 = n257 & n391 ;
  assign n466 = n257 | n391 ;
  assign n467 = ~n465 & n466 ;
  assign n468 = n349 & n467 ;
  assign n469 = n349 | n467 ;
  assign n470 = ~n468 & n469 ;
  assign n471 = ( n393 & n406 ) | ( n393 & n419 ) | ( n406 & n419 ) ;
  assign n472 = n395 & n398 ;
  assign n473 = n395 | n398 ;
  assign n474 = ~n472 & n473 ;
  assign n475 = ( n394 & n397 ) | ( n394 & n400 ) | ( n397 & n400 ) ;
  assign n476 = n474 & n475 ;
  assign n477 = n474 | n475 ;
  assign n478 = ~n476 & n477 ;
  assign n479 = n407 & n410 ;
  assign n480 = n407 | n410 ;
  assign n481 = ~n479 & n480 ;
  assign n482 = ( n409 & n412 ) | ( n409 & n416 ) | ( n412 & n416 ) ;
  assign n483 = n481 & n482 ;
  assign n484 = n481 | n482 ;
  assign n485 = ~n483 & n484 ;
  assign n486 = n478 & n485 ;
  assign n487 = n478 | n485 ;
  assign n488 = ~n486 & n487 ;
  assign n489 = n471 & n488 ;
  assign n490 = n471 | n488 ;
  assign n491 = ~n489 & n490 ;
  assign n492 = ( n392 & n425 ) | ( n392 & n458 ) | ( n425 & n458 ) ;
  assign n493 = n428 & n431 ;
  assign n494 = n428 | n431 ;
  assign n495 = ~n493 & n494 ;
  assign n496 = ( n427 & n430 ) | ( n427 & n433 ) | ( n430 & n433 ) ;
  assign n497 = n495 & n496 ;
  assign n498 = n495 | n496 ;
  assign n499 = ~n497 & n498 ;
  assign n500 = n441 & n444 ;
  assign n501 = n441 | n444 ;
  assign n502 = ~n500 & n501 ;
  assign n503 = ( n440 & n443 ) | ( n440 & n446 ) | ( n443 & n446 ) ;
  assign n504 = n502 & n503 ;
  assign n505 = n502 | n503 ;
  assign n506 = ~n504 & n505 ;
  assign n507 = n499 & n506 ;
  assign n508 = n499 | n506 ;
  assign n509 = ~n507 & n508 ;
  assign n510 = ( n426 & n439 ) | ( n426 & n452 ) | ( n439 & n452 ) ;
  assign n511 = n509 & n510 ;
  assign n512 = n509 | n510 ;
  assign n513 = ~n511 & n512 ;
  assign n514 = ( n491 & n492 ) | ( n491 & n513 ) | ( n492 & n513 ) ;
  assign n515 = ( n471 & n478 ) | ( n471 & n485 ) | ( n478 & n485 ) ;
  assign n516 = ( n395 & n398 ) | ( n395 & n475 ) | ( n398 & n475 ) ;
  assign n517 = ( n407 & n410 ) | ( n407 & n482 ) | ( n410 & n482 ) ;
  assign n518 = n516 & n517 ;
  assign n519 = n516 | n517 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = n515 & n520 ;
  assign n522 = n515 | n520 ;
  assign n523 = ~n521 & n522 ;
  assign n524 = ( n428 & n431 ) | ( n428 & n496 ) | ( n431 & n496 ) ;
  assign n525 = ( n441 & n444 ) | ( n441 & n503 ) | ( n444 & n503 ) ;
  assign n526 = n524 & n525 ;
  assign n527 = n524 | n525 ;
  assign n528 = ~n526 & n527 ;
  assign n529 = ( n499 & n506 ) | ( n499 & n510 ) | ( n506 & n510 ) ;
  assign n530 = n528 & n529 ;
  assign n531 = n528 | n529 ;
  assign n532 = ~n530 & n531 ;
  assign n533 = n523 & n532 ;
  assign n534 = n523 | n532 ;
  assign n535 = ~n533 & n534 ;
  assign n536 = n514 & n535 ;
  assign n537 = n514 | n535 ;
  assign n538 = ~n536 & n537 ;
  assign n539 = n259 | n348 ;
  assign n540 = ~n349 & n539 ;
  assign n541 = ( n515 & n516 ) | ( n515 & n517 ) | ( n516 & n517 ) ;
  assign n542 = ( n514 & n523 ) | ( n514 & n532 ) | ( n523 & n532 ) ;
  assign n543 = ( n524 & n525 ) | ( n524 & n529 ) | ( n525 & n529 ) ;
  assign n544 = ( n541 & n542 ) | ( n541 & n543 ) | ( n542 & n543 ) ;
  assign n545 = n491 & n513 ;
  assign n546 = n491 | n513 ;
  assign n547 = ~n545 & n546 ;
  assign n548 = n492 & n547 ;
  assign n549 = n492 | n547 ;
  assign n550 = ~n548 & n549 ;
  assign n551 = n541 & n543 ;
  assign n552 = n541 | n543 ;
  assign n553 = ~n551 & n552 ;
  assign n554 = n542 & n553 ;
  assign n555 = n542 | n553 ;
  assign n556 = ~n554 & n555 ;
  assign out_3_ = n464 ;
  assign out_2_ = n470 ;
  assign out_5_ = n538 ;
  assign out_1_ = n540 ;
  assign out_0_ = 1'b0 ;
  assign out_7_ = n544 ;
  assign out_4_ = n550 ;
  assign out_6_ = n556 ;
endmodule