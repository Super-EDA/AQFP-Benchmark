module c5315 (G1,G10,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G11,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G12,G120,G121,G122,G123,G124,G125,G126,G127,G128,G129,G13,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G14,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G15,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G16,G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G17,G170,G171,G172,G173,G174,G175,G176,G177,G178,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G6,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G7,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G8,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G9,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315);
  input G1,G10,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G11,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G12,G120,G121,G122,G123,G124,G125,G126,G127,G128,G129,G13,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G14,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G15,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G16,G160,G161,G162,G163,G164,G165,G166,G167,G168,G169,G17,G170,G171,G172,G173,G174,G175,G176,G177,G178,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G6,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G7,G70,G71,G72,G73,G74,G75,G76,G77,G78,G79,G8,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G9,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99;
  output G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315;
  wire _w_8986,_w_8985,_w_8983,_w_8978,_w_8974,_w_8972,_w_8971,_w_8963,_w_8961,_w_8956,_w_8955,_w_8952,_w_8951,_w_8948,_w_8947,_w_8943,_w_8941,_w_8936,_w_8935,_w_8928,_w_8925,_w_8924,_w_8922,_w_8921,_w_8920,_w_8918,_w_8913,_w_8903,_w_8901,_w_8896,_w_8893,_w_8888,_w_8887,_w_8886,_w_8881,_w_8879,_w_8877,_w_8876,_w_8875,_w_8874,_w_8873,_w_8872,_w_8870,_w_8868,_w_8866,_w_8865,_w_8863,_w_8861,_w_8859,_w_8858,_w_8856,_w_8852,_w_8851,_w_8850,_w_8849,_w_8844,_w_8838,_w_8836,_w_8835,_w_8834,_w_8831,_w_8828,_w_8827,_w_8826,_w_8823,_w_8822,_w_8817,_w_8816,_w_8813,_w_8810,_w_8806,_w_8805,_w_8804,_w_8799,_w_8797,_w_8794,_w_8793,_w_8792,_w_8790,_w_8788,_w_8787,_w_8786,_w_8783,_w_8781,_w_8777,_w_8776,_w_8772,_w_8771,_w_8770,_w_8769,_w_8768,_w_8764,_w_8763,_w_8758,_w_8751,_w_8748,_w_8744,_w_8743,_w_8740,_w_8738,_w_8732,_w_8730,_w_8728,_w_8727,_w_8721,_w_8720,_w_8719,_w_8718,_w_8717,_w_8709,_w_8708,_w_8789,_w_8707,_w_8706,_w_8700,_w_8692,_w_8691,_w_8690,_w_8689,_w_8688,_w_8686,_w_8681,_w_8679,_w_8675,_w_8672,_w_8671,_w_8668,_w_8664,_w_8745,_w_8663,_w_8659,_w_8653,_w_8929,_w_8651,_w_8650,_w_8649,_w_8648,_w_8647,_w_8644,_w_8643,_w_8641,_w_8639,_w_8637,_w_8634,_w_8726,_w_8633,_w_8632,_w_8631,_w_8629,_w_8627,_w_8623,_w_8622,_w_8621,_w_8620,_w_8619,_w_8613,_w_8612,_w_8611,_w_8609,_w_8606,_w_8605,_w_8601,_w_8600,_w_8597,_w_8596,_w_8595,_w_8594,_w_8592,_w_8590,_w_8589,_w_8584,_w_8581,_w_8580,_w_8578,_w_8577,_w_8573,_w_8567,_w_8564,_w_8563,_w_8559,_w_8556,_w_8553,_w_8552,_w_8547,_w_8546,_w_8543,_w_8541,_w_8538,_w_8536,_w_8535,_w_8533,_w_8529,_w_8969,_w_8528,_w_8527,_w_8526,_w_8525,_w_8524,_w_8522,_w_8518,_w_8516,_w_8515,_w_8514,_w_8511,_w_8510,_w_8508,_w_8507,_w_8506,_w_8569,_w_8505,_w_8504,_w_8503,_w_8502,_w_8499,_w_8498,_w_8497,_w_8493,_w_8485,_w_8484,_w_8482,_w_8479,_w_8478,_w_8477,_w_8473,_w_8469,_w_8468,_w_8466,_w_8464,_w_8461,_w_8458,_w_8457,_w_8455,_w_8453,_w_8451,_w_8446,_w_8445,_w_8438,_w_8431,_w_8427,_w_8426,_w_8424,_w_8421,_w_8419,_w_8415,_w_8414,_w_8410,_w_8406,_w_8402,_w_8401,_w_8398,_w_8396,_w_8393,_w_8392,_w_8387,_w_8386,_w_8385,_w_8383,_w_8381,_w_8380,_w_8377,_w_8953,_w_8376,_w_8375,_w_8374,_w_8371,_w_8367,_w_8359,_w_8358,_w_8354,_w_8353,_w_8351,_w_8348,_w_8347,_w_8423,_w_8346,_w_8910,_w_8341,_w_8340,_w_8339,_w_8338,_w_8765,_w_8334,_w_8333,_w_8331,_w_8329,_w_8327,_w_8325,_w_8323,_w_8320,_w_8418,_w_8318,_w_8315,_w_8314,_w_8312,_w_8311,_w_8413,_w_8310,_w_8308,_w_8307,_w_8303,_w_8302,_w_8296,_w_8293,_w_8291,_w_8289,_w_8572,_w_8286,_w_8283,_w_8736,_w_8279,_w_8276,_w_8275,_w_8274,_w_8273,_w_8272,_w_8271,_w_8269,_w_8300,_w_8267,_w_8266,_w_8265,_w_8264,_w_8684,_w_8262,_w_8261,_w_8260,_w_8259,_w_8258,_w_8257,_w_8256,_w_8255,_w_8737,_w_8254,_w_8890,_w_8253,_w_8250,_w_8249,_w_8247,_w_8391,_w_8245,_w_8244,_w_8243,_w_8242,_w_8239,_w_8238,_w_8234,_w_8233,_w_8232,_w_8231,_w_8228,_w_8226,_w_8224,_w_8223,_w_8222,_w_8220,_w_8550,_w_8218,_w_8212,_w_8211,_w_8208,_w_8204,_w_8198,_w_8193,_w_8192,_w_8191,_w_8190,_w_8188,_w_8660,_w_8181,_w_8179,_w_8178,_w_8177,_w_8174,_w_8173,_w_8905,_w_8171,_w_8163,_w_8160,_w_8491,_w_8159,_w_8158,_w_8156,_w_8155,_w_8154,_w_8153,_w_8152,_w_8382,_w_8149,_w_8147,_w_8143,_w_8196,_w_8140,_w_8135,_w_8305,_w_8134,_w_8132,_w_8130,_w_8129,_w_8125,_w_8119,_w_8117,_w_8294,_w_8115,_w_8113,_w_8112,_w_8111,_w_8110,_w_8108,_w_8101,_w_8099,_w_8097,_w_8096,_w_8092,_w_8090,_w_8089,_w_8087,_w_8084,_w_8082,_w_8080,_w_8079,_w_8270,_w_8078,_w_8076,_w_8906,_w_8074,_w_8070,_w_8065,_w_8062,_w_8059,_w_8057,_w_8475,_w_8055,_w_8676,_w_8054,_w_8053,_w_8966,_w_8066,_w_8052,_w_8049,_w_8041,_w_8040,_w_8038,_w_8037,_w_8033,_w_8031,_w_8025,_w_8023,_w_8022,_w_8021,_w_8020,_w_8019,_w_8018,_w_8016,_w_8014,_w_8013,_w_8004,_w_8001,_w_8625,_w_7999,_w_7998,_w_7997,_w_8741,_w_7992,_w_7990,_w_7989,_w_7987,_w_7986,_w_7985,_w_7981,_w_7980,_w_7978,_w_8586,_w_7977,_w_7976,_w_7975,_w_7974,_w_8091,_w_7972,_w_7968,_w_7965,_w_7964,_w_7963,_w_8862,_w_7962,_w_7960,_w_7959,_w_7957,_w_7956,_w_7955,_w_7953,_w_7954,_w_7952,_w_7951,_w_7950,_w_7947,_w_7945,_w_7942,_w_7941,_w_7939,_w_7931,_w_7929,_w_7925,_w_8420,_w_7924,_w_7919,_w_7918,_w_7915,_w_7912,_w_7911,_w_7910,_w_8072,_w_7909,_w_7908,_w_7906,_w_7905,_w_7904,_w_7900,_w_8105,_w_7897,_w_7896,_w_7895,_w_7892,_w_7891,_w_7887,_w_7886,_w_7885,_w_7883,_w_7882,_w_7880,_w_7878,_w_8448,_w_7877,_w_7874,_w_7871,_w_7869,_w_7867,_w_7865,_w_7961,_w_7864,_w_7861,_w_7860,_w_7857,_w_7855,_w_7853,_w_7851,_w_7850,_w_7848,_w_7847,_w_7846,_w_7845,_w_7844,_w_7840,_w_8742,_w_7839,_w_7838,_w_7837,_w_7832,_w_7831,_w_7830,_w_7828,_w_7827,_w_7823,_w_7820,_w_7819,_w_7818,_w_7817,_w_7814,_w_7813,_w_7808,_w_7807,_w_7806,_w_7804,_w_7803,_w_7802,_w_7800,_w_7792,_w_7788,_w_7787,_w_7786,_w_7784,_w_7783,_w_7782,_w_7781,_w_7780,_w_7776,_w_7773,_w_7772,_w_7771,_w_7769,_w_7768,_w_7767,_w_7766,_w_7764,_w_7761,_w_7760,_w_7759,_w_7758,_w_7756,_w_7752,_w_8460,_w_7750,_w_7748,_w_7747,_w_7746,_w_7739,_w_7735,_w_7751,_w_7733,_w_7732,_w_7731,_w_7730,_w_7729,_w_7727,_w_7726,_w_7725,_w_7723,_w_7719,_w_8045,_w_7718,_w_7715,_w_7712,_w_7709,_w_7704,_w_7701,_w_7698,_w_7695,_w_7693,_w_7692,_w_7691,_w_7690,_w_7688,_w_7687,_w_7684,_w_7683,_w_7682,_w_7681,_w_7678,_w_7675,_w_7674,_w_7669,_w_8801,_w_7667,_w_7666,_w_7661,_w_7659,_w_7657,_w_7656,_w_7655,_w_7653,_w_7651,_w_7650,_w_7648,_w_7647,_w_7641,_w_8313,_w_7639,_w_7638,_w_7633,_w_7632,_w_7631,_w_7630,_w_7629,_w_7628,_w_7627,_w_7619,_w_7618,_w_7616,_w_7613,_w_7611,_w_7607,_w_7606,_w_7598,_w_7596,_w_7593,_w_7589,_w_7588,_w_7586,_w_7583,_w_7582,_w_7580,_w_8853,_w_7578,_w_7575,_w_7574,_w_7573,_w_7572,_w_7570,_w_7566,_w_7565,_w_8699,_w_7564,_w_7563,_w_7557,_w_7556,_w_7555,_w_7552,_w_7551,_w_7549,_w_7543,_w_7542,_w_7539,_w_8452,_w_7537,_w_7535,_w_7534,_w_7533,_w_7531,_w_7529,_w_7526,_w_7518,_w_7516,_w_8395,_w_8126,_w_7515,_w_7513,_w_7510,_w_7508,_w_7507,_w_8968,_w_7506,_w_7505,_w_7502,_w_7499,_w_7497,_w_7495,_w_7490,_w_7487,_w_7485,_w_7484,_w_7995,_w_7480,_w_7478,_w_7473,_w_7471,_w_7465,_w_7464,_w_7463,_w_7462,_w_7461,_w_8009,_w_7459,_w_8361,_w_7456,_w_7452,_w_7451,_w_7450,_w_7446,_w_7444,_w_7438,_w_7437,_w_7434,_w_7431,_w_7429,_w_7428,_w_7424,_w_8210,_w_7423,_w_8297,_w_7421,_w_7420,_w_7416,_w_7415,_w_7612,_w_7408,_w_7407,_w_7406,_w_7404,_w_7403,_w_7402,_w_7399,_w_7397,_w_7395,_w_7393,_w_7392,_w_7386,_w_7385,_w_7384,_w_7381,_w_7380,_w_7378,_w_7377,_w_8011,_w_7376,_w_7375,_w_7374,_w_8120,_w_7371,_w_7370,_w_7365,_w_7362,_w_7360,_w_7359,_w_7357,_w_7351,_w_7350,_w_7344,_w_7343,_w_7342,_w_7339,_w_7337,_w_7336,_w_7335,_w_7331,_w_7330,_w_7329,_w_7449,_w_7324,_w_7323,_w_7319,_w_7315,_w_7314,_w_7312,_w_7311,_w_7310,_w_7306,_w_7585,_w_7304,_w_7303,_w_8523,_w_7298,_w_8815,_w_7297,_w_7296,_w_7295,_w_8287,_w_7294,_w_7293,_w_7292,_w_7287,_w_7285,_w_7281,_w_7280,_w_7279,_w_8561,_w_7278,_w_7277,_w_7276,_w_7274,_w_7272,_w_7271,_w_7269,_w_8891,_w_7268,_w_7267,_w_7265,_w_8871,_w_7264,_w_7261,_w_8914,_w_7260,_w_8680,_w_7258,_w_7821,_w_7255,_w_7250,_w_8433,_w_7248,_w_7247,_w_8372,_w_7246,_w_7241,_w_7239,_w_7238,_w_7237,_w_7236,_w_7235,_w_7232,_w_8298,_w_7230,_w_7228,_w_7227,_w_7226,_w_7364,_w_7225,_w_7224,_w_7220,_w_7217,_w_7213,_w_7211,_w_7210,_w_7209,_w_7207,_w_7206,_w_7203,_w_7201,_w_7196,_w_7195,_w_7193,_w_7192,_w_7189,_w_7186,_w_7184,_w_7183,_w_7182,_w_7181,_w_7180,_w_7178,_w_7176,_w_7175,_w_7174,_w_7172,_w_7171,_w_7170,_w_7169,_w_7168,_w_8463,_w_7166,_w_8897,_w_7165,_w_7162,_w_7160,_w_7159,_w_7157,_w_7156,_w_7154,_w_7153,_w_7498,_w_7151,_w_7145,_w_7369,_w_7141,_w_7140,_w_7139,_w_7137,_w_7136,_w_7135,_w_7134,_w_7132,_w_7129,_w_8615,_w_7576,_w_7550,_w_7128,_w_7127,_w_7126,_w_7125,_w_7123,_w_7671,_w_7120,_w_7118,_w_7117,_w_7115,_w_7114,_w_7113,_w_7112,_w_7111,_w_7110,_w_7108,_w_8093,_w_7107,_w_7106,_w_7098,_w_7097,_w_7096,_w_7095,_w_7194,_w_7094,_w_7092,_w_8624,_w_7089,_w_7088,_w_7087,_w_7086,_w_7084,_w_7083,_w_7958,_w_7822,_w_7080,_w_7079,_w_7077,_w_7073,_w_7072,_w_7475,_w_7071,_w_7067,_w_7066,_w_7212,_w_7065,_w_7063,_w_7062,_w_7061,_w_7060,_w_7400,_w_7396,_w_7059,_w_7057,_w_8237,_w_7054,_w_7050,_w_8591,_w_7049,_w_7048,_w_7046,_w_7045,_w_7042,_w_7040,_w_7039,_w_7038,_w_7030,_w_7029,_w_8927,_w_7026,_w_7025,_w_7024,_w_7022,_w_7546,_w_7021,_w_7020,_w_7019,_w_7018,_w_7017,_w_7016,_w_7013,_w_7012,_w_7009,_w_7008,_w_7006,_w_7005,_w_7003,_w_7000,_w_6999,_w_6998,_w_7663,_w_6997,_w_6996,_w_6995,_w_6993,_w_6991,_w_6989,_w_8962,_w_7051,_w_6988,_w_6987,_w_6986,_w_6982,_w_6980,_w_6976,_w_6975,_w_6974,_w_6971,_w_8430,_w_6966,_w_6965,_w_8982,_w_6964,_w_6963,_w_6962,_w_7011,_w_6960,_w_6956,_w_7624,_w_6955,_w_6952,_w_6950,_w_6948,_w_6947,_w_8599,_w_8189,_w_6945,_w_6944,_w_6940,_w_6938,_w_6933,_w_6932,_w_8284,_w_6928,_w_8425,_w_6927,_w_6926,_w_6924,_w_6923,_w_6920,_w_6919,_w_6914,_w_6913,_w_7479,_w_6912,_w_6910,_w_6909,_w_6908,_w_8860,_w_8176,_w_6906,_w_6905,_w_6903,_w_7971,_w_6901,_w_8839,_w_6898,_w_6896,_w_6887,_w_8756,_w_6886,_w_6885,_w_6884,_w_6883,_w_6882,_w_8199,_w_6879,_w_6878,_w_6877,_w_6876,_w_8885,_w_6875,_w_8626,_w_6873,_w_6872,_w_6871,_w_6870,_w_6868,_w_6867,_w_6866,_w_6864,_w_6863,_w_6862,_w_6959,_w_6861,_w_6858,_w_6857,_w_6855,_w_6850,_w_6845,_w_6844,_w_6843,_w_6840,_w_6839,_w_6838,_w_6837,_w_6836,_w_6835,_w_6834,_w_8122,_w_6833,_w_6832,_w_6830,_w_6829,_w_6827,_w_6826,_w_6825,_w_8958,_w_6824,_w_6822,_w_6821,_w_6819,_w_6816,_w_7881,_w_6815,_w_6811,_w_6810,_w_7474,_w_6809,_w_7155,_w_6807,_w_6806,_w_6804,_w_6802,_w_6798,_w_6797,_w_6796,_w_6792,_w_6791,_w_6789,_w_6787,_w_6786,_w_6785,_w_6784,_w_6782,_w_6779,_w_6778,_w_8902,_w_6776,_w_6775,_w_6773,_w_6772,_w_8350,_w_6771,_w_6767,_w_7041,_w_6766,_w_6765,_w_6764,_w_6761,_w_6759,_w_6756,_w_6755,_w_6754,_w_6751,_w_6750,_w_7317,_w_6749,_w_6747,_w_6745,_w_6744,_w_6743,_w_6742,_w_6741,_w_6740,_w_8946,_w_6739,_w_6738,_w_6737,_w_6736,_w_6735,_w_8889,_w_6733,_w_6732,_w_8973,_w_6730,_w_6729,_w_6727,_w_6725,_w_6722,_w_6721,_w_7333,_w_6720,_w_7685,_w_6719,_w_7584,_w_6718,_w_6714,_w_8854,_w_6712,_w_7577,_w_7321,_w_6711,_w_6710,_w_8086,_w_7677,_w_6708,_w_6707,_w_6706,_w_6704,_w_6705,_w_6701,_w_6700,_w_6699,_w_6697,_w_6695,_w_6694,_w_6693,_w_8638,_w_6690,_w_8548,_w_6689,_w_6688,_w_6686,_w_6685,_w_6683,_w_6847,_w_6682,_w_8207,_w_6681,_w_6679,_w_7932,_w_6678,_w_6676,_w_6675,_w_6669,_w_6668,_w_6667,_w_6663,_w_6662,_w_6659,_w_6658,_w_6655,_w_6654,_w_6651,_w_6650,_w_6649,_w_6671,_w_6645,_w_6644,_w_6643,_w_6641,_w_7348,_w_6640,_w_6637,_w_7982,_w_7494,_w_6632,_w_6631,_w_6630,_w_6628,_w_6627,_w_6626,_w_6625,_w_6623,_w_6780,_w_6622,_w_6621,_w_6620,_w_6618,_w_6888,_w_6616,_w_6615,_w_6614,_w_6611,_w_6609,_w_6608,_w_6606,_w_7469,_w_6605,_w_6604,_w_6603,_w_6596,_w_6595,_w_6594,_w_6591,_w_6590,_w_6589,_w_6588,_w_6587,_w_6584,_w_6581,_w_7825,_w_6579,_w_6577,_w_6572,_w_6571,_w_6569,_w_6564,_w_8095,_w_6562,_w_6560,_w_6555,_w_6554,_w_7245,_w_6552,_w_6549,_w_6545,_w_6544,_w_6543,_w_6542,_w_6538,_w_6535,_w_6532,_w_7500,_w_6531,_w_6530,_w_6529,_w_6526,_w_6525,_w_6524,_w_6522,_w_6521,_w_6520,_w_6519,_w_6518,_w_6517,_w_6515,_w_6513,_w_6512,_w_6509,_w_8830,_w_6507,_w_6506,_w_8544,_w_6504,_w_6502,_w_6500,_w_6499,_w_7001,_w_6498,_w_8304,_w_6493,_w_6491,_w_6489,_w_6488,_w_6486,_w_6483,_w_6481,_w_6479,_w_7410,_w_6477,_w_6476,_w_6474,_w_7243,_w_6471,_w_6469,_w_6465,_w_6464,_w_6463,_w_8818,_w_6461,_w_6458,_w_8230,_w_6454,_w_8558,_w_6452,_w_6451,_w_6449,_w_8121,_w_6448,_w_6447,_w_6450,_w_6446,_w_8976,_w_6445,_w_6444,_w_8051,_w_6443,_w_6442,_w_6441,_w_6440,_w_6680,_w_6439,_w_6438,_w_6436,_w_6434,_w_6427,_w_6426,_w_6425,_w_6647,_w_6424,_w_6421,_w_8227,_w_6420,_w_6419,_w_6417,_w_6415,_w_6413,_w_7216,_w_6412,_w_6411,_w_6410,_w_6408,_w_6406,_w_6405,_w_6401,_w_6400,_w_6398,_w_6397,_w_6396,_w_6395,_w_6391,_w_6387,_w_6598,_w_6385,_w_8195,_w_6381,_w_6380,_w_7251,_w_6379,_w_6377,_w_6375,_w_6374,_w_6372,_w_6370,_w_6369,_w_8585,_w_6366,_w_6364,_w_6362,_w_6360,_w_6358,_w_6353,_w_6352,_w_6351,_w_6350,_w_6342,_w_6341,_w_7514,_w_6340,_w_7753,_w_6339,_w_6333,_w_6332,_w_6328,_w_6327,_w_8899,_w_8867,_w_6321,_w_6318,_w_6533,_w_6317,_w_7640,_w_6315,_w_6313,_w_6312,_w_7105,_w_6311,_w_6310,_w_6305,_w_6303,_w_8531,_w_6666,_w_6302,_w_6301,_w_6300,_w_6299,_w_6298,_w_6296,_w_6295,_w_6586,_w_6293,_w_6292,_w_6289,_w_6287,_w_8166,_w_6286,_w_6282,_w_6281,_w_7544,_w_6280,_w_8290,_w_6277,_w_8467,_w_8071,_w_6276,_w_6273,_w_6271,_w_6270,_w_6269,_w_6268,_w_6265,_w_8335,_w_6264,_w_8560,_w_6263,_w_6261,_w_6254,_w_6249,_w_6247,_w_7679,_w_6245,_w_6244,_w_8046,_w_6243,_w_6235,_w_7069,_w_6233,_w_7554,_w_6232,_w_7873,_w_6497,_w_6231,_w_7662,_w_6238,_w_6228,_w_6226,_w_6225,_w_6220,_w_6218,_w_6217,_w_7757,_w_6214,_w_6213,_w_6211,_w_7435,_w_6210,_w_6208,_w_6205,_w_6204,_w_8472,_w_6203,_w_7634,_w_6202,_w_6201,_w_6200,_w_6198,_w_6241,_w_6197,_w_6196,_w_6194,_w_6191,_w_6190,_w_6189,_w_6184,_w_6182,_w_6179,_w_6176,_w_6174,_w_6173,_w_6172,_w_6255,_w_6170,_w_6169,_w_6167,_w_7401,_w_6166,_w_7700,_w_6164,_w_6163,_w_6162,_w_6161,_w_6159,_w_7673,_w_6157,_w_6156,_w_6155,_w_6154,_w_6153,_w_6152,_w_6146,_w_6144,_w_6143,_w_6142,_w_6140,_w_6138,_w_6136,_w_7522,_w_6134,_w_6132,_w_8894,_w_6131,_w_6378,_w_6130,_w_6129,_w_6219,_w_6126,_w_6125,_w_6119,_w_6117,_w_6115,_w_6114,_w_6112,_w_6111,_w_6110,_w_8798,_w_8368,_w_6108,_w_6107,_w_6106,_w_6105,_w_6104,_w_6384,_w_6103,_w_6102,_w_6101,_w_6098,_w_6093,_w_6092,_w_6091,_w_6088,_w_8628,_w_6087,_w_6086,_w_6084,_w_6083,_w_6081,_w_6079,_w_7922,_w_6077,_w_6075,_w_6072,_w_6371,_w_6070,_w_6069,_w_8169,_w_6067,_w_6062,_w_6060,_w_6059,_w_6058,_w_6057,_w_6056,_w_6055,_w_6052,_w_6051,_w_6047,_w_6046,_w_6045,_w_6044,_w_6043,_w_8301,_w_6042,_w_6039,_w_6038,_w_6033,_w_6639,_w_6031,_w_6027,_w_6985,_w_6026,_w_6022,_w_6018,_w_6017,_w_6860,_w_6013,_w_6008,_w_6550,_w_6007,_w_6006,_w_6003,_w_6001,_w_6000,_w_5999,_w_7829,_w_5997,_w_5993,_w_5992,_w_5989,_w_5987,_w_8187,_w_6734,_w_5985,_w_5984,_w_6215,_w_5982,_w_5981,_w_5980,_w_5979,_w_8251,_w_5977,_w_5976,_w_5974,_w_7711,_w_5972,_w_5971,_w_5968,_w_5967,_w_7791,_w_5960,_w_5958,_w_5957,_w_5956,_w_5955,_w_5953,_w_8405,_w_5951,_w_5950,_w_5948,_w_7644,_w_5944,_w_7191,_w_5943,_w_5942,_w_5941,_w_8909,_w_8449,_w_5940,_w_5937,_w_5936,_w_5933,_w_6516,_w_5932,_w_5931,_w_6762,_w_5926,_w_8157,_w_5924,_w_5922,_w_6256,_w_5920,_w_6967,_w_5919,_w_5918,_w_5917,_w_7707,_w_5916,_w_5915,_w_5913,_w_5911,_w_5910,_w_8443,_w_5906,_w_5905,_w_5903,_w_6171,_w_5902,_w_5901,_w_5899,_w_5898,_w_5895,_w_5894,_w_6540,_w_5893,_w_8432,_w_6376,_w_5892,_w_5890,_w_5889,_w_5888,_w_5886,_w_5885,_w_5879,_w_5878,_w_5876,_w_8696,_w_5875,_w_5873,_w_6902,_w_5872,_w_5870,_w_5868,_w_8537,_w_5866,_w_6199,_w_5865,_w_5864,_w_6336,_w_5863,_w_7273,_w_5862,_w_5861,_w_5858,_w_5857,_w_5856,_w_7091,_w_5952,_w_5853,_w_5874,_w_5852,_w_7934,_w_6236,_w_5850,_w_5845,_w_5843,_w_5842,_w_8566,_w_5840,_w_5839,_w_8026,_w_5837,_w_8654,_w_5835,_w_8588,_w_6324,_w_5834,_w_5832,_w_5831,_w_5830,_w_5823,_w_5821,_w_7928,_w_5819,_w_8184,_w_5818,_w_5816,_w_5815,_w_5814,_w_5810,_w_5809,_w_5808,_w_5806,_w_8767,_w_5935,_w_5805,_w_5804,_w_7161,_w_5803,_w_5801,_w_6670,_w_5802,_w_5800,_w_5797,_w_5938,_w_5796,_w_8833,_w_5795,_w_5794,_w_5792,_w_7252,_w_5791,_w_5786,_w_5784,_w_7722,_w_5783,_w_5782,_w_5780,_w_5779,_w_5778,_w_5777,_w_6757,_w_5773,_w_5848,_w_5772,_w_5771,_w_5770,_w_5769,_w_5768,_w_5765,_w_7411,_w_5764,_w_5763,_w_5760,_w_5758,_w_7509,_w_5757,_w_5884,_w_5756,_w_5754,_w_6346,_w_5750,_w_6801,_w_5749,_w_5748,_w_8106,_w_5747,_w_8217,_w_5745,_w_5744,_w_5743,_w_5738,_w_6691,_w_5736,_w_8213,_w_5735,_w_5731,_w_5730,_w_5729,_w_5728,_w_5727,_w_5726,_w_5725,_w_5722,_w_8557,_w_5721,_w_5720,_w_8162,_w_5719,_w_5717,_w_5716,_w_5714,_w_8750,_w_5712,_w_8666,_w_5711,_w_5709,_w_5708,_w_5707,_w_5705,_w_5703,_w_5702,_w_5697,_w_8702,_w_7361,_w_5696,_w_8565,_w_5695,_w_5692,_w_5691,_w_5687,_w_5685,_w_5684,_w_5683,_w_5682,_w_5681,_w_7138,_w_5680,_w_5679,_w_5678,_w_5676,_w_5675,_w_5674,_w_5670,_w_5667,_w_5666,_w_5665,_w_5663,_w_8603,_w_5662,_w_5660,_w_5658,_w_7608,_w_5656,_w_6893,_w_5654,_w_6978,_w_5652,_w_5650,_w_5649,_w_7426,_w_5648,_w_8949,_w_6558,_w_5646,_w_5645,_w_5644,_w_5641,_w_5640,_w_5638,_w_5637,_w_5636,_w_5635,_w_5633,_w_5630,_w_5629,_w_5628,_w_5627,_w_5623,_w_5619,_w_5617,_w_6547,_w_5616,_w_5615,_w_6800,_w_5610,_w_5609,_w_5608,_w_5606,_w_6672,_w_5605,_w_5602,_w_5601,_w_5599,_w_5597,_w_5596,_w_5594,_w_5591,_w_5590,_w_5589,_w_8575,_w_5588,_w_5587,_w_8047,_w_5586,_w_8285,_w_5579,_w_5577,_w_5575,_w_7579,_w_5574,_w_5573,_w_6267,_w_5570,_w_5568,_w_7143,_w_6954,_w_5567,_w_5565,_w_5563,_w_5560,_w_5558,_w_8412,_w_5557,_w_5556,_w_5555,_w_7177,_w_6338,_w_5553,_w_5690,_w_5551,_w_7567,_w_5549,_w_5545,_w_5543,_w_5541,_w_5537,_w_5536,_w_5534,_w_6537,_w_5531,_w_6230,_w_5781,_w_5530,_w_5529,_w_8869,_w_5528,_w_5526,_w_5523,_w_7372,_w_5522,_w_5521,_w_7834,_w_5518,_w_7489,_w_5515,_w_7242,_w_5514,_w_8695,_w_5512,_w_5511,_w_8662,_w_5510,_w_5799,_w_5508,_w_7436,_w_5505,_w_7204,_w_5504,_w_5502,_w_8481,_w_7015,_w_5849,_w_5500,_w_5499,_w_5497,_w_5491,_w_5490,_w_5489,_w_7988,_w_5488,_w_5486,_w_5485,_w_5482,_w_5481,_w_5476,_w_5475,_w_7221,_w_5474,_w_8409,_w_5473,_w_8015,_w_6150,_w_5472,_w_8640,_w_5975,_w_5468,_w_5463,_w_5462,_w_5461,_w_8545,_w_6949,_w_5459,_w_8321,_w_5458,_w_7870,_w_5457,_w_5456,_w_5455,_w_5454,_w_5453,_w_8549,_w_5451,_w_5450,_w_6459,_w_5448,_w_5446,_w_6151,_w_5444,_w_6004,_w_5441,_w_6209,_w_5440,_w_5438,_w_5883,_w_5437,_w_5435,_w_5430,_w_5429,_w_8761,_w_5659,_w_5428,_w_5427,_w_5425,_w_6856,_w_5424,_w_5422,_w_5421,_w_5420,_w_7898,_w_5418,_w_5417,_w_7717,_w_5416,_w_5415,_w_5934,_w_5412,_w_7425,_w_5410,_w_5408,_w_5407,_w_6472,_w_5406,_w_5405,_w_6580,_w_5403,_w_5402,_w_7483,_w_5400,_w_5398,_w_7208,_w_5397,_w_8500,_w_5396,_w_5395,_w_5394,_w_5391,_w_5390,_w_5389,_w_5388,_w_5387,_w_6551,_w_5386,_w_5385,_w_5382,_w_5381,_w_5379,_w_5375,_w_5373,_w_5372,_w_5366,_w_6661,_w_5363,_w_5362,_w_8008,_w_5361,_w_5358,_w_5507,_w_5356,_w_5355,_w_7602,_w_7561,_w_5353,_w_5352,_w_5350,_w_7736,_w_5349,_w_6473,_w_5346,_w_5357,_w_5345,_w_5344,_w_5342,_w_7749,_w_5341,_w_5339,_w_5338,_w_5337,_w_5336,_w_5335,_w_5742,_w_5334,_w_5332,_w_6636,_w_5331,_w_5329,_w_6818,_w_5326,_w_5320,_w_5318,_w_5315,_w_5313,_w_7884,_w_5312,_w_5311,_w_5307,_w_5869,_w_5304,_w_5301,_w_5299,_w_5294,_w_6227,_w_5293,_w_5718,_w_5292,_w_5291,_w_5290,_w_5288,_w_7053,_w_5287,_w_5286,_w_5285,_w_5283,_w_5282,_w_5775,_w_5281,_w_7453,_w_7387,_w_5280,_w_6983,_w_5278,_w_5277,_w_5276,_w_8800,_w_5274,_w_5273,_w_5272,_w_8124,_w_5270,_w_6234,_w_5269,_w_5268,_w_8225,_w_5267,_w_7263,_w_5266,_w_6599,_w_5265,_w_8530,_w_8456,_w_7334,_w_5261,_w_6262,_w_5260,_w_5259,_w_5258,_w_5256,_w_5254,_w_7816,_w_5253,_w_5251,_w_5374,_w_5250,_w_8005,_w_5248,_w_5246,_w_5244,_w_5243,_w_8064,_w_5242,_w_5241,_w_8205,_w_5240,_w_5238,_w_5237,_w_7737,_w_5236,_w_5234,_w_5232,_w_5231,_w_7504,_w_5230,_w_5229,_w_5228,_w_8697,_w_5227,_w_5419,_w_5225,_w_5224,_w_7458,_w_7035,_w_5223,_w_5222,_w_5221,_w_5218,_w_7023,_w_5216,_w_5214,_w_5211,_w_8185,_w_5210,_w_5209,_w_5207,_w_8268,_w_5206,_w_5205,_w_5202,_w_5201,_w_5200,_w_5198,_w_5197,_w_5196,_w_5195,_w_5194,_w_5487,_w_5193,_w_5192,_w_5891,_w_5189,_w_7124,_w_5188,_w_5677,_w_5184,_w_8970,_w_5183,_w_5969,_w_5182,_w_5181,_w_5180,_w_5178,_w_5177,_w_6422,_w_5639,_w_5176,_w_7824,_w_5173,_w_5172,_w_8277,_w_6931,_w_5171,_w_5170,_w_5169,_w_5168,_w_7313,_w_5166,_w_5164,_w_5162,_w_5161,_w_5160,_w_7390,_w_5159,_w_5158,_w_5157,_w_5153,_w_5152,_w_5150,_w_8824,_w_5149,_w_5147,_w_8602,_w_7070,_w_5146,_w_5145,_w_6344,_w_5144,_w_5142,_w_5141,_w_5138,_w_5137,_w_8551,_w_5135,_w_7521,_w_5134,_w_5131,_w_5130,_w_8131,_w_5127,_w_5126,_w_5125,_w_8734,_w_5467,_w_5124,_w_5123,_w_5284,_w_5122,_w_8916,_w_5121,_w_5119,_w_5118,_w_5115,_w_5113,_w_5112,_w_6494,_w_5111,_w_5109,_w_5108,_w_8100,_w_5105,_w_8878,_w_5100,_w_5099,_w_5097,_w_6192,_w_5096,_w_5095,_w_5094,_w_5090,_w_5089,_w_5088,G5250_3,n372_3,G170_3,G170_1,n783_1,n380_2,_w_4776,_w_7916,G177_26,_w_6388,G174_8,n552_1,_w_7254,G177_22,G177_18,G177_13,_w_5962,_w_4568,_w_8085,G177_9,_w_3622,_w_5807,G177_7,G172_10,_w_8501,_w_6768,_w_3611,_w_4578,_w_8960,_w_3745,G128_3,G172_3,_w_4634,G172_2,_w_6503,G172_0,G176_36,G173_27,G173_26,n695_0,_w_6382,n746_1,_w_6874,G173_25,n476,_w_8784,G173_24,G79_1,G173_23,_w_8932,G173_21,G173_20,_w_5600,G173_19,G128_1,_w_8667,_w_5793,G173_17,_w_8657,G117_7,G173_15,G173_13,n187,G173_12,G169_11,_w_6900,G163_14,_w_8332,G173_10,G173_9,_w_3941,G173_6,G173_3,_w_5959,G165_1,n544_0,G173_2,n246_3,n678,_w_5478,_w_3630,_w_7366,G3_1,_w_8780,G3_0,_w_6653,_w_4086,G174_23,_w_3677,_w_3878,_w_7689,G5257_1,_w_7056,G174_16,_w_6258,G174_11,G170_0,n402,_w_5298,G174_7,G174_5,n1013,_w_8203,_w_7863,_w_3602,_w_8248,G175_13,G175_12,_w_6665,n734_1,_w_7680,G175_6,n1222,_w_6239,G175_1,_w_7093,_w_6212,_w_3676,_w_6478,G132_0,_w_6894,n1277,n356_1,n356_0,n1179_1,n552_12,n1179_0,n1263_1,n406_0,_w_4161,G25_1,_w_7036,n1303_2,G168_3,_w_8352,_w_6063,G174_21,_w_4431,_w_5434,G113_2,n804,n400_0,_w_6573,G160_0,_w_8843,n375_3,_w_8407,n825,n375_0,G36_0,n552_2,_w_6897,n630_10,n630_5,_w_3997,_w_7075,_w_5813,n630_0,G86_1,G39_0,G98_19,n479_5,n1058,G171_1,G98_17,n1189,G98_12,_w_4330,n412_0,_w_8411,_w_8180,_w_5175,n307,_w_8757,G98_0,n478_0,_w_4529,G114_0,n655_1,n283,_w_7493,G4_0,G111_2,n722_0,G41_1,_w_5015,G41_0,_w_5321,_w_3619,G2_5,G126_11,G2_4,_w_5496,_w_5235,G172_7,n649,_w_3499,G2_0,_w_4923,G96_5,G96_0,n925,_w_7716,_w_5264,G99_1,_w_5051,n432_1,G174_24,_w_5829,G128_9,G128_8,_w_5376,G177_16,G128_7,_w_4636,_w_5003,_w_5252,G173_22,G5286_5,n346_3,n999,G144_6,G144_5,G6_0,n1074,n596,n630_6,_w_6482,n740_1,_w_4604,G174_18,_w_3679,_w_4810,G128_4,n510,_w_3365,_w_4335,n1443,n665,G139_3,_w_6005,G153_1,_w_5525,n457_0,G61_0,_w_8017,G68_0,n438_3,_w_8436,G163_12,n438_2,G5250_2,n542_1,_w_3460,n438_1,_w_8175,n249_2,_w_4121,n413_3,n697,_w_5576,G123_23,n216,_w_8356,n737_0,_w_8048,_w_4151,G123_19,G123_18,_w_4397,G175_8,_w_4532,G123_1,_w_8749,_w_6224,_w_4968,G70_1,_w_5187,_w_5104,G70_0,_w_5327,n634,n456_6,n465,G79_0,_w_3573,n456_0,_w_6032,n373_0,_w_5887,n409_3,n381_4,_w_5527,n1330,n804_11,_w_4600,_w_3753,_w_4594,n375_5,n381_0,G98_2,G176_19,_w_5061,_w_4557,n1187_0,G119_7,G88_5,_w_8655,n346_0,n326,G92_12,G92_11,_w_7318,n1303_1,n421_1,G92_7,n658,G101_18,G15_1,G92_5,_w_5737,n470,_w_8094,_w_4146,_w_6320,_w_5538,_w_4484,_w_6972,G176_46,_w_8216,G169_13,G169_12,G169_10,G86_0,n443_0,G169_6,n1337_0,G169_4,G175_4,_w_6842,_w_5262,n426_0,_w_3721,G169_3,G90_10,G169_2,G169_0,n537_6,n1280,G113_0,_w_3506,n537_2,n537_0,_w_6684,_w_6541,G5248_2,G5248_1,n1184_0,n1255,_w_3675,n565_1,_w_5480,_w_5371,n394_3,n1449,_w_8441,n249_0,_w_4835,n645_1,n645_0,G172_13,G137_5,_w_8394,n1272_1,G138_4,G175_3,_w_8032,G137_0,n388_1,_w_4162,_w_5143,G14_1,_w_4257,n474_0,_w_6657,n427_2,G80_1,_w_4426,G5243_1,_w_3450,_w_4322,G161_10,_w_6795,n445_1,G2_2,G96_7,G163_6,G138_3,_w_7801,n445_0,_w_3754,n693,G72_1,n587,_w_6180,n1272_0,_w_8937,G173_14,G5251_6,n1285_0,G5251_5,_w_6925,G5251_3,n455,_w_7325,n702,_w_8417,_w_7635,G101_17,G5251_1,_w_7100,G5238_0,G5251_0,n1370,n379_2,_w_4104,n379_0,_w_5880,G5254_3,G88_6,n428_2,G127_0,_w_3668,_w_5219,G149_6,_w_7836,_w_7720,G174_17,G149_5,G149_2,G149_1,_w_5755,_w_4076,_w_5068,_w_7418,G149_0,_w_3929,G5285_5,G5285_1,G5287_3,n469,G123_14,n463_4,G5287_2,_w_4489,_w_8422,G5287_0,n1223_0,_w_7043,_w_3834,G5288_4,n669,G5288_1,n552,n1447_1,G5249_4,G5249_1,_w_5351,n418_2,_w_4487,G5248_4,_w_6435,n379,_w_5668,n264,_w_8035,n1252_1,_w_7560,n804_9,G137_4,n301,n653_2,_w_4115,n653_1,_w_8492,_w_7743,n658_1,_w_7037,n1371_0,_w_8846,n430_1,_w_8067,n1313,_w_4525,G26_0,n409_0,n336,n442_1,n576,_w_5082,_w_4734,_w_8642,_w_6633,_w_5289,n678_1,_w_7007,n1122,_w_6957,n289_1,n588_10,n397_3,n397_1,_w_7055,n1073,_w_7697,n491_0,_w_5930,G5259_3,_w_7775,G5259_2,n780,_w_3620,_w_8429,G140_4,_w_4931,_w_7902,G71_1,G167_3,n758,G176_38,n378_1,n277_0,G5292_2,_w_7253,n243_1,G64_24,_w_8610,_w_8295,G173_7,G128_11,_w_4713,n246_1,_w_6460,n246_0,n637_1,_w_8170,_w_6025,n406_2,_w_5998,G5288_0,n407_1,n408_1,_w_5128,n298_1,_w_6648,G176_27,_w_5384,G2_3,_w_3597,_w_5550,n414_2,n414_1,G174_1,G160_23,_w_5907,G160_14,_w_7488,G113_3,G103_3,G25_0,_w_3695,_w_6799,_w_5877,G160_9,G160_7,_w_7476,_w_6803,G98_13,_w_6487,n1248,_w_3818,G160_5,_w_4934,G160_1,_w_4030,G172_8,G5290_5,_w_5519,n250_0,_w_4820,_w_7443,n630_7,G5249_2,_w_5186,_w_3923,n359,n375_4,G5290_0,_w_8957,G94_13,n884,n424_3,n572_0,n1252_0,_w_4462,n385_2,n318_1,n337,_w_7605,n385_1,n386_3,n394_5,_w_8128,n939,n318_0,n766,G127_1,_w_5954,_w_4016,n387_3,_w_4443,n1428,n643_0,G98_5,n426_3,_w_5136,G172_9,G174_19,_w_8864,n412_2,n704,_w_4475,_w_7967,n643_1,_w_7358,n415_0,G107_10,_w_6951,_w_3858,n1257_0,_w_4720,_w_4085,n435_3,n435_0,_w_7430,_w_6034,G5254_2,n1311_0,n784,n1170_1,_w_7477,G172_14,_w_3951,_w_4767,n1170_0,G177_25,n1184_1,n1125,n1298_1,_w_5604,n770,_w_7149,n409_4,_w_7326,n1298_0,_w_5423,_w_3708,n1214_1,n836,_w_5333,n1214_0,G161_14,n1254_0,n319,_w_3802,_w_4194,_w_6065,n1263_0,n1275_1,G146_3,_w_4365,n372_1,_w_4829,n1275_0,n1282_0,G5292_3,_w_5811,G88_0,n1297_0,_w_3430,n762,_w_6881,_w_6790,n1314_0,_w_8118,_w_7562,_w_4044,_w_6373,_w_6368,n1334_0,G66_5,_w_8480,n1337_1,_w_4658,n268_1,n1359_0,G124_18,_w_4466,n537_1,n698_0,n459,n1374_0,_w_5306,n796,_w_3605,G160_22,n1407_1,n1048,_w_8364,G176_0,_w_8752,_w_6534,n1416_0,n1425_1,n1475,_w_8036,n553,_w_8028,n1450,_w_6021,G124_5,_w_5559,n1425_0,n1431_1,n1431_0,_w_5603,n1440_1,n613,_w_8841,n469_6,n1444_1,G54_0,_w_5065,_w_8172,n479_4,n1447_0,n1394,G98_16,_w_4354,i_G151,_w_3570,_w_4210,n521_0,_w_5516,n1474,_w_8774,_w_7984,_w_4728,_w_5672,n1473,n1289,_w_6122,_w_3558,_w_7167,n1101,n1466,n398_1,_w_7383,n1465,_w_3420,n1464,_w_8733,n1461,_w_3940,n517,n403_2,n1458,_w_6917,n1457,_w_4749,n1456,n1469,n464_5,n1455,_w_6770,n1452,n1448,_w_6480,n1447,n1446,G135_6,G98_14,n1444,n1441,_w_7259,G117_2,n1440,_w_6137,_w_5155,n1439,n1398_0,i_G1,_w_5324,n1435,_w_7405,n1092,n403_1,G137_1,G103_13,n1429,_w_3793,_w_4481,_w_6221,n1427,n1426,_w_4399,_w_4081,_w_4515,n1421,n1420,n1419,n384_0,_w_6123,n347,n427,n1436,_w_5923,n1416,n1422,n1415,n813_0,_w_4135,_w_6322,n1413,G160_20,n1412,n1411,n1407,_w_3447,_w_8309,n1129,G167_13,n1406,_w_4792,_w_6343,n1359,n1237,G159_11,G140_3,_w_4723,_w_5694,n1399,G128_10,_w_4267,n1393,n692_0,_w_7147,n356,G167_5,_w_4480,n1386,_w_3786,_w_5439,G98_18,G123_0,n1383,_w_6082,n805,n639,n1382,G175_9,n1282_1,_w_4827,n574_0,_w_5359,n1374,n256_1,_w_8685,_w_6354,_w_6015,n1325,n1140,_w_5509,n1408,n1369,n1241,_w_3549,n1366,n1362,n1361,n1360,_w_7332,n386,n1352,n769,n1351,G124_7,n1349,_w_7652,n1345,n1341,n1340,n1339,n1234,_w_6511,_w_6290,n521_1,_w_7085,G143_4,_w_4266,_w_8715,_w_8437,n1337,_w_6272,G166_2,_w_6760,_w_3419,n1364,_w_8002,n303,G88_1,_w_6496,n1334,n1063,n1333,n1331,_w_6345,n341,_w_8646,G123_10,n1425,n1328,n1326,n434_0,n1318,_w_4826,n224_1,n1401,G145_1,_w_8489,n513,_w_4991,n1315,G123_17,_w_6096,n537,n1314,G172_12,_w_6899,n448_2,n415_5,_w_3579,n1309,_w_4025,n1305,n1407_0,n1168,n1120,n552_0,n1300,_w_3854,n1135,G102_5,n1362_1,n1297,n1295,_w_7538,_w_4128,n1292,G105_3,n388_2,n473_1,G173_5,n874,_w_7347,n1284,n445_2,n1283,_w_5693,_w_4184,n1282,n1359_1,n380,n1279,n1276,_w_7762,n1275,n1274,n1273,_w_5447,n1387,n407_0,n1271,n1132,_w_8712,G158_3,n1269,n1268,_w_5129,n1267,_w_8665,n1264,n441,n365_1,n1235_0,G84_1,_w_7798,n1270,n1262,n1226_1,n232,n728,_w_4570,n1254,G169_14,n1233,n1253,_w_6617,n603,_w_4851,n731_1,G123_4,_w_8447,n617_0,n1236,n1230,n820,_w_3578,_w_6066,n1226,G160_18,n1223,n1221,_w_6414,n1219,_w_6274,n1218,n1288_1,_w_7519,_w_6113,n1216,_w_6118,_w_3673,_w_5871,_w_4508,n1212,_w_8773,n1211,_w_5970,n1000,_w_6602,_w_4173,_w_5785,_w_4523,n1298,n1012,G139_6,n1210,n300,n1207,n435_4,_w_5449,n1377_1,n352,_w_4295,n1205,n1344,_w_6094,n1342,n1203,_w_5190,n401_1,G69_1,n504,n1208,n1200,_w_5657,n384_2,_w_5767,G126_10,_w_3742,n1199,n374_0,n243_0,n1198,G66_0,_w_4989,n1195,_w_5612,_w_4131,_w_6399,_w_4796,_w_8030,_w_7799,n1193,n1045,_w_4409,n1184,n1300_1,n1305_0,n1183,G175_7,n1182,G92_4,n1180,n1032,_w_4412,_w_4693,_w_7441,n1176,G121_10,n1228,n451_4,_w_6984,_w_5614,G114_1,G96_8,G113_1,_w_7943,n1311_1,_w_3513,n1173,_w_6990,n1170,n1165,_w_7398,_w_3785,_w_4863,n1164,n1162,n421_0,n1176_1,n1161,n1072,_w_4270,G160_21,n394_0,_w_7373,n1158,_w_7779,_w_5929,G23_1,n1157,_w_7417,_w_3455,n392_0,_w_3645,_w_7338,n1155,n409_1,n1153,n881,_w_8063,n1147,n1143,_w_8496,n1139,_w_4041,n1137,n1134,n1133,n268,n1128,n1423,_w_8579,_w_6492,n1126,G128_2,_w_4153,n1124,_w_5432,_w_5431,n1123,n1121,n537_3,_w_4848,n1119,_w_4975,n1301,n1117,_w_5552,_w_4585,n1113,_w_4564,G73_0,_w_4972,n1308,_w_3956,_w_6979,n1110,_w_7623,n665_1,n1105,G5254_0,_w_8194,n1311,_w_7379,n1167,n1103,n1099,n1098,n1430,n1316,n1097,_w_4057,_w_8900,_w_7625,_w_7200,n632_7,n1093,_w_8658,n1087,_w_5073,_w_8981,_w_6074,n1086,_w_8056,n1194,n1107,n1082,G123_8,n655_0,G166_7,n391_3,_w_7741,n804_7,_w_4590,_w_6392,n847,n1078,_w_8408,_w_7363,n964,n1077,n418_3,n433_0,_w_3417,_w_7765,_w_6709,n1346,_w_5365,n552_7,n1186,n1169,n1069,n815_3,_w_4929,_w_3375,n1066,n1064,_w_7491,G160_26,_w_7901,n667_0,G160_19,n1062,_w_8471,n435,G101_11,_w_6036,n1257,_w_8616,n648,_w_7604,n415,_w_5319,_w_6068,n525,G167_11,G111_1,_w_8568,_w_5572,G177_5,G160_3,G158_0,_w_3629,_w_4748,n1211_1,_w_6716,n1391,_w_3529,_w_4730,_w_6635,n494_1,_w_8630,_w_6308,G27_0,n652,_w_4384,_w_8944,n268_0,_w_3788,n426,n608,_w_4542,G158_16,_w_4378,_w_7670,n505,_w_4250,_w_4179,G24_0,_w_7354,n877,G148_6,n1213,_w_3503,n802_8,n318,n376,n1252,n1324_0,_w_6805,G174_14,_w_8344,n751,n1247_1,_w_4430,G5221_5,_w_4963,_w_8724,_w_5226,n1347,_w_3853,n986,n1395_1,n378_0,n632_5,_w_8954,n363,n434,_w_6777,_w_4948,_w_7368,_w_4062,_w_5927,n207,_w_8039,G90_13,_w_3463,n424,_w_5392,G172_11,_w_8912,n1268_1,_w_7734,n350,_w_5443,n413_0,n343,n653_0,G132_1,G176_52,n606,n425_1,G64_21,n335,_w_3617,_w_7010,n1308_0,n573,_w_4706,_w_8880,n799,G5242_1,n1384,_w_8895,n872,_w_8917,n1266,n1198_0,n526,_w_8103,_w_7322,n773_5,n323,_w_5117,n643,_w_5904,_w_4285,_w_4416,n322,_w_5404,n416,n357,n962,n802_7,_w_7496,n783,n1172,G5255_1,_w_5413,n320,_w_4836,_w_7597,G173_4,_w_7284,n417,n315,n1477,n401,n1192_1,_w_5774,n311,G150_2,_w_3528,n379_3,_w_7559,n491_1,n1227,_w_4819,n854,_w_6175,n1090,_w_5053,n857,n279,_w_5580,n1146,_w_6922,_w_4681,_w_8336,n1444_0,_w_4661,n297,n414,n298,G159_0,_w_4752,n523,_w_4216,_w_4000,n1096,n384_3,G92_3,n1037,G155_0,n951,G145_6,n287,n952,_w_6510,_w_4653,G96_12,_w_8379,n931,n302,_w_6109,_w_4026,G92_2,_w_7214,G14_0,G5245_0,_w_8083,n469_10,_w_6097,n278,n583,_w_8061,G150_5,G174_10,G96_2,n276,_w_4071,_w_4265,n407,n418,n943,n307_0,_w_6148,n208,_w_6020,n524_0,n273,_w_7283,n1053,_w_4965,_w_6029,_w_3864,_w_7547,n313,_w_6054,G173_1,n272,_w_5328,n711,_w_5087,n442_0,_w_3640,n267,_w_7614,n1338,_w_5535,n479,_w_3988,n856,_w_6071,G5243_0,G121_6,_w_6889,n1357,n1374_1,n258,n374,_w_7841,G142_3,_w_6361,_w_3698,G172_5,n255,_w_7970,_w_7854,G115_5,_w_5110,n252,_w_6237,n876,_w_8042,_w_6895,n863,_w_6961,G175_10,_w_5582,n924,n246,_w_8186,_w_7587,n463,_w_6490,n714,n378,_w_3795,_w_4113,G5248_0,_w_6485,n238,_w_7842,_w_4247,_w_7455,n1005,n243,_w_7745,n241,G88_3,n574_1,_w_8779,_w_8759,_w_7391,G5221_7,n289,G5292_1,G107_13,n239,n646,G177_6,n342,_w_7794,n477_1,n230,n229,G146_1,_w_5347,n1028,_w_6116,n228,_w_8710,n691,G177_0,_w_4145,n224,_w_5826,n1336,n450,n469_4,n651,_w_4372,_w_6553,_w_4640,n868,n865,_w_8326,n1251,_w_5539,_w_3659,_w_7492,n277_1,n214,_w_8043,_w_7532,n1322,_w_6257,G5249_5,n213,_w_6646,n1254_1,_w_4638,n1403,n211,G144_4,n221,_w_6095,_w_5084,_w_7724,_w_6329,n432,_w_5057,_w_5029,n430,G24_1,_w_3383,n1386_1,n392_1,n415_4,n1385,G5213_1,_w_3406,n1175,n193,n435_1,G123_11,_w_5383,n201,n412_3,n188,n266,_w_3946,_w_8980,_w_8241,_w_5249,_w_4902,_w_7668,n779_0,n887,_w_3515,_w_6828,_w_5049,n1398,n1260,n189,n406_3,G158_25,n1176_0,_w_8669,_w_5028,_w_4957,_w_8114,n815_10,_w_6612,n292,n521,_w_6278,n698,_w_8444,_w_5825,G174_3,_w_6078,G5288_3,n896,_w_3741,n403,_w_8898,_w_5554,n719_1,n1396,n1138,n1232,n752_0,n968,n802_3,n251,G162_0,n394_4,n196,G174_22,_w_6085,n1445,_w_4880,n377,_w_3875,_w_8360,G100_0,G145_4,_w_8614,_w_4998,n1365,_w_8450,n257,n349,n420_0,n500,_w_7058,_w_6943,_w_5414,n419_1,n632_6,_w_7300,G36_1,n222,_w_3886,_w_5963,_w_5380,_w_7923,n1332,_w_8775,_w_8716,_w_5626,_w_4122,n373_1,_w_4261,n442_2,G176_37,G177_24,n324,n614,_w_3958,_w_8146,G173_16,G177_15,n593,n766_1,_w_6035,G124_13,G5287_1,G18_0,n1018,_w_4123,_w_7713,n1323,_w_7231,_w_6283,n381_3,_w_3777,_w_6359,_w_4005,_w_7440,n463_3,G131_1,G128_0,n1467,n428,n405,_w_3393,n437,_w_8098,n1256,_w_7785,n1288,n1390,_w_3942,_w_5965,G123_12,n1141,n703,_w_5010,_w_5540,_w_4830,n664,n1148,_w_4895,_w_8366,G113_5,_w_4334,n1201_1,n1354,_w_4655,n1204,n773_6,n803,_w_7937,n445,n325,n1392,n670,n277,_w_8439,n637,G169_8,G96_3,_w_3680,_w_8000,G5254_1,_w_6812,_w_6127,G77_1,n667,n572_1,n1268_2,_w_5479,n404,_w_7299,G27_1,n588_2,n1244_0,_w_4028,n759,G94_2,G176_44,n361,n493,n945,_w_6723,n394,_w_6099,n642,G128_12,_w_4199,n1247,G142_1,_w_4857,n284,n612,n223,G98_3,_w_4220,n386_6,_w_7233,_w_4205,n565,n344,_w_6316,n364,_w_6970,n274,G158_2,G87_0,n1022,n294,G5285_0,_w_6808,n624,_w_4386,n392,G5260_5,n1377,_w_8145,n450_0,_w_3928,n917,n1379,_w_6953,G5287_4,_w_5973,_w_5016,_w_6852,n670_1,_w_3844,n853,_w_5445,_w_4353,_w_5257,G158_21,_w_4649,n1150,n930,n766_0,_w_8747,_w_7879,_w_7270,n494,n398_0,n254,n647,_w_5040,n695,G5260_3,_w_6934,_w_4764,_w_4888,_w_5023,_w_7790,_w_4526,G175_14,_w_4925,n263,_w_4171,_w_8984,G21_1,_w_7875,_w_4418,G126_8,n1211_0,n384_1,G123_20,n385_0,n707_0,_w_7014,_w_7101,_w_4479,_w_8678,G169_1,_w_8073,n312,n442,_w_5762,n998,n717,n1358,G77_0,G176_32,n328,_w_7355,_w_5348,n1160,n435_2,_w_5302,_w_4022,n330,_w_4700,_w_8434,n1187,_w_6323,n429,_w_3574,n1373,n824,n381,G5262_1,n514,G177_29,_w_6918,_w_6306,_w_5881,n686,_w_8416,n452,_w_6597,n227,G124_17,_w_7903,n802_0,n373,_w_6696,n502,G64_9,n456,n1306,n922,n802_10,n436,_w_7116,_w_4042,_w_5996,n334,_w_8540,n588_6,n1389,_w_8807,_w_6660,_w_5101,n339,G160_16,n413,G5290_3,_w_3790,_w_4349,n249,n321,n234,_w_5945,n438,_w_6484,_w_4853,_w_4970,G169_7,n1414,_w_8148,n1094,G81_1,G177_12,n556,G105_13,_w_7102,_w_4031,n378_2,G176_42,_w_8847,n259,n365_0,n224_2,_w_4038,n384,n1039,n1214,n1004,_w_7609,G174_26,_w_5986,n914,n1020,n395,n557,_w_8819,n632_4,n1195_0,n500_0,n556_1,n479_1,_w_3966,_w_4307,n240,_w_7523,n699,G5293_0,_w_7676,n630_9,_w_7610,G150_1,n403_0,_w_3413,_w_7222,_w_5584,_w_3738,n666,n218,G156_1,_w_8593,n365,_w_3688,_w_5079,_w_8722,_w_7307,_w_6061,n393_0,n346,_w_7991,n840,_w_6619,n1355,n366,_w_4290,_w_5494,_w_4800,n206,_w_6141,n399_0,_w_4050,_w_7198,G144_0,G100_15,n1272,n333,_w_5533,n903,_w_7078,G121_7,_w_5203,n386_2,_w_8513,_w_3774,_w_4240,_w_4245,n597_1,_w_4421,n1285,n1235_1,G5288_2,n830,n1334_1,n389,_w_7104,n332,n434_2,G175_0,_w_8608,_w_6325,G96_1,_w_7702,n686_1,n249_1,_w_8060,_w_5014,_w_4786,_w_8081,_w_4326,n400_5,n452_0,n655,_w_8215,n391,_w_7413,_w_3481,_w_7940,_w_6846,_w_5133,n1329,_w_3484,G83_1,_w_5377,n1317,_w_3382,n630,_w_3881,_w_4163,n419,G76_0,n684,n607_0,_w_4292,n375,G161_3,_w_5949,n692,G174_9,_w_3595,_w_7229,G5292_4,_w_4612,G158_12,n745,_w_4287,G160_17,n552_15,n834,n400,n950,G94_4,n1303,_w_8987,_w_7921,n314,G158_1,n1159,n601,_w_6363,n588,G5260_1,_w_3418,_w_8840,_w_7626,_w_5964,n767,n1453,n813_9,_w_7187,n707_1,_w_4391,_w_4319,_w_5116,n469_9,n1444_3,n379_1,n760,_w_6030,_w_3932,n546_1,_w_8975,_w_3792,_w_5034,n372_0,n1432,n519,n429_1,_w_5484,n1179,n281,n773,_w_3991,_w_7714,_w_5426,n456_2,_w_8476,G107_0,_w_3976,G123_22,n1191,_w_8142,G130_1,_w_4565,_w_8832,_w_6814,n354,_w_5370,n1307,n217,n1108,_w_7888,_w_6758,G143_1,_w_6794,_w_5309,_w_8337,_w_7738,n552_19,n740_0,n421_5,_w_4414,_w_5710,n492,n1332_1,n1055,_w_7527,_w_4268,_w_8731,n631,n592,n1363,_w_3387,n1061,n869,_w_3491,n508,_w_8582,_w_5367,G177_10,_w_7142,n413_1,n290,_w_8570,G81_0,_w_3678,_w_4813,_w_8959,n1085,_w_3378,_w_8576,_w_3986,G5290_1,_w_3479,n372,_w_7033,n630_4,_w_4662,_w_6120,n1235,_w_5156,_w_3807,_w_3931,_w_4187,n394_1,_w_5369,_w_4277,_w_5715,_w_5566,n1223_1,n744_2,n622,_w_8821,_w_4099,_w_4769,n661,n1204_0,_w_3749,_w_7466,n726,_w_4964,n286,_w_6347,n967,n755,_w_7540,_w_3971,_w_5013,n288,_w_8428,G124_0,_w_5909,n729,G5258_2,_w_8673,n414_0,n746,G5253_3,_w_6089,G177_1,n425_2,_w_3935,n1424,_w_7907,n970,_w_6009,_w_3718,n544,_w_8365,n993,_w_8319,n1250,_w_4259,_w_3510,n776,_w_8705,G5291_5,n678_0,_w_7482,_w_7244,n224_0,n563,n1111,_w_8539,_w_8136,n994,n225,n309,_w_3797,_w_7658,_w_6642,G149_4,_w_3731,_w_3643,_w_6582,G175_5,_w_5634,G159_12,_w_6158,G166_1,_w_5139,_w_7866,_w_7144,G107_3,_w_6916,_w_5163,n1112,_w_3817,n723,_w_3884,_w_8182,G69_0,_w_3706,n512,_w_6475,_w_4742,n1292_1,_w_7031,_w_4007,_w_4930,n497_1,n1166,_w_3707,_w_8012,G5250_0,_w_6958,n1024,G137_3,_w_8494,_w_4348,G5249_3,_w_3930,_w_7179,_w_4778,_w_4874,n399_1,_w_6793,n296,G100_1,_w_5624,_w_3964,_w_6593,n793,G169_5,_w_4312,_w_8150,n1303_0,_w_3663,n811,n1400,_w_3921,n531,n849,_w_7721,_w_6527,n1190,_w_3729,_w_7223,_w_5012,_w_5761,_w_4719,n1447_3,G5244_0,G121_11,_w_7843,n202,n1174,n598,_w_6266,n520,n933,_w_7219,_w_4854,n397_2,n1206,_w_8933,_w_3959,_w_6402,n1263,n497,n798,_w_7190,n398,n958,G160_10,n1226_0,_w_5075,n463_2,_w_7345,G98_6,n1372,n360,n415_1,G124_1,_w_8077,G5285_4,_w_5561,n1451,G5288_5,n1428_1,n716_1,n1310,n750,n983,n265,_w_8168,n421,_w_4553,_w_6831,_w_6145,n671,_w_5024,n391_1,G68_1,_w_3625,_w_3505,_w_4877,n372_2,_w_5470,n632_0,n532,n1290,n191,_w_6355,_w_3412,n785,_w_6656,n1247_0,_w_5547,G135_4,G5242_0,_w_3523,n233,_w_5578,_w_5007,_w_3638,_w_7858,_w_4966,_w_8892,_w_6557,n828,n810,n1149,n260,_w_4917,n1240,_w_8519,n367,G153_0,G98_8,n761,_w_8363,n443_1,G5253_4,_w_5074,n860,_w_6698,n348,G177_19,_w_5542,n305,n527,n1417,n637_0,_w_4624,G5260_4,_w_5035,_w_5812,G137_6,n1089,n295,n706,n870,n915,G130_3,_w_4982,n423,_w_7340,G100_3,n545_3,_w_3820,_w_7320,n1405,_w_5296,n375_2,_w_8683,_w_5713,_w_4206,_w_5154,G5285_2,G126_4,n1320_1,_w_7636,_w_5820,_w_8370,_w_6393,n590,_w_7705,_w_5595,n995,n736,n694,_w_3568,n406_1,_w_4125,G135_2,n1204_1,n1296,_w_3692,n253,G54_1,n963,n898,n539,G102_1,_w_3496,_w_3805,_w_7433,n744,G168_9,_w_4406,n1472,n1317_1,_w_4664,_w_7755,_w_8555,_w_8123,n842,G105_11,n465_0,G169_9,_w_8778,_w_7553,_w_5741,n439,_w_4906,n440,n291,n355,n749,n838,n289_0,_w_7412,_w_6848,G141_4,n1243,n638,n443,_w_7262,_w_5368,n1299,_w_8278,n269,n1114,n1368,n448,n555,n282,n446,_w_5492,G175_11,n447,n1312,_w_3733,n1356,_w_7185,G109_7,_w_4325,n451,_w_7740,G119_1,_w_4522,_w_4097,n716,n244,n453,_w_8825,n556_0,n681,_w_4652,n362,n454,n1258,_w_3697,_w_6222,G160_6,n879,_w_4080,n457,_w_4023,_w_5700,G132_2,n668,_w_4182,G92_9,n458,G174_6,n242,n674,_w_6854,n760_1,_w_5140,n1057,G113_6,n894,_w_5838,n461,_w_7763,n1071,n548,G176_6,G5290_4,_w_7291,n1377_0,n522,_w_4616,n467,_w_8027,_w_6437,n689,G1_1,n908,_w_6774,_w_4137,n329,_w_7558,n609,n433_2,n471,n794,_w_5064,n472,n878,n516,_w_5483,n942,_w_7234,_w_7511,n511,n474,n1350_0,_w_6050,_w_5107,G98_9,n1319,_w_5501,n464,n1196,n1434,n837,n475,n480,_w_3511,n481,_w_5620,G161_8,_w_4758,n426_2,_w_7708,_w_5860,n483,G18_1,n375_1,_w_6731,G166_9,G5253_1,_w_3879,n484,_w_4117,G98_4,G92_6,_w_4714,n485,n1409,G121_2,n358,_w_7367,_w_3458,n478,n594,_w_4832,n400_1,_w_6076,_w_5671,n552_6,n487,n449_0,_w_7811,_w_3796,n370,n489,_w_8704,n403_3,n490,n1054,_w_8050,G96_6,n1156,n310,n491,n298_0,_w_7595,n498,_w_7571,n237,n388_0,n426_1,n499,n501,G161_2,_w_3943,_w_4815,n503,_w_3799,_w_5625,n641,_w_4939,G5286_3,n209,n507,n535,n515,n777,_w_8288,_w_6470,_w_4429,n923,n1220,_w_8674,_w_8574,_w_5698,G101_0,_w_4839,_w_5360,n409_5,G5213_0,_w_7815,_w_4535,_w_6251,n428_1,n1371_1,G5199_1,_w_8645,_w_5966,G167_7,_w_3624,_w_7868,n848,G160_4,n686_0,n524,_w_8240,_w_5330,G161_4,n381_5,n530,n732,n1038,n534,n1302,n786_1,G121_8,n408,n381_2,n540,n368,G174_27,n541,_w_7899,n708,_w_4346,n415_3,G166_13,n629,n547,n549,G158_10,n818,n459_0,G177_8,G168_4,n1268_0,_w_4688,n559,n438_0,n560,_w_3666,_w_7044,_w_6508,n1343,G160_12,_w_7286,n567,n256,n957,n744_5,_w_4464,n306,_w_8459,n562,_w_5030,n1106,n571,G5248_3,_w_3672,G160_11,n1238,n1115,n944,_w_7826,_w_5041,n537_4,G177_2,_w_6539,_w_5882,G140_2,_w_7257,G5291_4,_w_4309,n660,G103_2,_w_5631,n1289_0,_w_8746,G176_10,n1151,n575,_w_3606,_w_7796,n580,n735,_w_8390,_w_7081,n584,_w_6259,_w_4356,n1079,n1246,_w_5751,n626,_w_5055,G177_20,n940,_w_3798,n1044,n1281,_w_8440,G100_20,_w_6090,n585,_w_3536,G5248_5,n542,n424_2,G126_5,n1014,_w_7849,G177_23,n1041,_w_3850,_w_6935,n727,n960,_w_4699,n589,_w_4799,n595,_w_6389,n1459,_w_8598,_w_4177,n597,_w_4866,_w_6505,n212,_w_7486,n599,_w_7930,G174_0,n1008,n600,_w_8292,_w_3544,G21_0,n1046,_w_8785,n722_1,n632,n1195_1,n602,_w_5643,n1084,n1288_0,n1030,_w_6284,n204,n701_0,n607,n700,n432_0,n1297_1,n1202,_w_4574,n610,n815_11,G123_13,n616,G42_1,_w_7309,n617,_w_4588,n619,n424_1,_w_7481,_w_4953,n621,n1250_1,n779,n623,G149_3,n800,_w_4677,_w_5753,_w_5611,G160_25,n327,G98_15,n959_1,n628,n636,n1016,G176_8,_w_4785,_w_6674,_w_5928,n427_1,n640,n1065,_w_3762,n419_0,n399,n791,n542_0,n219,n1317_0,n444,n935,n656,_w_7592,_w_4609,n662,G5286_1,n415_2,n890,_w_4350,n1178,n712,_w_8714,_w_4201,_w_3650,n380_1,n1060,n672,G92_1,n673,_w_5673,_w_3962,G96_11,n862,n765,G40_0,_w_4120,_w_5080,_w_6462,n1209,n676,_w_3400,n586_11,_w_8583,n677,_w_8384,_w_3768,_w_8144,n695_1,_w_4223,_w_5004,_w_4843,n679,n680,n402_1,_w_4881,_w_5300,_w_3642,_w_4238,n488,n682,_w_7002,n826,_w_8908,n913,_w_3980,_w_3725,G144_2,n690,G17_1,G6_1,_w_7744,_w_6335,_w_6048,n701,n410,n705,_w_6570,_w_3865,n738,_w_6941,_w_4339,n391_2,_w_8532,n845,n715,_w_6813,G94_1,n1479,_w_7122,G16_0,_w_7301,n719,G123_2,_w_5789,n316,_w_5247,n813_10,n720,G98_11,_w_4147,_w_6702,_w_4320,n1224,_w_7275,n721,G39_1,n748,n1468,n1292_0,n731,_w_4239,_w_8197,G144_3,n381_1,G147_0,n734,n737,n786,n477,_w_6428,_w_5085,n778,n742,G160_24,_w_8931,n768,n1070,n463_5,G72_0,n1088,_w_7672,n753,G177_27,_w_4817,_w_6566,n754,G92_13,_w_5817,n966,n1348,n1229,n1010,n757,G5287_5,_w_3434,n1164_1,n1201,n904,_w_5571,_w_4438,n973,n891,n772,n787,_w_5308,n248,_w_4552,n409_2,n552_14,n383,_w_8355,n953,_w_3646,_w_8404,n1378,_w_4497,n873,_w_6386,G88_4,n812,_w_8462,G176_12,n817,n781,G5249_0,n722,n408_0,G5257_5,n788,G96_10,_w_5990,n1460,_w_4824,_w_4745,n789,n1042,n790,_w_4056,_w_4021,n1017,_w_3833,n433_1,n792,n1287,n488_1,_w_5827,n1177,_w_6859,_w_4805,n424_0,n378_3,_w_5867,n515_1,_w_5279,n1116,G100_13,_w_4900,n801,_w_6365,n802,_w_3832,_w_4269,_w_5613,n948,_w_6149,n807,_w_4083,G74_1,_w_4357,n420_1,n809,_w_5532,n769_1,n956,n813,_w_8534,_w_7442,G23_0,_w_5393,n888,_w_6781,G107_1,G109_4,_w_7933,n815,G73_1,n1244,_w_4260,n473,n816,n387_0,n716_0,G88_7,n1040,n821,_w_7594,n981,_w_3950,n422,_w_3488,n823,G168_11,n829,_w_6892,_w_5409,_w_4422,n839,G5259_0,G135_0,G167_9,n844,_w_4884,_w_4440,n696,n588_3,n846,G5221_9,_w_3767,n850,n1285_1,n880,G64_18,n882,n463_1,_w_5854,_w_4980,n889,_w_5978,G103_0,_w_4018,_w_4141,_w_5378,G177_4,n402_0,n1225,_w_4538,n893,G166_10,_w_6936,n895,_w_5787,_w_5471,n897,n1049,n558,n905,G5257_2,n307_1,n380_0,n907,_w_8562,_w_7914,_w_5132,_w_4444,_w_4907,_w_6357,_w_4977,n1304,n909,_w_7993,G17_0,n927,G90_12,_w_4899,n916,_w_7835,n822,G158_23,_w_3489,n430_0,_w_4891,_w_7686,G163_1,n220,G5286_4,_w_4231,G22_1,n926,_w_4949,_w_8808,n578,_w_4419,n692_1,n654,n804_2,n929,_w_4850,_w_8796,_w_7603,G2_1,n1080,_w_4448,n932,G5285_3,_w_8104,n630_3,_w_3894,_w_6023,n375_6,n413_2,n934,G128_13,G123_21,n1231,n813_1,n941,_w_6195,_w_5036,n947,n782,_w_4575,n959,n1197,n961,n1031,_w_7996,n418_1,n965,n449,n815_8,G98_1,n971,G123_16,n833,_w_7622,_w_3509,_w_7983,n1478,n744_1,G5258_4,_w_8006,_w_7812,n1291,n976,_w_4078,_w_8802,G176_17,G105_0,n980,_w_4610,_w_8820,_w_7852,n1362_0,n985,_w_6423,G5293_3,_w_3804,n250_1,n987,_w_5297,n756,n451_3,G174_25,n574,_w_3588,n989,_w_6841,_w_3540,_w_3770,_w_8791,n921,n740,_w_4176,_w_8670,G123_15,n804_4,G139_2,n1192,_w_4852,G121_0,n815_4,G84_0,n724,n1026,_w_6783,n1002,n763,n1025,n1006,n586_1,_w_8915,_w_7615,_w_5651,_w_4014,n1007,_w_4994,G173_8,n795,n912,_w_4317,n1011,G5251_4,n317,n1047,n1023,G74_0,G98_7,n246_2,_w_8151,_w_4215,n1029,G143_6,_w_6556,_w_5607,_w_5498,_w_4892,n1034,n451_2,_w_8587,n528,G160_27,G5_1,G101_1,n1164_0,_w_4066,n1402,n1050,G5254_4,_w_5469,n1404,n1052,_w_6652,n959_2,_w_8934,n1056,n1286,G5250_4,_w_8698,G5250_5,_w_4241,_w_6100,G167_0,_w_7862,_w_4571,_w_8369,G167_1,_w_5790,n586_10,G92_10,G167_2,G167_4,G167_6,_w_5701,_w_3911,G5259_4,G167_8,n899,_w_3377,n975,G167_12,_w_3960,_w_6307,G166_3,_w_8183,n547_0,G166_4,G166_5,G166_6,_w_7389,n1036,G166_8,n435_5,_w_4124,G166_11,G166_12,G119_3,G166_14,_w_6677,G80_0,G165_0,_w_7938,_w_5664,G147_6,n813_3,n538,G117_0,G117_3,G117_4,_w_3861,G117_5,G117_6,n988,_w_4958,G5257_0,G5257_3,G5257_4,n746_0,_w_5517,n425_0,n425_3,G147_4,G168_12,n546_0,n456_4,_w_3810,_w_5464,_w_3600,n1245,n544_1,_w_3913,_w_4646,_w_8474,_w_3696,G146_0,_w_5303,G146_2,_w_7649,n1395_0,_w_8299,_w_7524,G156_0,n776_0,_w_8911,_w_7004,G161_0,G161_1,_w_5855,_w_3623,G161_7,_w_4401,_w_5018,_w_5524,G161_9,_w_6367,G161_11,_w_3869,G161_12,_w_3667,G161_13,G158_4,_w_5005,G158_5,_w_3372,_w_4582,G158_7,n468,G158_8,_w_6016,G177_21,G158_9,_w_5047,G158_11,_w_5506,_w_4889,G158_13,_w_4342,G158_14,G158_17,G61_1,G155_1,_w_7382,_w_6139,_w_5411,G158_19,G158_20,_w_8003,G158_22,_w_3398,_w_7778,G107_2,_w_3456,_w_6457,G107_4,G107_5,G94_6,_w_6468,G107_6,_w_4580,G107_8,G107_9,G107_11,_w_8652,G5291_0,G5291_1,G176_23,_w_4160,n253_0,_w_4809,G5291_2,G176_50,_w_5546,n747,G5291_3,_w_8693,_w_3664,_w_6565,n954,G5221_0,_w_7581,n1476,_w_3814,G5221_1,G5221_2,_w_3684,G5221_3,_w_4912,G5221_4,G103_8,_w_5988,_w_3938,n1249,G5221_6,G5221_8,_w_7664,_w_6523,_w_5732,_w_3555,_w_3583,G85_0,_w_7215,_w_7150,_w_5503,_w_4486,G85_1,n804_1,G158_24,G159_2,G159_3,_w_7994,G66_1,G159_4,n400_2,n773_1,_w_6433,_w_5585,_w_5493,G168_0,G159_7,n1434_0,G102_0,_w_8682,n666_0,_w_5323,G159_9,G141_1,n331,G159_13,_w_8044,_w_6177,G159_14,G152_0,_w_6610,_w_4648,_w_4059,G150_0,G150_3,_w_6820,G82_1,n741,G150_6,_w_4333,_w_4060,n512_0,n512_1,G160_8,n607_2,n704_0,n704_1,_w_6331,G148_0,n1033,G102_2,G148_2,_w_6431,_w_3874,G148_3,_w_7742,n1259,G148_4,_w_7927,_w_6019,G145_0,G145_2,G145_3,G145_5,n936,G163_0,_w_7282,G163_4,_w_6664,G163_5,_w_4455,G163_7,_w_6288,G163_8,G163_10,G163_11,G173_18,G124_14,_w_3952,_w_8490,G143_0,G143_3,G143_5,G87_1,G141_0,G141_2,G141_3,_w_5174,G141_5,_w_3885,G117_1,G141_6,G130_2,n773_3,G130_4,_w_7173,_w_4765,n1332_0,_w_7188,n476_1,_w_4381,G138_0,n1418,n552_5,G138_1,_w_8495,_w_4735,_w_7349,G138_5,G94_0,n1433,_w_4395,G138_6,_w_3371,_w_8209,G143_2,_w_3560,G135_1,G135_3,_w_3628,_w_6728,G135_5,G64_22,n632_1,n552_3,_w_6080,_w_3593,n552_4,n552_8,n552_10,G124_12,_w_4053,n552_11,n552_13,_w_7472,_w_6578,_w_3896,G124_19,n552_17,_w_7809,_w_7133,_w_3766,_w_3473,n552_18,n552_20,n552_9,n552_21,_w_4583,_w_4595,n552_22,_w_4940,n552_24,_w_7660,n769_0,_w_4380,n497_0,G101_8,G168_1,G168_2,_w_4347,G168_5,_w_7926,G168_6,G168_8,_w_8811,G168_13,_w_5322,G26_1,_w_7290,_w_3715,_w_4108,_w_6865,n402_2,n543,_w_3615,G126_0,_w_7805,G126_2,_w_6466,G126_3,_w_6285,_w_3880,n620,G126_6,_w_3392,G126_7,G126_12,G126_13,G64_11,_w_6638,G92_8,_w_4193,_w_4306,n421_3,n421_4,n386_5,G125_0,_w_6187,G140_5,G125_2,_w_8202,_w_8068,n387_1,n630_1,G167_10,G157_0,G157_1,G157_3,G131_0,G140_6,n632_2,n632_3,_w_8723,n630_8,_w_4367,n632_9,n632_10,_w_6432,_w_3653,_w_8322,n1187_1,G105_7,n632_11,n472_4,_w_4771,G124_3,_w_8729,_w_7569,_w_5851,n813_7,G124_4,_w_8754,G101_7,G171_0,G124_8,G124_9,_w_7427,_w_6880,G124_10,G124_11,_w_8330,G173_0,n813_2,G124_15,n775,G150_4,G124_20,G124_21,G124_22,G124_23,_w_7356,_w_5946,G124_24,_w_8812,_w_4736,G124_25,_w_7797,_w_4211,n299,n1388,G121_1,_w_5091,n730,G121_3,_w_4355,G121_4,_w_8939,G121_5,G121_9,_w_7770,G121_12,G121_13,n233_0,n233_1,_w_4606,G16_1,n233_2,_w_7601,_w_4601,G5239_0,_w_6133,G100_9,_w_8795,_w_8677,G78_0,_w_8137,_w_5739,_w_5148,n1353,G4_1,G159_10,G78_1,G119_0,_w_5069,_w_4114,G119_2,G119_4,_w_7645,_w_4236,G119_5,n256_0,G119_6,n1278,_w_3893,_w_7637,n1192_0,_w_5746,n1416_1,G11_0,_w_7448,G11_1,G109_0,n382,_w_4566,G109_1,n399_2,G100_5,_w_8221,_w_6673,G109_2,_w_8753,_w_3871,G109_3,n779_1,_w_5569,G109_5,G109_6,G109_8,G109_10,G99_0,_w_4680,G5292_0,G109_12,_w_8904,G109_13,_w_5618,n1201_0,G105_1,n1444_2,G105_2,G105_10,n409,G105_6,_w_8306,G105_8,G5290_2,_w_4478,n866,G105_9,G105_12,G101_4,G5286_0,_w_6501,_w_3391,G5286_2,_w_5093,G140_0,_w_7249,_w_3542,_w_8509,n463_0,G140_1,n406,G129_0,_w_8024,_w_5562,n644,_w_4200,G103_4,_w_8760,_w_3530,_w_6583,G103_5,G103_6,_w_6216,G103_7,_w_7099,n776_1,G103_9,_w_7341,n1437,G103_10,_w_6429,_w_3780,G103_11,_w_8755,G101_2,_w_8842,_w_7454,_w_3702,G101_3,_w_8141,n1257_1,G101_9,_w_8554,n464_3,G101_12,G101_15,_w_8919,_w_5598,G101_16,_w_7617,G101_6,_w_4794,_w_7308,n462,G101_19,n804_8,G100_2,G100_4,_w_6763,G92_0,n710_0,_w_6073,_w_3427,G100_7,_w_6314,G159_8,G100_8,G100_11,_w_8940,_w_6430,_w_4527,G100_14,n1181,G100_16,_w_6724,_w_3978,G100_17,G100_19,G109_11,G100_18,G100_21,_w_3846,_w_7969,_w_7646,_w_6559,n991,n253_3,n744_0,n744_3,_w_6514,n744_4,G5293_2,_w_4273,n439_0,G100_6,G159_1,_w_4170,n439_1,_w_8782,_w_5343,n439_2,n439_3,G126_1,n749_1,n442_3,n442_5,n802_6,_w_6939,_w_4500,_w_7795,n442_6,n443_2,_w_3591,n443_3,n448_0,n448_1,_w_4313,n448_3,G5253_0,_w_8950,G5253_5,_w_4387,n450_1,_w_4784,G5260_0,_w_4091,G5260_2,n486,n451_0,G159_6,n451_5,n1239,n452_1,n453_0,n453_1,_w_5103,n457_1,_w_5776,_w_3632,n568,n457_2,n458_0,n458_1,_w_8102,_w_3963,n458_2,G105_5,n459_1,n459_2,_w_3462,n462_1,_w_4244,n462_2,_w_7076,n462_3,_w_8735,_w_6390,_w_4715,n464_0,n464_1,_w_4727,G161_5,n464_2,_w_5686,n465_3,n1152,_w_4075,n466_0,_w_7859,n345,n466_1,_w_6011,G166_0,n618,_w_3917,_w_8075,_w_4511,n476_2,n1289_1,_w_3641,n689_0,_w_8965,n271,_w_4837,n469_2,n469_3,_w_5295,n469_5,_w_4544,_w_4847,_w_4962,_w_6165,_w_3397,_w_4207,n472_0,n472_1,_w_5239,G5261_1,_w_5011,G90_4,n472_2,_w_6240,n472_3,_w_8138,_w_4683,_w_8766,n472_5,_w_4563,n472_6,n710,n472_7,n473_0,_w_4476,n1440_0,n474_1,n1434_1,_w_4909,n485_0,n466,n478_1,_w_4650,_w_4976,n594_0,_w_8161,_w_4724,_w_3994,n594_1,n763_0,_w_6853,n763_1,n503_0,n503_1,_w_6869,G139_0,_w_4288,n728_1,_w_7694,G139_4,_w_6416,G139_5,_w_6946,n600_1,n728_0,n974,G5255_2,_w_8977,_w_5991,_w_4679,_w_7789,G5255_3,G5255_4,G5255_5,_w_7470,n509_0,_w_8967,_w_8139,_w_7394,G5262_0,_w_4140,n387,n509_1,G64_0,_w_3474,G64_1,_w_7889,_w_7501,_w_5317,G100_10,_w_3809,_w_4228,_w_4696,G64_3,_w_3689,_w_3863,_w_4747,_w_4589,G64_5,n645,_w_4159,_w_5325,n1068,n900,G64_6,_w_5921,_w_5002,G64_7,G64_8,G64_13,G64_14,G98_10,G64_15,_w_8635,G64_16,G64_17,n1470,G159_5,G64_19,G64_20,G64_23,_w_7890,n997,_w_4280,G64_25,G94_3,_w_8809,_w_8235,G94_5,G94_7,_w_6326,_w_5092,G94_8,_w_3368,n542_2,G94_9,G94_11,G94_12,_w_4869,n465_2,n518_1,G5254_5,n524_1,_w_5669,n337_1,n530_0,n530_1,n1081,_w_3634,n534_0,_w_6563,_w_4695,n534_1,n547_1,_w_8517,_w_3445,G66_2,_w_3933,_w_4951,G66_3,G177_11,_w_4425,G94_10,_w_3877,n476_0,G66_4,G163_2,_w_4106,n586_0,_w_3512,n394_2,_w_4149,_w_4603,n586_2,n586_3,n586_4,n586_5,_w_4618,n586_6,n198,_w_3965,_w_8328,_w_7920,n586_7,_w_5828,_w_3655,n542_4,_w_5752,_w_3907,n1431,n542_5,n588_0,n588_1,_w_4705,n588_4,n588_5,n588_7,_w_6467,_w_6188,n449_1,n588_8,_w_4697,n588_11,G5293_1,G5293_4,n597_0,G123_3,n597_2,_w_6168,G5293_5,_w_3982,G115_0,_w_7665,G115_1,_w_4323,_w_6456,G115_3,_w_7591,G115_4,n607_3,_w_5513,n731_0,G172_4,_w_3563,n226,_w_4711,n390,n610_0,n610_1,n617_1,n485_1,n620_0,n620_1,_w_5824,G15_0,n327_0,_w_7090,n327_1,n640_0,_w_8703,_w_7158,_w_5022,G5258_1,n640_1,_w_6040,_w_5581,n640_2,G40_1,_w_4449,_w_5151,n444_1,_w_6692,_w_4774,n665_0,_w_6981,n666_1,n488_0,n1303_3,G82_0,G5250_1,n686_2,n1095,n886,n686_3,_w_6403,n744_6,_w_3648,_w_4296,_w_8282,n401_0,_w_7710,G90_8,n346_2,n701_1,_w_4635,_w_8349,_w_6915,n918,n710_1,n1395,n719_0,_w_5433,_w_4351,_w_3836,_w_4675,G76_1,n734_0,_w_6601,n737_1,_w_3751,_w_4908,_w_6703,n786_0,_w_7777,_w_3532,_w_4084,_w_5305,n477_0,G144_1,n752_1,G163_3,n760_0,_w_7599,n773_0,_w_5213,_w_3416,n773_2,n773_4,_w_4926,_w_6207,_w_4452,n773_7,_w_3999,n1324_1,_w_5520,_w_4470,_w_5255,n527_0,G177_28,_w_3838,n527_1,n789_0,_w_4521,_w_3415,_w_3467,_w_4403,_w_8964,n412,_w_4996,n789_1,G75_0,G101_13,_w_3609,G75_1,_w_7548,G111_0,n1350_1,n802_1,_w_6968,n802_4,n802_5,_w_3743,_w_7460,n1320_0,n858,_w_4175,n802_9,_w_6185,_w_4860,_w_6624,_w_6574,n802_11,G130_0,n804_0,_w_7517,_w_6455,n804_3,_w_5548,_w_4345,n1215,n804_5,_w_4039,n804_6,n804_10,_w_6356,n813_4,n813_5,_w_8855,n659,n813_11,n813_6,n813_8,n815_1,_w_3750,n911,n815_2,n275,n815_5,n815_6,_w_6453,n815_7,n815_9,n1244_1,n902,n393_1,_w_6930,G142_0,G161_6,G142_2,_w_4999,G176_1,_w_5844,G176_2,G176_3,G176_4,_w_8317,_w_7068,_w_6291,G176_7,_w_3537,n569,n231,G176_9,n577,G176_11,G176_13,G176_14,G176_15,_w_4008,G176_16,G176_18,n831,G176_20,G176_21,G176_22,_w_5185,G176_24,n1250_0,_w_5046,_w_3794,_w_8373,G176_25,G176_26,_w_8389,G1_0,G176_29,n689_1,G176_30,_w_7979,_w_7754,G176_31,n632_8,G176_33,n496,_w_3590,G176_34,G128_5,G176_35,_w_4271,G176_39,_w_8848,G176_40,_w_4065,_w_4415,G176_41,G176_45,n1327,G176_47,G176_48,_w_4614,G176_49,_w_4283,G176_51,G176_53,G102_3,_w_4483,_w_7388,_w_3831,G102_4,G102_7,G102_8,G102_9,G102_10,_w_3898,_w_6726,G102_11,G102_13,_w_8388,G130_5,G102_14,_w_5442,n607_1,n536,G102_15,_w_8403,n545,G102_16,G102_17,_w_4946,n397,G102_18,G90_0,_w_3441,_w_7525,G90_1,G90_2,G90_3,G101_14,G90_5,G90_6,G90_11,_w_6851,G5_0,_w_8739,_w_8442,_w_8164,n959_0,n386_1,n203,n386_4,G147_1,_w_4315,_w_7973,G147_2,G177_3,G147_3,_w_6349,_w_4390,G147_5,_w_8342,_w_4088,_w_7074,n545_0,n545_1,n545_2,_w_4642,G64_10,_w_3364,G128_6,_w_3366,_w_7706,_w_5642,_w_3367,_w_6994,_w_3953,_w_6260,_w_3370,_w_7948,_w_3373,_w_8470,_w_7447,_w_3376,_w_4956,_w_3379,_w_7103,n992,_w_3380,_w_5460,_w_3381,_w_5477,_w_3384,_w_3385,_w_3386,_w_3559,_w_8884,_w_3682,_w_3389,_w_6407,_w_3390,_w_5593,_w_3394,_w_5766,n391_0,n1463,_w_4152,_w_3395,n518,_w_3396,_w_3399,_w_5120,_w_3401,_w_3402,_w_3403,_w_5908,G102_6,_w_3404,_w_3405,_w_3407,_w_4096,_w_3466,_w_6969,n764,_w_3408,n1397,_w_3409,n630_11,_w_3411,_w_6002,_w_3414,_w_8687,G123_6,n749_0,_w_3421,_w_3422,_w_4687,_w_3423,_w_8316,_w_3424,n586,_w_4491,_w_4015,_w_5621,n1398_1,_w_4672,n293,_w_3425,_w_7774,_w_4739,_w_3426,_w_8133,_w_3429,_w_3431,n374_1,_w_3432,n861,_w_3433,_w_3435,_w_3436,_w_4311,_w_3437,n442_4,_w_3438,_w_3439,_w_6536,n346_1,_w_3440,_w_4298,_w_3442,n308,_w_3443,_w_4037,_w_8604,_w_5102,_w_3444,_w_3448,_w_8883,_w_3449,_w_4788,_w_3451,_w_7703,_w_4922,_w_3452,_w_4738,_w_4218,n1321,_w_3454,_w_3457,_w_3461,_w_3564,G123_7,n337_0,_w_3464,_w_3465,_w_3468,_w_6634,_w_3469,_w_3470,_w_3889,_w_3471,_w_6746,_w_3472,n1335,_w_3475,_w_3476,G174_20,_w_3477,_w_7163,_w_3478,n566,n841,_w_3902,_w_3480,G158_15,_w_3482,n456_1,_w_4997,_w_7541,_w_3483,_w_8219,_w_3485,_w_3487,n429_0,_w_3490,_w_6613,_w_3492,_w_3493,_w_6548,_w_3494,_w_3497,_w_5191,_w_3498,_w_8465,_w_6252,_w_5167,_w_3500,_w_3501,_w_6546,_w_3575,_w_3502,_w_6823,_w_3504,n515_0,_w_5044,_w_5364,_w_3507,_w_8926,_w_7917,_w_7536,_w_6600,_w_3765,G5292_5,_w_3508,_w_3654,n564,_w_3514,_w_7793,_w_3516,_w_3517,_w_7445,_w_3518,_w_4849,_w_3519,G96_4,_w_3520,_w_3521,_w_5045,_w_8837,_w_5465,G5258_0,G5261_0,_w_3522,n1294,i_G114,_w_3524,_w_3525,n421_2,_w_3526,_w_3541,_w_3531,_w_5466,_w_4628,_w_3533,_w_3534,_w_8845,G5251_2,G126_9,_w_3926,_w_3538,_w_6973,n752,_w_3539,_w_3543,_w_8200,_w_3545,_w_4914,_w_3546,_w_3550,_w_7205,_w_3712,_w_7530,_w_3551,_w_3552,n698_1,_w_3553,_w_3734,n552_25,_w_3554,_w_3556,_w_5704,_w_3557,_w_3562,_w_3658,_w_8281,n582,G124_16,_w_4541,_w_3565,_w_7696,_w_4105,_w_6904,_w_4130,_w_3566,n630_2,G5253_2,_w_3567,G90_9,_w_3569,_w_6753,_w_3571,_w_3453,_w_3576,_w_3580,_w_3581,_w_3582,_w_7316,_w_3584,_w_4027,n687,_w_3585,_w_4979,_w_3587,n456_5,_w_3589,_w_5653,_w_3592,_w_8711,G5221_10,_w_4457,_w_3594,_w_7457,_w_3596,_w_3598,_w_8069,_w_3599,_w_6334,_w_3603,_w_6183,_w_3604,_w_4945,n469_8,_w_5072,G96_9,G139_1,_w_3607,n554,_w_4885,_w_3608,_w_3610,_w_3612,_w_4089,_w_3613,_w_4343,_w_3614,_w_3616,n412_1,_w_3621,_w_4110,n495,_w_4225,n1371,_w_3626,G113_4,_w_3631,_w_7028,_w_6181,n397_0,_w_3633,_w_4262,_w_8571,_w_3635,_w_8400,_w_3637,_w_5316,n1102,G22_0,G105_4,_w_3639,_w_3644,_w_6124,_w_4189,_w_3647,_w_3649,_w_4932,_w_3651,_w_8930,_w_5947,_w_3652,_w_6014,_w_3656,_w_7409,_w_5632,_w_5271,n234_1,_w_4671,_w_4913,_w_8617,_w_3660,_w_3586,_w_3661,G103_12,_w_3662,_w_3665,_w_3669,_w_7422,_w_3671,_w_4540,_w_8483,_w_3674,n234_0,_w_3681,_w_7346,_w_3683,n949,_w_3685,_w_3687,_w_3690,_w_3691,_w_3915,_w_3693,_w_3694,_w_3699,n906,_w_3700,_w_7913,_w_3744,n806,n1188,_w_4494,_w_3701,_w_4684,_w_8694,_w_3703,_w_4607,G64_12,n386_0,_w_3704,_w_3705,_w_4782,_w_3968,_w_3710,n250,_w_3711,_w_8923,_w_8007,_w_3713,_w_3714,_w_3716,_w_6193,n633,_w_3717,_w_3719,_w_6929,_w_4814,_w_3722,_w_3723,_w_3724,_w_3726,_w_7621,_w_3727,n479_2,_w_3728,_w_3730,_w_4197,G158_6,_w_4665,_w_7728,G5229_0,_w_3813,_w_3732,_w_8280,_w_8229,n462_0,_w_4772,G5258_5,_w_3735,_w_5212,G107_12,_w_3737,_w_3739,_w_3746,_w_8857,_w_3748,_w_3752,_w_3755,_w_3756,_w_8397,_w_3757,n1300_0,n1410,_w_5031,_w_3758,n920,_w_3759,_w_3760,_w_4064,_w_8345,_w_7966,_w_3761,n1217,_w_4142,_w_3764,_w_8246,_w_4901,n253_1,_w_4087,_w_5706,n236,_w_3771,G157_2,_w_5019,_w_8713,_w_5086,_w_5354,G174_2,n270,_w_3772,_w_3775,_w_3776,_w_8945,_w_5165,_w_3778,_w_3779,_w_3781,_w_3782,_w_3783,_w_5914,_w_3784,_w_3787,_w_6567,_w_3789,_w_5452,_w_3800,G160_15,_w_3801,_w_5020,_w_3410,_w_3803,_w_6383,_w_3374,_w_3806,_w_3808,_w_8487,_w_3812,_w_3815,n451_1,_w_3816,_w_5912,_w_3819,_w_3821,_w_4804,_w_8979,_w_8656,_w_7353,_w_6561,_w_6053,_w_3428,_w_3822,_w_3823,_w_3824,_w_3904,n1001,n739,_w_3825,_w_6128,G174_15,_w_3826,_w_3827,n855,n852,_w_3829,_w_3830,G125_1,_w_3835,_w_4528,n411,_w_3837,_w_3839,_w_8088,_w_7512,n537_5,_w_3840,_w_5544,_w_4126,_w_3841,_w_6575,_w_3842,_w_3843,n420,_w_3601,_w_4436,_w_4620,_w_3845,_w_3847,_w_7064,_w_3848,n465_1,_w_3849,_w_8814,_w_4435,_w_5897,_w_3851,n1131,n247,_w_3852,_w_6717,_w_3855,_w_6010,n1130,_w_3856,G101_5,_w_3857,_w_6294,_w_3859,G100_12,_w_3860,_w_5564,_w_3862,_w_8938,_w_6279,_w_6160,_w_3866,_w_8252,_w_3867,_w_7642,_w_5060,n588_9,_w_3868,_w_7467,_w_5220,n1308_1,_w_3870,_w_3872,_w_6528,_w_3873,_w_3876,_w_6064,_w_3882,_w_3883,_w_3887,_w_5655,_w_4751,_w_3888,_w_3890,_w_7240,_w_3891,_w_3892,_w_3900,_w_4501,_w_3895,n351,_w_5043,_w_3897,_w_4924,_w_8454,_w_3899,_w_3903,n433,_w_3905,_w_3906,_w_3908,_w_3909,_w_5310,_w_3910,_w_6348,_w_4519,_w_3912,_w_3916,_w_6246,_w_4656,_w_3918,n469_7,_w_3919,_w_5263,_w_4226,_w_3773,_w_4405,_w_3920,_w_7520,_w_3924,_w_3927,_w_3934,_w_3936,_w_6135,G148_5,_w_3939,_w_7503,_w_3944,n529,_w_4127,G172_6,_w_3945,_w_3947,_w_4188,_w_4382,n245,_w_3948,n774,_w_3949,_w_3954,_w_4773,_w_5399,_w_3955,_w_4838,_w_3957,_w_4488,_w_7620,_w_3961,_w_8486,_w_4641,_w_8661,_w_3967,_w_3970,_w_3763,_w_4674,n1375,_w_3740,_w_3972,_w_8725,_w_3973,_w_3974,_w_3975,_w_3977,_w_3979,_w_6248,_w_3981,_w_6907,_w_3983,_w_3984,_w_3985,_w_3987,_w_3989,_w_8167,_w_7654,_w_7305,_w_5841,_w_3990,_w_6495,_w_5401,n1380,_w_3992,_w_6769,n418_0,n1324,G124_2,_w_3993,n1019,_w_3995,_w_8512,_w_3996,_w_6942,_w_3998,n518_0,_w_4001,_w_4002,_w_6748,_w_4003,_w_7266,_w_5436,_w_5179,_w_4004,_w_4154,_w_4006,_w_4009,_w_4012,_w_5983,n832,_w_4013,_w_6713,_w_4959,_w_4019,_w_5759,_w_4020,_w_4024,_w_4032,_w_8107,_w_7936,_w_3925,_w_4033,_w_4272,_w_4034,_w_3736,_w_4129,_w_4036,_w_4040,n340,_w_4046,G177_17,_w_4808,_w_4047,_w_4214,_w_4048,_w_4049,_w_4052,_w_6992,_w_4054,_w_7352,_w_6275,_w_4055,_w_4058,_w_3922,_w_4801,_w_7643,_w_4061,_w_4063,_w_4067,n261,_w_4068,_w_7082,_w_4274,_w_4069,_w_4070,_w_4072,_w_4894,_w_4073,_w_4631,_w_4074,_w_4845,n600_0,G109_9,_w_4077,_w_3670,_w_4082,_w_4090,_w_8378,_w_8236,_w_5098,n653,_w_4092,_w_4477,_w_4463,_w_4093,_w_4094,_w_4095,_w_4098,_w_6752,_w_4100,_w_4101,_w_6788,_w_4102,_w_4107,_w_7419,_w_4954,_w_3577,_w_4109,_w_6817,_w_3769,_w_4111,G64_2,_w_4112,_w_4116,n444_0,_w_4118,_w_8762,_w_4868,_w_4119,_w_5199,_w_4132,_w_3657,_w_4134,_w_4136,_w_4138,_w_4139,_w_5204,_w_4143,n500_1,_w_4208,G158_27,_w_4682,_w_5724,_w_4144,_w_8343,_w_4592,_w_4148,_w_6186,n1142,_w_4150,_w_4896,_w_3548,_w_4155,_w_5859,_w_4941,_w_4156,G115_2,_w_4157,G101_10,_w_4158,_w_4043,_w_4164,n709,_w_4166,_w_4167,_w_4168,G83_0,_w_4371,n542_3,_w_4169,_w_4172,_w_4174,_w_4178,_w_4235,_w_5052,_w_8618,_w_7432,_w_4181,_w_8701,_w_6687,G71_0,n938,_w_4183,_w_4185,_w_7121,n1386_0,_w_4186,n1198_1,_w_4190,_w_4327,n1293,_w_4191,_w_5009,_w_3527,_w_4192,_w_4195,_w_5833,n1261,G123_5,_w_4512,_w_4196,_w_8907,n304,_w_4198,_w_4787,_w_4202,_w_6037,G170_2,G174_13,G158_26,_w_4203,n670_0,_w_4204,_w_4209,_w_4212,_w_6890,_w_4783,_w_4217,_w_4222,_w_7032,_w_4224,_w_3369,_w_4227,_w_4229,G137_2,_w_4337,_w_5740,_w_4230,_w_7699,_w_5275,_w_4275,_w_4232,n552_16,_w_4233,_w_4234,_w_7833,_w_4237,_w_4242,_w_5961,_w_3901,n1104,n388,_w_4243,_w_7468,_w_4246,_w_4249,_w_4252,_w_4219,_w_4253,_w_4255,n1305_1,_w_4256,_w_4258,n658_0,_w_4263,_w_4264,_w_7893,_w_4276,_w_4278,_w_4279,_w_8034,_w_5622,_w_4281,n425,_w_4282,_w_8263,G163_9,_w_4284,_w_5733,_w_4791,_w_4286,n643_2,G138_2,_w_4289,_w_6297,n371,_w_4254,_w_4291,_w_4293,_w_4505,_w_4294,n1428_0,_w_4297,_w_6242,_w_4921,_w_4299,_w_6394,_w_4555,_w_3561,_w_4622,_w_8214,_w_4300,_w_4301,_w_4865,n718,_w_4302,_w_4551,_w_4303,_w_4947,_w_4304,_w_4305,_w_4308,_w_4310,_w_8116,_w_4314,_w_6977,_w_4316,_w_5689,_w_4318,_w_4324,_w_6319,_w_4328,n1185,n977,_w_4329,_w_5846,_w_5245,_w_3388,_w_4668,n387_2,_w_4332,_w_5217,_w_4336,_w_4424,_w_4338,n604,_w_4340,_w_4341,G176_43,_w_4344,_w_6250,_w_4657,_w_4352,_w_4359,_w_6049,_w_3828,_w_4493,_w_4360,G174_4,n1350,_w_4361,_w_5836,_w_4362,_w_4461,_w_4363,_w_4364,_w_6404,n783_0,_w_4366,_w_4368,_w_4369,_w_4370,_w_7027,_w_4374,_w_7328,n1171,_w_4375,_w_8803,_w_4376,_w_4377,_w_4379,_w_4383,_w_4385,_w_6921,_w_4388,_w_4389,_w_4392,_w_4393,_w_6409,_w_4394,_w_5083,_w_4035,_w_4396,_w_5995,_w_5925,_w_4398,_w_4400,G42_0,_w_4402,_w_8357,_w_4404,_w_4407,G124_6,_w_4408,_w_4410,_w_6937,_w_3636,_w_4411,_w_4413,_w_4417,G96_13,_w_4420,_w_8488,_w_4423,_w_6568,_w_4427,_w_5688,_w_5114,n460,_w_4428,_w_4432,_w_4010,_w_4433,_w_4434,n815_0,_w_4437,_w_4439,_w_3720,_w_4890,_w_4441,_w_7146,_w_6337,_w_4180,_w_4442,_w_7119,_w_4446,_w_4447,n197,_w_4743,_w_6178,_w_4450,_w_7109,n199,_w_4451,_w_7944,_w_7047,_w_5900,_w_4051,_w_4453,_w_7148,n707,_w_4454,_w_4456,n427_0,_w_4458,_w_4633,n586_8,_w_4459,G103_1,_w_4460,_w_5106,_w_4465,_w_4467,n685,_w_4468,n1381,_w_4471,_w_4472,n479_3,_w_4473,n688,_w_4474,_w_7856,n235,_w_4482,G102_12,_w_4485,_w_4530,_w_4490,_w_4690,_w_4762,_w_4492,n469_1,_w_4495,_w_5233,_w_4496,n509,_w_4498,_w_4499,_w_5847,_w_5583,_w_4502,_w_4987,_w_4503,_w_8324,_w_3937,_w_4504,_w_4011,_w_4506,_w_4509,_w_5340,_w_4510,_w_4816,n1367,n469_0,_w_4513,_w_5734,_w_4017,_w_4221,_w_4514,_w_4873,_w_4516,G66_6,_w_4517,G148_1,_w_4518,_w_4520,_w_4524,_w_4531,n1438,_w_4533,_w_4673,_w_7894,_w_4507,_w_4534,_w_7876,_w_4536,_w_6309,G168_7,_w_4537,_w_4539,_w_7545,_w_7218,n733,_w_4543,_w_4545,_w_4546,_w_4547,n1314_1,_w_4248,_w_4548,_w_4549,_w_6330,_w_4550,_w_4554,_w_8542,_w_4556,_w_4558,_w_6147,_w_4732,_w_4559,_w_4933,n464_4,_w_4560,n565_0,_w_4561,_w_7197,_w_4562,_w_4567,_w_4569,_w_4572,_w_4573,_w_4576,_w_4469,_w_3535,_w_4577,_w_4581,_w_4584,_w_4586,n353,G162_1,_w_4596,n627,_w_4587,n479_0,_w_4591,_w_4593,_w_6715,G88_2,_w_4597,_w_4598,_w_4599,_w_8109,_w_4602,_w_4605,G5199_0,_w_4678,_w_8521,_w_6253,_w_4608,n802_2,_w_4611,_w_4613,_w_4445,_w_4615,_w_6121,_w_4617,_w_4619,G123_9,_w_4621,_w_4623,_w_4625,_w_4626,_w_4644,_w_4712,_w_4627,_w_6592,_w_5798,_w_4629,_w_4630,n725,_w_4918,_w_6849,n400_4,_w_4632,_w_4637,_w_4639,_w_6229,_w_6024,n667_1,_w_4643,_w_4645,_w_7949,_w_5994,_w_4647,_w_4919,_w_7528,_w_4651,_w_4251,_w_4654,_w_3747,_w_3618,_w_4659,_w_4660,_w_3547,_w_4936,_w_4663,_w_4666,n285,_w_4667,_w_3459,_w_4669,_w_8520,_w_7202,_w_4670,_w_4676,_w_4685,_w_4686,n1447_2,_w_4689,_w_4691,_w_4692,_w_6304,_w_4694,_w_4698,_w_5008,_w_4701,_w_6911,_w_4759,_w_6028,_w_4702,n1076,_w_4775,_w_7872,_w_5006,_w_5896,_w_4703,_w_4704,n871,_w_4707,_w_4708,n814,_w_4103,_w_4709,_w_4859,_w_4710,_w_6012,_w_4716,_w_7052,n253_2,_w_4717,_w_8829,_w_8010,_w_4718,G176_5,_w_4721,G173_11,_w_4722,_w_8127,_w_4725,_w_5788,_w_4726,_w_3686,_w_4729,G5255_0,_w_4731,_w_8362,_w_4733,_w_7289,_w_5215,_w_4737,_w_3709,_w_4740,_w_7256,n1376,_w_4741,_w_5939,_w_4744,_w_5314,G5258_3,_w_4079,n552_23,_w_4746,_w_4750,_w_5495,_w_4753,G5259_1,_w_4755,G174_12,_w_4756,n442_7,_w_4757,_w_4760,_w_8942,_w_6418,_w_4331,_w_4761,_w_7590,_w_4763,G177_14,_w_4766,_w_7568,_w_4768,G163_13,_w_4770,G160_13,_w_3627,_w_4777,_w_4779,_w_4780,_w_4781,_w_4789,_w_8201,_w_6041,n885,_w_4790,_w_7130,n725_1,_w_4793,n434_1,n979,_w_4795,_w_4797,_w_8029,_w_5208,_w_4798,_w_4802,_w_4803,_w_4165,_w_4806,_w_4807,_w_4811,_w_4812,_w_7164,_w_4818,_w_8435,_w_4821,_w_4822,_w_4823,_w_4825,_w_7152,n396,_w_4828,_w_4831,_w_6223,_w_4833,n428_0,_w_4834,_w_5592,n393,_w_4358,_w_4840,_w_4841,_w_4842,n546,_w_4844,_w_8636,_w_7935,_w_4846,_w_4855,G107_7,_w_4856,_w_7199,_w_4858,_w_4861,_w_7034,_w_4862,_w_7288,_w_4864,_w_4867,_w_8165,_w_4870,_w_5058,_w_4871,_w_4579,_w_4872,_w_4373,_w_4875,_w_4876,n725_0,G64_4,_w_4878,_w_3572,_w_4879,_w_8399,_w_4882,_w_4754,_w_4883,_w_4886,n338,_w_4887,_w_4893,_w_4321,_w_4897,_w_4898,_w_4903,_w_4133,_w_4904,n262,_w_4905,_w_4910,_w_7810,_w_4911,_w_4915,_w_7302,_w_3486,_w_4916,_w_4920,n192,_w_4927,n1144,_w_4928,_w_7327,n385,_w_4935,_w_4937,_w_8058,n864,_w_4938,_w_4942,_w_6585,_w_3811,_w_4943,_w_5822,G129_1,_w_4944,_w_7131,_w_6891,_w_4213,_w_4950,_w_7439,_w_5723,_w_4952,n1242,_w_4955,_w_7946,n456_3,_w_4961,_w_5699,_w_4960,n494_0,_w_4967,_w_4029,_w_4969,_w_6607,_w_4971,n1320,_w_4973,_w_6629,_w_4974,G175_2,_w_4978,_w_4981,_w_4045,_w_4983,_w_6206,G176_28,_w_5067,_w_4984,n982,_w_4985,_w_4986,n400_3,_w_4988,_w_4990,_w_7600,_w_4992,_w_4993,_w_3791,_w_4995,_w_5000,_w_8206,G90_7,_w_5001,_w_3446,n657,_w_5017,_w_3495,G5259_5,_w_5021,_w_5025,_w_5026,G172_1,n572,_w_3914,_w_5027,_w_5032,_w_6576,G168_10,_w_5033,_w_8607,_w_7414,_w_5037,_w_5038,_w_5647,_w_5039,_w_8882,_w_5042,n611,_w_5048,_w_3969,_w_5050,G160_2,n432_2,_w_5054,_w_5056,G158_18,_w_5059,_w_5062,_w_5063,_w_5066,n586_9,_w_5070,_w_5071,_w_5076,_w_5077,_w_5661,_w_5078,_w_5081;

  bfr _b_7561(.a(_w_8986),.q(_w_8987));
  bfr _b_7559(.a(_w_8984),.q(_w_8985));
  bfr _b_7555(.a(_w_8980),.q(_w_8981));
  bfr _b_7550(.a(_w_8975),.q(_w_8976));
  bfr _b_7548(.a(_w_8973),.q(_w_8974));
  bfr _b_7545(.a(_w_8970),.q(_w_8971));
  bfr _b_7544(.a(_w_8969),.q(_w_8970));
  bfr _b_7542(.a(_w_8967),.q(_w_8968));
  bfr _b_7539(.a(_w_8964),.q(_w_8965));
  bfr _b_7538(.a(_w_8963),.q(_w_8964));
  bfr _b_7534(.a(_w_8959),.q(_w_8960));
  bfr _b_7533(.a(_w_8958),.q(_w_8959));
  bfr _b_7531(.a(G99),.q(_w_8957));
  bfr _b_7530(.a(G98),.q(_w_8955));
  bfr _b_7529(.a(_w_8954),.q(_w_8952));
  bfr _b_7528(.a(_w_8953),.q(_w_8954));
  bfr _b_7527(.a(G97),.q(_w_8953));
  bfr _b_7525(.a(G95),.q(_w_8951));
  bfr _b_7523(.a(G93),.q(_w_8949));
  bfr _b_7520(.a(_w_8945),.q(_w_8944));
  bfr _b_7519(.a(G9),.q(_w_8945));
  bfr _b_7518(.a(_w_8943),.q(_w_8942));
  bfr _b_7517(.a(G89),.q(_w_8943));
  bfr _b_7510(.a(_w_8935),.q(_w_8936));
  bfr _b_7507(.a(_w_8932),.q(_w_8933));
  bfr _b_7504(.a(_w_8929),.q(_w_8930));
  bfr _b_7503(.a(_w_8928),.q(_w_8929));
  bfr _b_7500(.a(_w_8925),.q(_w_8926));
  bfr _b_7497(.a(_w_8922),.q(_w_8923));
  bfr _b_7495(.a(_w_8920),.q(_w_8921));
  bfr _b_7494(.a(_w_8919),.q(_w_8920));
  bfr _b_7493(.a(_w_8918),.q(_w_8919));
  bfr _b_7492(.a(_w_8917),.q(_w_8918));
  bfr _b_7491(.a(_w_8916),.q(_w_8917));
  bfr _b_7490(.a(_w_8915),.q(_w_8916));
  bfr _b_7487(.a(_w_8912),.q(_w_8913));
  bfr _b_7484(.a(_w_8909),.q(_w_8910));
  bfr _b_7481(.a(_w_8906),.q(_w_8907));
  bfr _b_7476(.a(_w_8901),.q(_w_8902));
  bfr _b_7475(.a(_w_8900),.q(_w_8901));
  bfr _b_7473(.a(_w_8898),.q(_w_8899));
  bfr _b_7471(.a(_w_8896),.q(_w_8897));
  bfr _b_7470(.a(_w_8895),.q(_w_8896));
  bfr _b_7469(.a(_w_8894),.q(_w_8895));
  bfr _b_7463(.a(_w_8888),.q(_w_8889));
  bfr _b_7461(.a(_w_8886),.q(_w_8887));
  bfr _b_7459(.a(_w_8884),.q(_w_8885));
  bfr _b_7457(.a(_w_8882),.q(_w_8883));
  bfr _b_7456(.a(_w_8881),.q(_w_8882));
  bfr _b_7454(.a(_w_8879),.q(_w_8880));
  bfr _b_7453(.a(_w_8878),.q(_w_8879));
  bfr _b_7452(.a(_w_8877),.q(_w_8878));
  bfr _b_7450(.a(G86),.q(_w_8876));
  bfr _b_7441(.a(_w_8866),.q(_w_8867));
  bfr _b_7437(.a(_w_8862),.q(_w_8863));
  bfr _b_7436(.a(_w_8861),.q(_w_8862));
  bfr _b_7434(.a(_w_8859),.q(_w_8860));
  bfr _b_7425(.a(_w_8850),.q(_w_8851));
  bfr _b_7423(.a(_w_8848),.q(_w_8849));
  bfr _b_7421(.a(_w_8846),.q(_w_8847));
  bfr _b_7420(.a(_w_8845),.q(_w_8846));
  bfr _b_7415(.a(_w_8840),.q(_w_8807));
  bfr _b_7414(.a(_w_8839),.q(_w_8840));
  bfr _b_7411(.a(_w_8836),.q(_w_8837));
  bfr _b_7409(.a(_w_8834),.q(_w_8835));
  bfr _b_7408(.a(_w_8833),.q(_w_8834));
  bfr _b_7406(.a(_w_8831),.q(_w_8832));
  bfr _b_7404(.a(_w_8829),.q(_w_8830));
  bfr _b_7403(.a(_w_8828),.q(_w_8829));
  bfr _b_7402(.a(_w_8827),.q(_w_8828));
  bfr _b_7401(.a(_w_8826),.q(_w_8827));
  bfr _b_7397(.a(_w_8822),.q(_w_8823));
  bfr _b_7396(.a(_w_8821),.q(_w_8822));
  bfr _b_7395(.a(_w_8820),.q(_w_8821));
  bfr _b_7394(.a(_w_8819),.q(_w_8820));
  bfr _b_7393(.a(_w_8818),.q(_w_8819));
  bfr _b_7392(.a(_w_8817),.q(_w_8818));
  bfr _b_7389(.a(_w_8814),.q(_w_8815));
  bfr _b_7387(.a(_w_8812),.q(_w_8813));
  bfr _b_7386(.a(_w_8811),.q(_w_8812));
  bfr _b_7381(.a(_w_8806),.q(_w_8773));
  bfr _b_7379(.a(_w_8804),.q(_w_8805));
  bfr _b_7376(.a(_w_8801),.q(_w_8802));
  bfr _b_7373(.a(_w_8798),.q(_w_8799));
  bfr _b_7372(.a(_w_8797),.q(_w_8798));
  bfr _b_7369(.a(_w_8794),.q(_w_8795));
  bfr _b_7368(.a(_w_8793),.q(_w_8794));
  bfr _b_7367(.a(_w_8792),.q(_w_8793));
  bfr _b_7365(.a(_w_8790),.q(_w_8791));
  bfr _b_7361(.a(_w_8786),.q(_w_8787));
  bfr _b_7360(.a(_w_8785),.q(_w_8786));
  bfr _b_7357(.a(_w_8782),.q(_w_8783));
  bfr _b_7486(.a(_w_8911),.q(_w_8912));
  bfr _b_7355(.a(_w_8780),.q(_w_8781));
  bfr _b_7350(.a(_w_8775),.q(_w_8776));
  bfr _b_7349(.a(_w_8774),.q(_w_8775));
  bfr _b_7347(.a(_w_8772),.q(_w_8739));
  bfr _b_7345(.a(_w_8770),.q(_w_8771));
  bfr _b_7340(.a(_w_8765),.q(_w_8766));
  bfr _b_7335(.a(_w_8760),.q(_w_8761));
  bfr _b_7334(.a(_w_8759),.q(_w_8760));
  bfr _b_7333(.a(_w_8758),.q(_w_8759));
  bfr _b_7332(.a(_w_8757),.q(_w_8758));
  bfr _b_7331(.a(_w_8756),.q(_w_8757));
  bfr _b_7329(.a(_w_8754),.q(_w_8755));
  bfr _b_7328(.a(_w_8753),.q(_w_8754));
  bfr _b_7326(.a(_w_8751),.q(_w_8752));
  bfr _b_7325(.a(_w_8750),.q(_w_8751));
  bfr _b_7322(.a(_w_8747),.q(_w_8748));
  bfr _b_7319(.a(_w_8744),.q(_w_8745));
  bfr _b_7313(.a(_w_8738),.q(_w_8706));
  bfr _b_7312(.a(_w_8737),.q(_w_8738));
  bfr _b_7308(.a(_w_8733),.q(_w_8734));
  bfr _b_7307(.a(_w_8732),.q(_w_8733));
  bfr _b_7306(.a(_w_8731),.q(_w_8732));
  bfr _b_7303(.a(_w_8728),.q(_w_8729));
  bfr _b_7302(.a(_w_8727),.q(_w_8728));
  bfr _b_7301(.a(_w_8726),.q(_w_8727));
  bfr _b_7300(.a(_w_8725),.q(_w_8726));
  bfr _b_7295(.a(_w_8720),.q(_w_8721));
  bfr _b_7293(.a(_w_8718),.q(_w_8719));
  bfr _b_7291(.a(_w_8716),.q(_w_8717));
  bfr _b_7289(.a(_w_8714),.q(_w_8715));
  bfr _b_7288(.a(_w_8713),.q(_w_8714));
  bfr _b_7286(.a(_w_8711),.q(_w_8712));
  bfr _b_7280(.a(_w_8705),.q(_w_8673));
  bfr _b_7279(.a(_w_8704),.q(_w_8705));
  bfr _b_7278(.a(_w_8703),.q(_w_8704));
  bfr _b_7275(.a(_w_8700),.q(_w_8701));
  bfr _b_7273(.a(_w_8698),.q(_w_8699));
  bfr _b_7271(.a(_w_8696),.q(_w_8697));
  bfr _b_7266(.a(_w_8691),.q(_w_8692));
  bfr _b_7264(.a(_w_8689),.q(_w_8690));
  bfr _b_7263(.a(_w_8688),.q(_w_8689));
  bfr _b_7260(.a(_w_8685),.q(_w_8686));
  bfr _b_7255(.a(_w_8680),.q(_w_8681));
  bfr _b_7254(.a(_w_8679),.q(_w_8680));
  bfr _b_7251(.a(_w_8676),.q(_w_8677));
  bfr _b_7247(.a(_w_8672),.q(_w_8671));
  bfr _b_7242(.a(_w_8667),.q(_w_8668));
  bfr _b_7240(.a(_w_8665),.q(_w_8666));
  bfr _b_7239(.a(_w_8664),.q(_w_8665));
  bfr _b_7238(.a(_w_8663),.q(_w_8664));
  bfr _b_7237(.a(_w_8662),.q(_w_8663));
  bfr _b_7236(.a(_w_8661),.q(_w_8662));
  bfr _b_7235(.a(_w_8660),.q(_w_8661));
  bfr _b_7234(.a(_w_8659),.q(_w_8660));
  bfr _b_7231(.a(_w_8656),.q(_w_8657));
  bfr _b_7230(.a(_w_8655),.q(_w_8656));
  bfr _b_7229(.a(_w_8654),.q(_w_8655));
  bfr _b_7226(.a(_w_8651),.q(_w_8652));
  bfr _b_7223(.a(_w_8648),.q(_w_8649));
  bfr _b_7222(.a(_w_8647),.q(_w_8648));
  bfr _b_7216(.a(_w_8641),.q(_w_8642));
  bfr _b_7215(.a(_w_8640),.q(_w_8641));
  bfr _b_7212(.a(G79),.q(_w_8638));
  bfr _b_7211(.a(_w_8636),.q(_w_8603));
  bfr _b_7210(.a(_w_8635),.q(_w_8636));
  bfr _b_7200(.a(_w_8625),.q(_w_8626));
  bfr _b_7198(.a(_w_8623),.q(_w_8624));
  bfr _b_7196(.a(_w_8621),.q(_w_8622));
  bfr _b_7195(.a(_w_8620),.q(_w_8621));
  bfr _b_7192(.a(_w_8617),.q(_w_8618));
  bfr _b_7190(.a(_w_8615),.q(_w_8616));
  bfr _b_7188(.a(_w_8613),.q(_w_8614));
  bfr _b_7187(.a(_w_8612),.q(_w_8613));
  bfr _b_7186(.a(_w_8611),.q(_w_8612));
  bfr _b_7176(.a(_w_8601),.q(_w_8602));
  bfr _b_7175(.a(_w_8600),.q(_w_8601));
  bfr _b_7209(.a(_w_8634),.q(_w_8635));
  bfr _b_7174(.a(_w_8599),.q(_w_8600));
  bfr _b_7173(.a(_w_8598),.q(_w_8599));
  bfr _b_7170(.a(_w_8595),.q(_w_8596));
  bfr _b_7168(.a(_w_8593),.q(_w_8594));
  bfr _b_7166(.a(_w_8591),.q(_w_8592));
  bfr _b_7163(.a(_w_8588),.q(_w_8589));
  bfr _b_7162(.a(_w_8587),.q(_w_8588));
  bfr _b_7161(.a(_w_8586),.q(_w_8587));
  bfr _b_7160(.a(_w_8585),.q(_w_8586));
  bfr _b_7157(.a(_w_8582),.q(_w_8583));
  bfr _b_7155(.a(_w_8580),.q(_w_8581));
  bfr _b_7154(.a(_w_8579),.q(_w_8580));
  bfr _b_7153(.a(_w_8578),.q(_w_8579));
  bfr _b_7151(.a(_w_8576),.q(_w_8577));
  bfr _b_7149(.a(_w_8574),.q(_w_8575));
  bfr _b_7148(.a(_w_8573),.q(_w_8574));
  bfr _b_7147(.a(_w_8572),.q(_w_8573));
  bfr _b_7139(.a(_w_8564),.q(_w_8565));
  bfr _b_7136(.a(_w_8561),.q(_w_8562));
  bfr _b_7135(.a(_w_8560),.q(_w_8561));
  bfr _b_7297(.a(_w_8722),.q(_w_8723));
  bfr _b_7134(.a(_w_8559),.q(_w_8560));
  bfr _b_7133(.a(_w_8558),.q(_w_8559));
  bfr _b_7132(.a(_w_8557),.q(_w_8558));
  bfr _b_7131(.a(_w_8556),.q(_w_8557));
  bfr _b_7130(.a(_w_8555),.q(_w_8556));
  bfr _b_7129(.a(_w_8554),.q(_w_8555));
  bfr _b_7128(.a(_w_8553),.q(_w_8554));
  bfr _b_7124(.a(_w_8549),.q(_w_8550));
  bfr _b_7122(.a(_w_8547),.q(_w_8548));
  bfr _b_7121(.a(_w_8546),.q(_w_8547));
  bfr _b_7119(.a(_w_8544),.q(_w_8545));
  bfr _b_7118(.a(_w_8543),.q(_w_8544));
  bfr _b_7552(.a(_w_8977),.q(_w_8978));
  bfr _b_7114(.a(_w_8539),.q(_w_8540));
  bfr _b_7113(.a(_w_8538),.q(_w_8539));
  bfr _b_7111(.a(G76),.q(_w_8537));
  bfr _b_7110(.a(_w_8535),.q(_w_8502));
  bfr _b_7108(.a(_w_8533),.q(_w_8534));
  bfr _b_7105(.a(_w_8530),.q(_w_8531));
  bfr _b_7102(.a(_w_8527),.q(_w_8528));
  bfr _b_7094(.a(_w_8519),.q(_w_8520));
  bfr _b_7093(.a(_w_8518),.q(_w_8519));
  bfr _b_7092(.a(_w_8517),.q(_w_8518));
  bfr _b_7090(.a(_w_8515),.q(_w_8516));
  bfr _b_7087(.a(_w_8512),.q(_w_8513));
  bfr _b_7086(.a(_w_8511),.q(_w_8512));
  bfr _b_7083(.a(_w_8508),.q(_w_8509));
  bfr _b_7078(.a(_w_8503),.q(_w_8504));
  bfr _b_7077(.a(G75),.q(_w_8503));
  bfr _b_7076(.a(_w_8501),.q(_w_8468));
  bfr _b_7075(.a(_w_8500),.q(_w_8501));
  bfr _b_7073(.a(_w_8498),.q(_w_8499));
  bfr _b_7072(.a(_w_8497),.q(_w_8498));
  bfr _b_7100(.a(_w_8525),.q(_w_8526));
  bfr _b_7069(.a(_w_8494),.q(_w_8495));
  bfr _b_7068(.a(_w_8493),.q(_w_8494));
  bfr _b_7067(.a(_w_8492),.q(_w_8493));
  bfr _b_7064(.a(_w_8489),.q(_w_8490));
  bfr _b_7063(.a(_w_8488),.q(_w_8489));
  bfr _b_7062(.a(_w_8487),.q(_w_8488));
  bfr _b_7061(.a(_w_8486),.q(_w_8487));
  bfr _b_7057(.a(_w_8482),.q(_w_8483));
  bfr _b_7056(.a(_w_8481),.q(_w_8482));
  bfr _b_7465(.a(_w_8890),.q(_w_8891));
  bfr _b_7055(.a(_w_8480),.q(_w_8481));
  bfr _b_7050(.a(_w_8475),.q(_w_8476));
  bfr _b_7049(.a(_w_8474),.q(_w_8475));
  bfr _b_7048(.a(_w_8473),.q(_w_8474));
  bfr _b_7046(.a(_w_8471),.q(_w_8472));
  bfr _b_7045(.a(_w_8470),.q(_w_8471));
  bfr _b_7043(.a(G74),.q(_w_8469));
  bfr _b_7041(.a(_w_8466),.q(_w_8467));
  bfr _b_7039(.a(_w_8464),.q(_w_8465));
  bfr _b_7038(.a(_w_8463),.q(_w_8464));
  bfr _b_7037(.a(_w_8462),.q(_w_8463));
  bfr _b_7036(.a(_w_8461),.q(_w_8462));
  bfr _b_7035(.a(_w_8460),.q(_w_8461));
  bfr _b_7034(.a(_w_8459),.q(_w_8460));
  bfr _b_7032(.a(_w_8457),.q(_w_8458));
  bfr _b_7031(.a(_w_8456),.q(_w_8457));
  bfr _b_7028(.a(_w_8453),.q(_w_8454));
  bfr _b_7027(.a(_w_8452),.q(_w_8453));
  bfr _b_7026(.a(_w_8451),.q(_w_8452));
  bfr _b_7023(.a(_w_8448),.q(_w_8449));
  bfr _b_7020(.a(_w_8445),.q(_w_8446));
  bfr _b_7019(.a(_w_8444),.q(_w_8445));
  bfr _b_7017(.a(_w_8442),.q(_w_8443));
  bfr _b_7016(.a(_w_8441),.q(_w_8442));
  bfr _b_7015(.a(_w_8440),.q(_w_8441));
  bfr _b_7014(.a(_w_8439),.q(_w_8440));
  bfr _b_7217(.a(_w_8642),.q(_w_8643));
  bfr _b_7013(.a(_w_8438),.q(_w_8439));
  bfr _b_7009(.a(G73),.q(_w_8435));
  bfr _b_7007(.a(_w_8432),.q(_w_8433));
  bfr _b_7006(.a(_w_8431),.q(_w_8432));
  bfr _b_7005(.a(_w_8430),.q(_w_8431));
  bfr _b_7004(.a(_w_8429),.q(_w_8430));
  bfr _b_7003(.a(_w_8428),.q(_w_8429));
  bfr _b_7024(.a(_w_8449),.q(_w_8450));
  bfr _b_7002(.a(_w_8427),.q(_w_8428));
  bfr _b_7001(.a(_w_8426),.q(_w_8427));
  bfr _b_7000(.a(_w_8425),.q(_w_8426));
  bfr _b_6999(.a(_w_8424),.q(_w_8425));
  bfr _b_6998(.a(_w_8423),.q(_w_8424));
  bfr _b_6997(.a(_w_8422),.q(_w_8423));
  bfr _b_6994(.a(_w_8419),.q(_w_8420));
  bfr _b_6993(.a(_w_8418),.q(_w_8419));
  bfr _b_6992(.a(_w_8417),.q(_w_8418));
  bfr _b_6989(.a(_w_8414),.q(_w_8415));
  bfr _b_6988(.a(_w_8413),.q(_w_8414));
  bfr _b_6987(.a(_w_8412),.q(_w_8413));
  bfr _b_6986(.a(_w_8411),.q(_w_8412));
  bfr _b_6985(.a(_w_8410),.q(_w_8411));
  bfr _b_6981(.a(_w_8406),.q(_w_8407));
  bfr _b_6977(.a(_w_8402),.q(_w_8403));
  bfr _b_6975(.a(G72),.q(_w_8401));
  bfr _b_6974(.a(_w_8399),.q(_w_8366));
  bfr _b_7448(.a(_w_8873),.q(_w_8874));
  bfr _b_6973(.a(_w_8398),.q(_w_8399));
  bfr _b_6971(.a(_w_8396),.q(_w_8397));
  bfr _b_6968(.a(_w_8393),.q(_w_8394));
  bfr _b_6967(.a(_w_8392),.q(_w_8393));
  bfr _b_6964(.a(_w_8389),.q(_w_8390));
  bfr _b_6962(.a(_w_8387),.q(_w_8388));
  bfr _b_6961(.a(_w_8386),.q(_w_8387));
  bfr _b_6960(.a(_w_8385),.q(_w_8386));
  bfr _b_6959(.a(_w_8384),.q(_w_8385));
  bfr _b_6957(.a(_w_8382),.q(_w_8383));
  bfr _b_6955(.a(_w_8380),.q(_w_8381));
  bfr _b_6954(.a(_w_8379),.q(_w_8380));
  bfr _b_6950(.a(_w_8375),.q(_w_8376));
  bfr _b_7371(.a(_w_8796),.q(_w_8797));
  bfr _b_6949(.a(_w_8374),.q(_w_8375));
  bfr _b_6947(.a(_w_8372),.q(_w_8373));
  bfr _b_6946(.a(_w_8371),.q(_w_8372));
  bfr _b_6941(.a(G71),.q(_w_8367));
  bfr _b_6938(.a(_w_8363),.q(_w_8364));
  bfr _b_6936(.a(_w_8361),.q(_w_8362));
  bfr _b_6934(.a(_w_8359),.q(_w_8360));
  bfr _b_6933(.a(_w_8358),.q(_w_8359));
  bfr _b_6931(.a(_w_8356),.q(_w_8357));
  bfr _b_6927(.a(_w_8352),.q(_w_8353));
  bfr _b_6926(.a(_w_8351),.q(_w_8352));
  bfr _b_6925(.a(_w_8350),.q(_w_8351));
  bfr _b_6923(.a(_w_8348),.q(_w_8349));
  bfr _b_6922(.a(_w_8347),.q(_w_8348));
  bfr _b_6918(.a(_w_8343),.q(_w_8344));
  bfr _b_7123(.a(_w_8548),.q(_w_8549));
  bfr _b_6913(.a(_w_8338),.q(_w_8339));
  bfr _b_6911(.a(_w_8336),.q(_w_8337));
  bfr _b_6909(.a(_w_8334),.q(_w_8335));
  bfr _b_6908(.a(_w_8333),.q(_w_8334));
  bfr _b_6905(.a(G7),.q(_w_8331));
  bfr _b_6902(.a(_w_8327),.q(_w_8328));
  bfr _b_6900(.a(_w_8325),.q(_w_8326));
  bfr _b_6897(.a(_w_8322),.q(_w_8323));
  bfr _b_6895(.a(_w_8320),.q(_w_8321));
  bfr _b_6892(.a(_w_8317),.q(_w_8318));
  bfr _b_6891(.a(_w_8316),.q(_w_8317));
  bfr _b_6889(.a(_w_8314),.q(_w_8315));
  bfr _b_6882(.a(_w_8307),.q(_w_8308));
  bfr _b_6876(.a(_w_8301),.q(_w_8302));
  bfr _b_6875(.a(_w_8300),.q(_w_8301));
  bfr _b_6873(.a(_w_8298),.q(_w_8299));
  bfr _b_6870(.a(_w_8295),.q(_w_8262));
  bfr _b_6869(.a(_w_8294),.q(_w_8295));
  bfr _b_6868(.a(_w_8293),.q(_w_8294));
  bfr _b_6867(.a(_w_8292),.q(_w_8293));
  bfr _b_6866(.a(_w_8291),.q(_w_8292));
  bfr _b_6864(.a(_w_8289),.q(_w_8290));
  bfr _b_6863(.a(_w_8288),.q(_w_8289));
  bfr _b_6862(.a(_w_8287),.q(_w_8288));
  bfr _b_6861(.a(_w_8286),.q(_w_8287));
  bfr _b_6857(.a(_w_8282),.q(_w_8283));
  bfr _b_6854(.a(_w_8279),.q(_w_8280));
  bfr _b_6853(.a(_w_8278),.q(_w_8279));
  bfr _b_6852(.a(_w_8277),.q(_w_8278));
  bfr _b_6851(.a(_w_8276),.q(_w_8277));
  bfr _b_6850(.a(_w_8275),.q(_w_8276));
  bfr _b_6848(.a(_w_8273),.q(_w_8274));
  bfr _b_6847(.a(_w_8272),.q(_w_8273));
  bfr _b_6845(.a(_w_8270),.q(_w_8271));
  bfr _b_6841(.a(_w_8266),.q(_w_8267));
  bfr _b_6840(.a(_w_8265),.q(_w_8266));
  bfr _b_6839(.a(_w_8264),.q(_w_8265));
  bfr _b_6837(.a(G68),.q(_w_8263));
  bfr _b_7515(.a(_w_8940),.q(_w_8941));
  bfr _b_6836(.a(_w_8261),.q(_w_8224));
  bfr _b_6835(.a(_w_8260),.q(_w_8261));
  bfr _b_6834(.a(_w_8259),.q(_w_8260));
  bfr _b_6833(.a(_w_8258),.q(_w_8259));
  bfr _b_6831(.a(_w_8256),.q(_w_8257));
  bfr _b_6829(.a(_w_8254),.q(_w_8255));
  bfr _b_6826(.a(_w_8251),.q(_w_8252));
  bfr _b_6825(.a(_w_8250),.q(_w_8251));
  bfr _b_6820(.a(_w_8245),.q(_w_8246));
  bfr _b_6819(.a(_w_8244),.q(_w_8245));
  bfr _b_6817(.a(_w_8242),.q(_w_8243));
  bfr _b_6814(.a(_w_8239),.q(_w_8240));
  bfr _b_6813(.a(_w_8238),.q(_w_8239));
  bfr _b_6812(.a(_w_8237),.q(_w_8238));
  bfr _b_6810(.a(_w_8235),.q(_w_8236));
  bfr _b_6808(.a(_w_8233),.q(_w_8234));
  bfr _b_6807(.a(_w_8232),.q(_w_8233));
  bfr _b_6805(.a(_w_8230),.q(_w_8231));
  bfr _b_6803(.a(_w_8228),.q(_w_8229));
  bfr _b_7468(.a(_w_8893),.q(_w_8894));
  bfr _b_6802(.a(_w_8227),.q(_w_8228));
  bfr _b_6798(.a(_w_8223),.q(_w_8187));
  bfr _b_7079(.a(_w_8504),.q(_w_8505));
  bfr _b_6793(.a(_w_8218),.q(_w_8219));
  bfr _b_6791(.a(_w_8216),.q(_w_8217));
  bfr _b_6789(.a(_w_8214),.q(_w_8215));
  bfr _b_6788(.a(_w_8213),.q(_w_8214));
  bfr _b_6787(.a(_w_8212),.q(_w_8213));
  bfr _b_6786(.a(_w_8211),.q(_w_8212));
  bfr _b_6785(.a(_w_8210),.q(_w_8211));
  bfr _b_6784(.a(_w_8209),.q(_w_8210));
  bfr _b_7169(.a(_w_8594),.q(_w_8595));
  bfr _b_6783(.a(_w_8208),.q(_w_8209));
  bfr _b_6781(.a(_w_8206),.q(_w_8207));
  bfr _b_6777(.a(_w_8202),.q(_w_8203));
  bfr _b_6775(.a(_w_8200),.q(_w_8201));
  bfr _b_6774(.a(_w_8199),.q(_w_8200));
  bfr _b_6773(.a(_w_8198),.q(_w_8199));
  bfr _b_6772(.a(_w_8197),.q(_w_8198));
  bfr _b_6770(.a(_w_8195),.q(_w_8196));
  bfr _b_6767(.a(_w_8192),.q(_w_8193));
  bfr _b_6766(.a(_w_8191),.q(_w_8192));
  bfr _b_6764(.a(_w_8189),.q(_w_8190));
  bfr _b_6762(.a(G66),.q(_w_8188));
  bfr _b_6761(.a(_w_8186),.q(_w_8184));
  bfr _b_6760(.a(_w_8185),.q(_w_8186));
  bfr _b_7320(.a(_w_8745),.q(_w_8746));
  bfr _b_6759(.a(G65),.q(_w_8185));
  bfr _b_6753(.a(_w_8178),.q(_w_8179));
  bfr _b_6751(.a(_w_8176),.q(_w_8177));
  bfr _b_6750(.a(_w_8175),.q(_w_8176));
  bfr _b_6747(.a(_w_8172),.q(_w_8173));
  bfr _b_6746(.a(_w_8171),.q(_w_8172));
  bfr _b_6745(.a(_w_8170),.q(_w_8171));
  bfr _b_6743(.a(_w_8168),.q(_w_8169));
  bfr _b_6742(.a(_w_8167),.q(_w_8168));
  bfr _b_6741(.a(_w_8166),.q(_w_8167));
  bfr _b_6740(.a(_w_8165),.q(_w_8166));
  bfr _b_6737(.a(_w_8162),.q(_w_8163));
  bfr _b_6736(.a(_w_8161),.q(_w_8162));
  bfr _b_6734(.a(_w_8159),.q(_w_8160));
  bfr _b_6733(.a(_w_8158),.q(_w_8159));
  bfr _b_6732(.a(_w_8157),.q(_w_8158));
  bfr _b_6731(.a(_w_8156),.q(_w_8157));
  bfr _b_6729(.a(_w_8154),.q(_w_8155));
  bfr _b_6727(.a(_w_8152),.q(_w_8153));
  bfr _b_6726(.a(_w_8151),.q(_w_8152));
  bfr _b_6722(.a(G63),.q(_w_8147));
  bfr _b_6720(.a(_w_8145),.q(_w_8146));
  bfr _b_6719(.a(_w_8144),.q(_w_8145));
  bfr _b_6718(.a(_w_8143),.q(_w_8144));
  bfr _b_6717(.a(_w_8142),.q(_w_8143));
  bfr _b_6715(.a(_w_8140),.q(_w_8141));
  bfr _b_6714(.a(_w_8139),.q(_w_8140));
  bfr _b_7557(.a(_w_8982),.q(_w_8983));
  bfr _b_6713(.a(_w_8138),.q(_w_8139));
  bfr _b_6712(.a(_w_8137),.q(_w_8138));
  bfr _b_6711(.a(_w_8136),.q(_w_8137));
  bfr _b_6723(.a(G64),.q(_w_8149));
  bfr _b_6710(.a(_w_8135),.q(_w_8136));
  bfr _b_6706(.a(_w_8131),.q(_w_8132));
  bfr _b_6705(.a(_w_8130),.q(_w_8131));
  bfr _b_6701(.a(_w_8126),.q(_w_8127));
  bfr _b_6699(.a(_w_8124),.q(_w_8125));
  bfr _b_6697(.a(_w_8122),.q(_w_8123));
  bfr _b_6696(.a(_w_8121),.q(_w_8122));
  bfr _b_6695(.a(_w_8120),.q(_w_8121));
  bfr _b_6694(.a(_w_8119),.q(_w_8120));
  bfr _b_6693(.a(_w_8118),.q(_w_8119));
  bfr _b_6806(.a(_w_8231),.q(_w_8232));
  bfr _b_6689(.a(_w_8114),.q(_w_8115));
  bfr _b_6687(.a(_w_8112),.q(_w_8080));
  bfr _b_6686(.a(_w_8111),.q(_w_8112));
  bfr _b_6685(.a(_w_8110),.q(_w_8111));
  bfr _b_7298(.a(_w_8723),.q(_w_8724));
  bfr _b_6681(.a(_w_8106),.q(_w_8107));
  bfr _b_6680(.a(_w_8105),.q(_w_8106));
  bfr _b_6678(.a(_w_8103),.q(_w_8104));
  bfr _b_6676(.a(_w_8101),.q(_w_8102));
  bfr _b_6675(.a(_w_8100),.q(_w_8101));
  bfr _b_7324(.a(_w_8749),.q(_w_8750));
  bfr _b_6670(.a(_w_8095),.q(_w_8096));
  bfr _b_7501(.a(_w_8926),.q(_w_8927));
  bfr _b_6666(.a(_w_8091),.q(_w_8092));
  bfr _b_6661(.a(_w_8086),.q(_w_8087));
  bfr _b_6660(.a(_w_8085),.q(_w_8086));
  bfr _b_6659(.a(_w_8084),.q(_w_8085));
  bfr _b_6658(.a(_w_8083),.q(_w_8084));
  bfr _b_6656(.a(_w_8081),.q(_w_8082));
  bfr _b_6655(.a(G6),.q(_w_8081));
  bfr _b_6653(.a(_w_8078),.q(_w_8079));
  bfr _b_6651(.a(_w_8076),.q(_w_8077));
  bfr _b_6649(.a(_w_8074),.q(_w_8075));
  bfr _b_6648(.a(_w_8073),.q(_w_8074));
  bfr _b_6645(.a(_w_8070),.q(_w_8071));
  bfr _b_6642(.a(_w_8067),.q(_w_8068));
  bfr _b_6641(.a(_w_8066),.q(_w_8067));
  bfr _b_6640(.a(_w_8065),.q(_w_8066));
  bfr _b_6639(.a(_w_8064),.q(_w_8065));
  bfr _b_6888(.a(_w_8313),.q(_w_8314));
  bfr _b_6638(.a(_w_8063),.q(_w_8064));
  bfr _b_6637(.a(_w_8062),.q(_w_8063));
  bfr _b_6636(.a(_w_8061),.q(_w_8062));
  bfr _b_6634(.a(_w_8059),.q(_w_8060));
  bfr _b_6629(.a(_w_8054),.q(_w_8055));
  bfr _b_6628(.a(_w_8053),.q(_w_8054));
  bfr _b_6627(.a(_w_8052),.q(_w_8053));
  bfr _b_6626(.a(_w_8051),.q(_w_8052));
  bfr _b_6625(.a(_w_8050),.q(_w_8051));
  bfr _b_6623(.a(_w_8048),.q(_w_8049));
  bfr _b_6622(.a(_w_8047),.q(_w_8048));
  bfr _b_6621(.a(_w_8046),.q(_w_8047));
  bfr _b_6620(.a(_w_8045),.q(_w_8046));
  bfr _b_6619(.a(_w_8044),.q(_w_8045));
  bfr _b_6618(.a(_w_8043),.q(_w_8044));
  bfr _b_6778(.a(_w_8203),.q(_w_8204));
  bfr _b_6616(.a(_w_8041),.q(_w_8042));
  bfr _b_7305(.a(_w_8730),.q(_w_8731));
  bfr _b_6613(.a(_w_8038),.q(_w_8039));
  bfr _b_6611(.a(G58),.q(_w_8037));
  bfr _b_6610(.a(_w_8035),.q(_w_8015));
  bfr _b_6609(.a(_w_8034),.q(_w_8035));
  bfr _b_6608(.a(_w_8033),.q(_w_8034));
  bfr _b_6607(.a(_w_8032),.q(_w_8033));
  bfr _b_6979(.a(_w_8404),.q(_w_8405));
  bfr _b_6604(.a(_w_8029),.q(_w_8030));
  bfr _b_7370(.a(_w_8795),.q(_w_8796));
  bfr _b_6603(.a(_w_8028),.q(_w_8029));
  bfr _b_6600(.a(_w_8025),.q(_w_8026));
  bfr _b_6599(.a(_w_8024),.q(_w_8025));
  bfr _b_6598(.a(_w_8023),.q(_w_8024));
  bfr _b_6597(.a(_w_8022),.q(_w_8023));
  bfr _b_6596(.a(_w_8021),.q(_w_8022));
  bfr _b_6595(.a(_w_8020),.q(_w_8021));
  bfr _b_6592(.a(_w_8017),.q(_w_8018));
  bfr _b_6589(.a(_w_8014),.q(_w_7994));
  bfr _b_6928(.a(_w_8353),.q(_w_8354));
  bfr _b_6588(.a(_w_8013),.q(_w_8014));
  bfr _b_6583(.a(_w_8008),.q(_w_8009));
  bfr _b_7514(.a(_w_8939),.q(_w_8940));
  bfr _b_6582(.a(_w_8007),.q(_w_8008));
  bfr _b_6581(.a(_w_8006),.q(_w_8007));
  bfr _b_6579(.a(_w_8004),.q(_w_8005));
  bfr _b_6578(.a(_w_8003),.q(_w_8004));
  bfr _b_6576(.a(_w_8001),.q(_w_8002));
  bfr _b_6575(.a(_w_8000),.q(_w_8001));
  bfr _b_6574(.a(_w_7999),.q(_w_8000));
  bfr _b_6571(.a(_w_7996),.q(_w_7997));
  bfr _b_6566(.a(_w_7991),.q(_w_7992));
  bfr _b_6562(.a(_w_7987),.q(_w_7988));
  bfr _b_6593(.a(_w_8018),.q(_w_8019));
  bfr _b_6561(.a(_w_7986),.q(_w_7987));
  bfr _b_6560(.a(_w_7985),.q(_w_7986));
  bfr _b_6558(.a(_w_7983),.q(_w_7984));
  bfr _b_6556(.a(_w_7981),.q(_w_7982));
  bfr _b_6796(.a(_w_8221),.q(_w_8222));
  bfr _b_6554(.a(_w_7979),.q(_w_7980));
  bfr _b_6549(.a(_w_7974),.q(_w_7975));
  bfr _b_7464(.a(_w_8889),.q(_w_8890));
  bfr _b_6548(.a(G55),.q(_w_7974));
  bfr _b_6547(.a(_w_7972),.q(_w_7961));
  bfr _b_6546(.a(_w_7971),.q(_w_7972));
  bfr _b_6541(.a(_w_7966),.q(_w_7967));
  bfr _b_6539(.a(_w_7964),.q(_w_7965));
  bfr _b_6537(.a(_w_7962),.q(_w_7963));
  bfr _b_6536(.a(G54),.q(_w_7962));
  bfr _b_6535(.a(_w_7960),.q(_w_7939));
  bfr _b_6530(.a(_w_7955),.q(_w_7956));
  bfr _b_6529(.a(_w_7954),.q(_w_7955));
  bfr _b_6594(.a(_w_8019),.q(_w_8020));
  bfr _b_6528(.a(_w_7953),.q(_w_7954));
  bfr _b_6527(.a(_w_7952),.q(_w_7953));
  bfr _b_6526(.a(_w_7951),.q(_w_7952));
  bfr _b_6522(.a(_w_7947),.q(_w_7948));
  bfr _b_6521(.a(_w_7946),.q(_w_7947));
  bfr _b_6520(.a(_w_7945),.q(_w_7946));
  bfr _b_6519(.a(_w_7944),.q(_w_7945));
  bfr _b_6518(.a(_w_7943),.q(_w_7944));
  bfr _b_6516(.a(_w_7941),.q(_w_7942));
  bfr _b_6513(.a(_w_7938),.q(_w_7918));
  bfr _b_6511(.a(_w_7936),.q(_w_7937));
  bfr _b_6508(.a(_w_7933),.q(_w_7934));
  bfr _b_6506(.a(_w_7931),.q(_w_7932));
  bfr _b_6505(.a(_w_7930),.q(_w_7931));
  bfr _b_6503(.a(_w_7928),.q(_w_7929));
  bfr _b_6501(.a(_w_7926),.q(_w_7927));
  bfr _b_6500(.a(_w_7925),.q(_w_7926));
  bfr _b_7256(.a(_w_8681),.q(_w_8682));
  bfr _b_6885(.a(_w_8310),.q(_w_8311));
  bfr _b_6498(.a(_w_7923),.q(_w_7924));
  bfr _b_6496(.a(_w_7921),.q(_w_7922));
  bfr _b_6494(.a(_w_7919),.q(_w_7920));
  bfr _b_6493(.a(G52),.q(_w_7919));
  bfr _b_6492(.a(_w_7917),.q(_w_7897));
  bfr _b_6491(.a(_w_7916),.q(_w_7917));
  bfr _b_6490(.a(_w_7915),.q(_w_7916));
  bfr _b_6488(.a(_w_7913),.q(_w_7914));
  bfr _b_6485(.a(_w_7910),.q(_w_7911));
  bfr _b_6484(.a(_w_7909),.q(_w_7910));
  bfr _b_6482(.a(_w_7907),.q(_w_7908));
  bfr _b_6481(.a(_w_7906),.q(_w_7907));
  bfr _b_6477(.a(_w_7902),.q(_w_7903));
  bfr _b_6474(.a(_w_7899),.q(_w_7900));
  bfr _b_6473(.a(_w_7898),.q(_w_7899));
  bfr _b_7274(.a(_w_8699),.q(_w_8700));
  bfr _b_6471(.a(_w_7896),.q(_w_7875));
  bfr _b_6470(.a(_w_7895),.q(_w_7896));
  bfr _b_6469(.a(_w_7894),.q(_w_7895));
  bfr _b_6468(.a(_w_7893),.q(_w_7894));
  bfr _b_6466(.a(_w_7891),.q(_w_7892));
  bfr _b_6463(.a(_w_7888),.q(_w_7889));
  bfr _b_6502(.a(_w_7927),.q(_w_7928));
  bfr _b_6462(.a(_w_7887),.q(_w_7888));
  bfr _b_6461(.a(_w_7886),.q(_w_7887));
  bfr _b_6460(.a(_w_7885),.q(_w_7886));
  bfr _b_7311(.a(_w_8736),.q(_w_8737));
  bfr _b_6459(.a(_w_7884),.q(_w_7885));
  bfr _b_6458(.a(_w_7883),.q(_w_7884));
  bfr _b_6457(.a(_w_7882),.q(_w_7883));
  bfr _b_6456(.a(_w_7881),.q(_w_7882));
  bfr _b_6453(.a(_w_7878),.q(_w_7879));
  bfr _b_6452(.a(_w_7877),.q(_w_7878));
  bfr _b_6451(.a(_w_7876),.q(_w_7877));
  bfr _b_6450(.a(G50),.q(_w_7876));
  bfr _b_6449(.a(_w_7874),.q(_w_7842));
  bfr _b_6448(.a(_w_7873),.q(_w_7874));
  bfr _b_6446(.a(_w_7871),.q(_w_7872));
  bfr _b_6444(.a(_w_7869),.q(_w_7870));
  bfr _b_6443(.a(_w_7868),.q(_w_7869));
  bfr _b_6441(.a(_w_7866),.q(_w_7867));
  bfr _b_6440(.a(_w_7865),.q(_w_7866));
  bfr _b_6437(.a(_w_7862),.q(_w_7863));
  bfr _b_6887(.a(_w_8312),.q(_w_8313));
  bfr _b_6436(.a(_w_7861),.q(_w_7862));
  bfr _b_6434(.a(_w_7859),.q(_w_7860));
  bfr _b_7467(.a(_w_8892),.q(_w_8893));
  bfr _b_6472(.a(G51),.q(_w_7898));
  bfr _b_6432(.a(_w_7857),.q(_w_7858));
  bfr _b_6428(.a(_w_7853),.q(_w_7854));
  bfr _b_6427(.a(_w_7852),.q(_w_7853));
  bfr _b_6423(.a(_w_7848),.q(_w_7849));
  bfr _b_6422(.a(_w_7847),.q(_w_7848));
  bfr _b_6421(.a(_w_7846),.q(_w_7847));
  bfr _b_6419(.a(_w_7844),.q(_w_7845));
  bfr _b_7022(.a(_w_8447),.q(_w_8448));
  bfr _b_6417(.a(G5),.q(_w_7843));
  bfr _b_6415(.a(_w_7840),.q(_w_7841));
  bfr _b_6414(.a(_w_7839),.q(_w_7840));
  bfr _b_6413(.a(_w_7838),.q(_w_7839));
  bfr _b_7502(.a(_w_8927),.q(_w_8928));
  bfr _b_6412(.a(_w_7837),.q(_w_7838));
  bfr _b_6410(.a(_w_7835),.q(_w_7836));
  bfr _b_6407(.a(_w_7832),.q(_w_7833));
  bfr _b_6404(.a(_w_7829),.q(_w_7830));
  bfr _b_6402(.a(_w_7827),.q(_w_7828));
  bfr _b_6401(.a(_w_7826),.q(_w_7827));
  bfr _b_6400(.a(_w_7825),.q(_w_7826));
  bfr _b_6396(.a(G49),.q(_w_7822));
  bfr _b_6393(.a(_w_7818),.q(_w_7819));
  bfr _b_6391(.a(_w_7816),.q(_w_7817));
  bfr _b_6388(.a(_w_7813),.q(_w_7814));
  bfr _b_6387(.a(_w_7812),.q(_w_7813));
  bfr _b_6386(.a(_w_7811),.q(_w_7812));
  bfr _b_6385(.a(_w_7810),.q(_w_7811));
  bfr _b_6384(.a(_w_7809),.q(_w_7810));
  bfr _b_6381(.a(_w_7806),.q(_w_7807));
  bfr _b_6380(.a(_w_7805),.q(_w_7806));
  bfr _b_6379(.a(_w_7804),.q(_w_7805));
  bfr _b_6378(.a(_w_7803),.q(_w_7804));
  bfr _b_6377(.a(_w_7802),.q(_w_7803));
  bfr _b_6374(.a(G48),.q(_w_7800));
  bfr _b_6373(.a(_w_7798),.q(_w_7778));
  bfr _b_6372(.a(_w_7797),.q(_w_7798));
  bfr _b_6370(.a(_w_7795),.q(_w_7796));
  bfr _b_6367(.a(_w_7792),.q(_w_7793));
  bfr _b_7336(.a(_w_8761),.q(_w_8762));
  bfr _b_6366(.a(_w_7791),.q(_w_7792));
  bfr _b_6364(.a(_w_7789),.q(_w_7790));
  bfr _b_6361(.a(_w_7786),.q(_w_7787));
  bfr _b_6744(.a(_w_8169),.q(_w_8170));
  bfr _b_6359(.a(_w_7784),.q(_w_7785));
  bfr _b_6358(.a(_w_7783),.q(_w_7784));
  bfr _b_6357(.a(_w_7782),.q(_w_7783));
  bfr _b_6356(.a(_w_7781),.q(_w_7782));
  bfr _b_6353(.a(G47),.q(_w_7779));
  bfr _b_6352(.a(_w_7777),.q(_w_7757));
  bfr _b_6351(.a(_w_7776),.q(_w_7777));
  bfr _b_6350(.a(_w_7775),.q(_w_7776));
  bfr _b_6348(.a(_w_7773),.q(_w_7774));
  bfr _b_6346(.a(_w_7771),.q(_w_7772));
  bfr _b_6345(.a(_w_7770),.q(_w_7771));
  bfr _b_6339(.a(_w_7764),.q(_w_7765));
  bfr _b_6338(.a(_w_7763),.q(_w_7764));
  bfr _b_6335(.a(_w_7760),.q(_w_7761));
  bfr _b_6333(.a(_w_7758),.q(_w_7759));
  bfr _b_6332(.a(G46),.q(_w_7758));
  bfr _b_6331(.a(_w_7756),.q(_w_7736));
  bfr _b_6330(.a(_w_7755),.q(_w_7756));
  bfr _b_7197(.a(_w_8622),.q(_w_8623));
  bfr _b_6329(.a(_w_7754),.q(_w_7755));
  bfr _b_6480(.a(_w_7905),.q(_w_7906));
  bfr _b_6328(.a(_w_7753),.q(_w_7754));
  bfr _b_6327(.a(_w_7752),.q(_w_7753));
  bfr _b_6325(.a(_w_7750),.q(_w_7751));
  bfr _b_7146(.a(_w_8571),.q(_w_8572));
  bfr _b_6324(.a(_w_7749),.q(_w_7750));
  bfr _b_6322(.a(_w_7747),.q(_w_7748));
  bfr _b_6318(.a(_w_7743),.q(_w_7744));
  bfr _b_6943(.a(_w_8368),.q(_w_8369));
  bfr _b_6317(.a(_w_7742),.q(_w_7743));
  bfr _b_6315(.a(_w_7740),.q(_w_7741));
  bfr _b_6312(.a(_w_7737),.q(_w_7738));
  bfr _b_6311(.a(G45),.q(_w_7737));
  bfr _b_6550(.a(_w_7975),.q(_w_7976));
  bfr _b_6310(.a(_w_7735),.q(_w_7715));
  bfr _b_6823(.a(_w_8248),.q(_w_8249));
  bfr _b_6309(.a(_w_7734),.q(_w_7735));
  bfr _b_6307(.a(_w_7732),.q(_w_7733));
  bfr _b_6827(.a(_w_8252),.q(_w_8253));
  bfr _b_6304(.a(_w_7729),.q(_w_7730));
  bfr _b_6303(.a(_w_7728),.q(_w_7729));
  bfr _b_6301(.a(_w_7726),.q(_w_7727));
  bfr _b_6299(.a(_w_7724),.q(_w_7725));
  bfr _b_6298(.a(_w_7723),.q(_w_7724));
  bfr _b_6297(.a(_w_7722),.q(_w_7723));
  bfr _b_6295(.a(_w_7720),.q(_w_7721));
  bfr _b_6292(.a(_w_7717),.q(_w_7718));
  bfr _b_6290(.a(G44),.q(_w_7716));
  bfr _b_6289(.a(_w_7714),.q(_w_7694));
  bfr _b_6285(.a(_w_7710),.q(_w_7711));
  bfr _b_6284(.a(_w_7709),.q(_w_7710));
  bfr _b_6283(.a(_w_7708),.q(_w_7709));
  bfr _b_6282(.a(_w_7707),.q(_w_7708));
  bfr _b_6279(.a(_w_7704),.q(_w_7705));
  bfr _b_6278(.a(_w_7703),.q(_w_7704));
  bfr _b_6277(.a(_w_7702),.q(_w_7703));
  bfr _b_6274(.a(_w_7699),.q(_w_7700));
  bfr _b_6273(.a(_w_7698),.q(_w_7699));
  bfr _b_6272(.a(_w_7697),.q(_w_7698));
  bfr _b_6270(.a(_w_7695),.q(_w_7696));
  bfr _b_6268(.a(_w_7693),.q(_w_7661));
  bfr _b_6267(.a(_w_7692),.q(_w_7693));
  bfr _b_6263(.a(_w_7688),.q(_w_7689));
  bfr _b_6792(.a(_w_8217),.q(_w_8218));
  bfr _b_6262(.a(_w_7687),.q(_w_7688));
  bfr _b_7140(.a(_w_8565),.q(_w_8566));
  bfr _b_6260(.a(_w_7685),.q(_w_7686));
  bfr _b_6257(.a(_w_7682),.q(_w_7683));
  bfr _b_6255(.a(_w_7680),.q(_w_7681));
  bfr _b_6254(.a(_w_7679),.q(_w_7680));
  bfr _b_6251(.a(_w_7676),.q(_w_7677));
  bfr _b_6250(.a(_w_7675),.q(_w_7676));
  bfr _b_6249(.a(_w_7674),.q(_w_7675));
  bfr _b_6248(.a(_w_7673),.q(_w_7674));
  bfr _b_6244(.a(_w_7669),.q(_w_7670));
  bfr _b_6241(.a(_w_7666),.q(_w_7667));
  bfr _b_6240(.a(_w_7665),.q(_w_7666));
  bfr _b_7483(.a(G87),.q(_w_8909));
  bfr _b_6239(.a(_w_7664),.q(_w_7665));
  bfr _b_6483(.a(_w_7908),.q(_w_7909));
  bfr _b_6238(.a(_w_7663),.q(_w_7664));
  bfr _b_6231(.a(_w_7656),.q(_w_7657));
  bfr _b_6230(.a(_w_7655),.q(_w_7656));
  bfr _b_6228(.a(_w_7653),.q(_w_7654));
  bfr _b_6227(.a(_w_7652),.q(_w_7653));
  bfr _b_6226(.a(_w_7651),.q(_w_7652));
  bfr _b_6224(.a(_w_7649),.q(_w_7650));
  bfr _b_6223(.a(_w_7648),.q(_w_7649));
  bfr _b_6222(.a(_w_7647),.q(_w_7648));
  bfr _b_6219(.a(_w_7644),.q(_w_7645));
  bfr _b_6217(.a(_w_7642),.q(_w_7643));
  bfr _b_6214(.a(_w_7639),.q(_w_7640));
  bfr _b_6207(.a(_w_7632),.q(_w_7633));
  bfr _b_6206(.a(_w_7631),.q(_w_7632));
  bfr _b_6205(.a(_w_7630),.q(_w_7631));
  bfr _b_6204(.a(_w_7629),.q(_w_7630));
  bfr _b_7152(.a(_w_8577),.q(_w_8578));
  bfr _b_6203(.a(G41),.q(_w_7629));
  bfr _b_6202(.a(_w_7627),.q(_w_7595));
  bfr _b_6201(.a(_w_7626),.q(_w_7627));
  bfr _b_6199(.a(_w_7624),.q(_w_7625));
  bfr _b_6197(.a(_w_7622),.q(_w_7623));
  bfr _b_6195(.a(_w_7620),.q(_w_7621));
  bfr _b_6194(.a(_w_7619),.q(_w_7620));
  bfr _b_6193(.a(_w_7618),.q(_w_7619));
  bfr _b_6191(.a(_w_7616),.q(_w_7617));
  bfr _b_6190(.a(_w_7615),.q(_w_7616));
  bfr _b_6189(.a(_w_7614),.q(_w_7615));
  bfr _b_6188(.a(_w_7613),.q(_w_7614));
  bfr _b_6183(.a(_w_7608),.q(_w_7609));
  bfr _b_6182(.a(_w_7607),.q(_w_7608));
  bfr _b_6180(.a(_w_7605),.q(_w_7606));
  bfr _b_6178(.a(_w_7603),.q(_w_7604));
  bfr _b_6725(.a(_w_8150),.q(_w_8151));
  bfr _b_6172(.a(_w_7597),.q(_w_7598));
  bfr _b_6171(.a(_w_7596),.q(_w_7597));
  bfr _b_6170(.a(G40),.q(_w_7596));
  bfr _b_7203(.a(_w_8628),.q(_w_8629));
  bfr _b_6169(.a(_w_7594),.q(_w_7562));
  bfr _b_6165(.a(_w_7590),.q(_w_7591));
  bfr _b_6162(.a(_w_7587),.q(_w_7588));
  bfr _b_6161(.a(_w_7586),.q(_w_7587));
  bfr _b_6160(.a(_w_7585),.q(_w_7586));
  bfr _b_6159(.a(_w_7584),.q(_w_7585));
  bfr _b_6531(.a(_w_7956),.q(_w_7957));
  bfr _b_6158(.a(_w_7583),.q(_w_7584));
  bfr _b_6153(.a(_w_7578),.q(_w_7579));
  bfr _b_6152(.a(_w_7577),.q(_w_7578));
  bfr _b_6151(.a(_w_7576),.q(_w_7577));
  bfr _b_6150(.a(_w_7575),.q(_w_7576));
  bfr _b_6147(.a(_w_7572),.q(_w_7573));
  bfr _b_6145(.a(_w_7570),.q(_w_7571));
  bfr _b_6144(.a(_w_7569),.q(_w_7570));
  bfr _b_6143(.a(_w_7568),.q(_w_7569));
  bfr _b_6141(.a(_w_7566),.q(_w_7567));
  bfr _b_6135(.a(_w_7560),.q(_w_7561));
  bfr _b_6133(.a(_w_7558),.q(_w_7559));
  bfr _b_6132(.a(_w_7557),.q(_w_7558));
  bfr _b_6128(.a(_w_7553),.q(_w_7554));
  bfr _b_6126(.a(_w_7551),.q(_w_7552));
  bfr _b_6124(.a(_w_7549),.q(_w_7550));
  bfr _b_6123(.a(_w_7548),.q(_w_7549));
  bfr _b_7281(.a(G81),.q(_w_8707));
  bfr _b_6122(.a(_w_7547),.q(_w_7548));
  bfr _b_6121(.a(_w_7546),.q(_w_7547));
  bfr _b_7480(.a(_w_8905),.q(_w_8906));
  bfr _b_6120(.a(_w_7545),.q(_w_7546));
  bfr _b_6115(.a(_w_7540),.q(_w_7541));
  bfr _b_6112(.a(_w_7537),.q(_w_7538));
  bfr _b_6111(.a(_w_7536),.q(_w_7537));
  bfr _b_6569(.a(G56),.q(_w_7995));
  bfr _b_6110(.a(_w_7535),.q(_w_7536));
  bfr _b_7430(.a(_w_8855),.q(_w_8856));
  bfr _b_6108(.a(_w_7533),.q(_w_7534));
  bfr _b_6107(.a(_w_7532),.q(_w_7533));
  bfr _b_6103(.a(_w_7528),.q(_w_7510));
  bfr _b_6102(.a(_w_7527),.q(_w_7528));
  bfr _b_6101(.a(_w_7526),.q(_w_7527));
  bfr _b_7318(.a(_w_8743),.q(_w_8744));
  bfr _b_6100(.a(_w_7525),.q(_w_7526));
  bfr _b_6097(.a(_w_7522),.q(_w_7523));
  bfr _b_6092(.a(_w_7517),.q(_w_7518));
  bfr _b_6090(.a(_w_7515),.q(_w_7516));
  bfr _b_6086(.a(_w_7511),.q(_w_7512));
  bfr _b_6085(.a(G38),.q(_w_7511));
  bfr _b_6083(.a(_w_7508),.q(_w_7509));
  bfr _b_6081(.a(_w_7506),.q(_w_7507));
  bfr _b_6080(.a(_w_7505),.q(_w_7506));
  bfr _b_6078(.a(_w_7503),.q(_w_7504));
  bfr _b_6076(.a(_w_7501),.q(_w_7502));
  bfr _b_6075(.a(_w_7500),.q(_w_7501));
  bfr _b_6074(.a(_w_7499),.q(_w_7500));
  bfr _b_6073(.a(_w_7498),.q(_w_7499));
  bfr _b_6072(.a(_w_7497),.q(_w_7498));
  bfr _b_6070(.a(_w_7495),.q(_w_7496));
  bfr _b_6069(.a(_w_7494),.q(_w_7495));
  bfr _b_6068(.a(_w_7493),.q(_w_7494));
  bfr _b_6067(.a(_w_7492),.q(_w_7493));
  bfr _b_6065(.a(_w_7490),.q(_w_7458));
  bfr _b_6064(.a(_w_7489),.q(_w_7490));
  bfr _b_6063(.a(_w_7488),.q(_w_7489));
  bfr _b_6061(.a(_w_7486),.q(_w_7487));
  bfr _b_6059(.a(_w_7484),.q(_w_7485));
  bfr _b_6058(.a(_w_7483),.q(_w_7484));
  bfr _b_6055(.a(_w_7480),.q(_w_7481));
  bfr _b_6054(.a(_w_7479),.q(_w_7480));
  bfr _b_6053(.a(_w_7478),.q(_w_7479));
  bfr _b_6052(.a(_w_7477),.q(_w_7478));
  bfr _b_6047(.a(_w_7472),.q(_w_7473));
  bfr _b_6703(.a(_w_8128),.q(_w_8129));
  bfr _b_6045(.a(_w_7470),.q(_w_7471));
  bfr _b_6044(.a(_w_7469),.q(_w_7470));
  bfr _b_6043(.a(_w_7468),.q(_w_7469));
  bfr _b_6042(.a(_w_7467),.q(_w_7468));
  bfr _b_6040(.a(_w_7465),.q(_w_7466));
  bfr _b_6039(.a(_w_7464),.q(_w_7465));
  bfr _b_6038(.a(_w_7463),.q(_w_7464));
  bfr _b_6037(.a(_w_7462),.q(_w_7463));
  bfr _b_7532(.a(_w_8957),.q(_w_8958));
  bfr _b_6036(.a(_w_7461),.q(_w_7462));
  bfr _b_6035(.a(_w_7460),.q(_w_7461));
  bfr _b_6033(.a(G36),.q(_w_7459));
  bfr _b_6031(.a(G35),.q(_w_7457));
  bfr _b_6030(.a(G34),.q(_w_7455));
  bfr _b_6027(.a(_w_7452),.q(_w_7449));
  bfr _b_6025(.a(_w_7450),.q(_w_7451));
  bfr _b_6024(.a(G32),.q(_w_7450));
  bfr _b_6019(.a(_w_7444),.q(_w_7413));
  bfr _b_6015(.a(_w_7440),.q(_w_7441));
  bfr _b_6013(.a(_w_7438),.q(_w_7439));
  bfr _b_6008(.a(_w_7433),.q(_w_7434));
  bfr _b_6006(.a(_w_7431),.q(_w_7432));
  bfr _b_6005(.a(_w_7430),.q(_w_7431));
  bfr _b_6003(.a(_w_7428),.q(_w_7429));
  bfr _b_6002(.a(_w_7427),.q(_w_7428));
  bfr _b_6001(.a(_w_7426),.q(_w_7427));
  bfr _b_5998(.a(_w_7423),.q(_w_7424));
  bfr _b_5996(.a(_w_7421),.q(_w_7422));
  bfr _b_6014(.a(_w_7439),.q(_w_7440));
  bfr _b_5995(.a(_w_7420),.q(_w_7421));
  bfr _b_5994(.a(_w_7419),.q(_w_7420));
  bfr _b_7541(.a(_w_8966),.q(_w_8967));
  bfr _b_5993(.a(_w_7418),.q(_w_7419));
  bfr _b_5991(.a(_w_7416),.q(_w_7417));
  bfr _b_5989(.a(_w_7414),.q(_w_7415));
  bfr _b_5988(.a(G3),.q(_w_7414));
  bfr _b_5986(.a(G29),.q(_w_7412));
  bfr _b_5983(.a(_w_7408),.q(_w_7376));
  bfr _b_5982(.a(_w_7407),.q(_w_7408));
  bfr _b_5980(.a(_w_7405),.q(_w_7406));
  bfr _b_5978(.a(_w_7403),.q(_w_7404));
  bfr _b_5977(.a(_w_7402),.q(_w_7403));
  bfr _b_5976(.a(_w_7401),.q(_w_7402));
  bfr _b_5974(.a(_w_7399),.q(_w_7400));
  bfr _b_5970(.a(_w_7395),.q(_w_7396));
  bfr _b_5969(.a(_w_7394),.q(_w_7395));
  bfr _b_5968(.a(_w_7393),.q(_w_7394));
  bfr _b_5967(.a(_w_7392),.q(_w_7393));
  bfr _b_5965(.a(_w_7390),.q(_w_7391));
  bfr _b_5962(.a(_w_7387),.q(_w_7388));
  bfr _b_5961(.a(_w_7386),.q(_w_7387));
  bfr _b_5958(.a(_w_7383),.q(_w_7384));
  bfr _b_5957(.a(_w_7382),.q(_w_7383));
  bfr _b_5955(.a(_w_7380),.q(_w_7381));
  bfr _b_5952(.a(_w_7377),.q(_w_7378));
  bfr _b_5948(.a(_w_7373),.q(_w_7374));
  bfr _b_5946(.a(_w_7371),.q(_w_7372));
  bfr _b_7081(.a(_w_8506),.q(_w_8507));
  bfr _b_5945(.a(_w_7370),.q(_w_7371));
  bfr _b_5944(.a(_w_7369),.q(_w_7370));
  bfr _b_5943(.a(_w_7368),.q(_w_7369));
  bfr _b_5940(.a(_w_7365),.q(_w_7366));
  bfr _b_5939(.a(_w_7364),.q(_w_7365));
  bfr _b_6568(.a(_w_7993),.q(_w_7973));
  bfr _b_5937(.a(_w_7362),.q(_w_7363));
  bfr _b_5936(.a(_w_7361),.q(_w_7362));
  bfr _b_5931(.a(_w_7356),.q(_w_7357));
  bfr _b_5929(.a(_w_7354),.q(_w_7355));
  bfr _b_5925(.a(_w_7350),.q(_w_7351));
  bfr _b_6586(.a(_w_8011),.q(_w_8012));
  bfr _b_5921(.a(_w_7346),.q(_w_7347));
  bfr _b_5917(.a(_w_7342),.q(_w_7310));
  bfr _b_5915(.a(_w_7340),.q(_w_7341));
  bfr _b_6821(.a(_w_8246),.q(_w_8247));
  bfr _b_5913(.a(_w_7338),.q(_w_7339));
  bfr _b_5912(.a(_w_7337),.q(_w_7338));
  bfr _b_7419(.a(_w_8844),.q(_w_8845));
  bfr _b_5909(.a(_w_7334),.q(_w_7335));
  bfr _b_5907(.a(_w_7332),.q(_w_7333));
  bfr _b_5964(.a(_w_7389),.q(_w_7390));
  bfr _b_5906(.a(_w_7331),.q(_w_7332));
  bfr _b_5905(.a(_w_7330),.q(_w_7331));
  bfr _b_5904(.a(_w_7329),.q(_w_7330));
  bfr _b_5903(.a(_w_7328),.q(_w_7329));
  bfr _b_5902(.a(_w_7327),.q(_w_7328));
  bfr _b_5901(.a(_w_7326),.q(_w_7327));
  bfr _b_5900(.a(_w_7325),.q(_w_7326));
  bfr _b_5899(.a(_w_7324),.q(_w_7325));
  bfr _b_5898(.a(_w_7323),.q(_w_7324));
  bfr _b_5896(.a(_w_7321),.q(_w_7322));
  bfr _b_5895(.a(_w_7320),.q(_w_7321));
  bfr _b_5894(.a(_w_7319),.q(_w_7320));
  bfr _b_6756(.a(_w_8181),.q(_w_8182));
  bfr _b_5893(.a(_w_7318),.q(_w_7319));
  bfr _b_5892(.a(_w_7317),.q(_w_7318));
  bfr _b_5890(.a(_w_7315),.q(_w_7316));
  bfr _b_5889(.a(_w_7314),.q(_w_7315));
  bfr _b_5888(.a(_w_7313),.q(_w_7314));
  bfr _b_5886(.a(_w_7311),.q(_w_7312));
  bfr _b_5884(.a(_w_7309),.q(_w_7277));
  bfr _b_5881(.a(_w_7306),.q(_w_7307));
  bfr _b_7202(.a(_w_8627),.q(_w_8628));
  bfr _b_5876(.a(_w_7301),.q(_w_7302));
  bfr _b_6192(.a(_w_7617),.q(_w_7618));
  bfr _b_5872(.a(_w_7297),.q(_w_7298));
  bfr _b_5866(.a(_w_7291),.q(_w_7292));
  bfr _b_6157(.a(_w_7582),.q(_w_7583));
  bfr _b_5865(.a(_w_7290),.q(_w_7291));
  bfr _b_5861(.a(_w_7286),.q(_w_7287));
  bfr _b_5860(.a(_w_7285),.q(_w_7286));
  bfr _b_5859(.a(_w_7284),.q(_w_7285));
  bfr _b_5857(.a(_w_7282),.q(_w_7283));
  bfr _b_5855(.a(_w_7280),.q(_w_7281));
  bfr _b_5853(.a(_w_7278),.q(_w_7279));
  bfr _b_5848(.a(_w_7273),.q(_w_7274));
  bfr _b_5845(.a(_w_7270),.q(_w_7271));
  bfr _b_5843(.a(_w_7268),.q(_w_7269));
  bfr _b_5840(.a(_w_7265),.q(_w_7266));
  bfr _b_5839(.a(_w_7264),.q(_w_7265));
  bfr _b_5838(.a(_w_7263),.q(_w_7264));
  bfr _b_5835(.a(_w_7260),.q(_w_7261));
  bfr _b_5942(.a(_w_7367),.q(_w_7368));
  bfr _b_5834(.a(_w_7259),.q(_w_7260));
  bfr _b_5832(.a(_w_7257),.q(_w_7258));
  bfr _b_7337(.a(_w_8762),.q(_w_8763));
  bfr _b_5831(.a(_w_7256),.q(_w_7257));
  bfr _b_5830(.a(_w_7255),.q(_w_7256));
  bfr _b_5828(.a(_w_7253),.q(_w_7254));
  bfr _b_5827(.a(_w_7252),.q(_w_7253));
  bfr _b_5824(.a(_w_7249),.q(_w_7250));
  bfr _b_5823(.a(_w_7248),.q(_w_7249));
  bfr _b_5821(.a(_w_7246),.q(_w_7247));
  bfr _b_5820(.a(_w_7245),.q(_w_7246));
  bfr _b_5819(.a(G23),.q(_w_7245));
  bfr _b_5818(.a(_w_7243),.q(_w_7212));
  bfr _b_5816(.a(_w_7241),.q(_w_7242));
  bfr _b_5815(.a(_w_7240),.q(_w_7241));
  bfr _b_5813(.a(_w_7238),.q(_w_7239));
  bfr _b_5812(.a(_w_7237),.q(_w_7238));
  bfr _b_5811(.a(_w_7236),.q(_w_7237));
  bfr _b_5810(.a(_w_7235),.q(_w_7236));
  bfr _b_5808(.a(_w_7233),.q(_w_7234));
  bfr _b_5807(.a(_w_7232),.q(_w_7233));
  bfr _b_5804(.a(_w_7229),.q(_w_7230));
  bfr _b_5802(.a(_w_7227),.q(_w_7228));
  bfr _b_5801(.a(_w_7226),.q(_w_7227));
  bfr _b_5799(.a(_w_7224),.q(_w_7225));
  bfr _b_5798(.a(_w_7223),.q(_w_7224));
  bfr _b_5973(.a(_w_7398),.q(_w_7399));
  bfr _b_5796(.a(_w_7221),.q(_w_7222));
  bfr _b_5792(.a(_w_7217),.q(_w_7218));
  bfr _b_5790(.a(_w_7215),.q(_w_7216));
  bfr _b_6797(.a(_w_8222),.q(_w_8223));
  bfr _b_5789(.a(_w_7214),.q(_w_7215));
  bfr _b_5786(.a(_w_7211),.q(_w_7205));
  bfr _b_7029(.a(_w_8454),.q(_w_8455));
  bfr _b_5785(.a(_w_7210),.q(_w_7211));
  bfr _b_5784(.a(_w_7209),.q(_w_7210));
  bfr _b_5783(.a(_w_7208),.q(_w_7209));
  bfr _b_5782(.a(_w_7207),.q(_w_7208));
  bfr _b_6344(.a(_w_7769),.q(_w_7770));
  bfr _b_5780(.a(G21),.q(_w_7206));
  bfr _b_5779(.a(_w_7204),.q(_w_7184));
  bfr _b_5778(.a(_w_7203),.q(_w_7204));
  bfr _b_5772(.a(_w_7197),.q(_w_7198));
  bfr _b_5771(.a(_w_7196),.q(_w_7197));
  bfr _b_6431(.a(_w_7856),.q(_w_7857));
  bfr _b_5769(.a(_w_7194),.q(_w_7195));
  bfr _b_6486(.a(_w_7911),.q(_w_7912));
  bfr _b_5767(.a(_w_7192),.q(_w_7193));
  bfr _b_5766(.a(_w_7191),.q(_w_7192));
  bfr _b_5765(.a(_w_7190),.q(_w_7191));
  bfr _b_5758(.a(_w_7183),.q(_w_7175));
  bfr _b_5757(.a(_w_7182),.q(_w_7183));
  bfr _b_5756(.a(_w_7181),.q(_w_7182));
  bfr _b_5755(.a(_w_7180),.q(_w_7181));
  bfr _b_5754(.a(_w_7179),.q(_w_7180));
  bfr _b_5753(.a(_w_7178),.q(_w_7179));
  bfr _b_5752(.a(_w_7177),.q(_w_7178));
  bfr _b_5747(.a(_w_7172),.q(_w_7173));
  bfr _b_5742(.a(_w_7167),.q(_w_7168));
  bfr _b_5737(.a(_w_7162),.q(_w_7163));
  bfr _b_5734(.a(_w_7159),.q(_w_7160));
  bfr _b_5733(.a(_w_7158),.q(_w_7159));
  bfr _b_5731(.a(_w_7156),.q(_w_7157));
  bfr _b_6119(.a(_w_7544),.q(_w_7545));
  bfr _b_5730(.a(_w_7155),.q(_w_7156));
  bfr _b_5724(.a(_w_7149),.q(_w_7150));
  bfr _b_5880(.a(_w_7305),.q(_w_7306));
  bfr _b_5723(.a(_w_7148),.q(_w_7149));
  bfr _b_5721(.a(_w_7146),.q(_w_7147));
  bfr _b_5719(.a(_w_7144),.q(_w_7145));
  bfr _b_5718(.a(_w_7143),.q(_w_7144));
  bfr _b_5717(.a(_w_7142),.q(_w_7143));
  bfr _b_5715(.a(_w_7140),.q(_w_7141));
  bfr _b_5714(.a(_w_7139),.q(_w_7140));
  bfr _b_5713(.a(_w_7138),.q(_w_7139));
  bfr _b_5711(.a(_w_7136),.q(_w_7137));
  bfr _b_5710(.a(_w_7135),.q(_w_7136));
  bfr _b_5707(.a(_w_7132),.q(_w_7133));
  bfr _b_5704(.a(_w_7129),.q(_w_7130));
  bfr _b_5703(.a(_w_7128),.q(_w_7129));
  bfr _b_5919(.a(_w_7344),.q(_w_7345));
  bfr _b_5702(.a(_w_7127),.q(_w_7128));
  bfr _b_7040(.a(_w_8465),.q(_w_8466));
  bfr _b_6545(.a(_w_7970),.q(_w_7971));
  bfr _b_5701(.a(_w_7126),.q(_w_7127));
  bfr _b_5697(.a(_w_7122),.q(_w_7123));
  bfr _b_5695(.a(G18),.q(_w_7121));
  bfr _b_5693(.a(_w_7118),.q(_w_7119));
  bfr _b_5692(.a(_w_7117),.q(_w_7118));
  bfr _b_5691(.a(_w_7116),.q(_w_7117));
  bfr _b_5689(.a(_w_7114),.q(_w_7115));
  bfr _b_5688(.a(_w_7113),.q(_w_7114));
  bfr _b_5685(.a(_w_7110),.q(_w_7111));
  bfr _b_7178(.a(G78),.q(_w_8604));
  bfr _b_5683(.a(_w_7108),.q(_w_7109));
  bfr _b_5680(.a(_w_7105),.q(_w_7106));
  bfr _b_5679(.a(G177),.q(_w_7105));
  bfr _b_5678(.a(_w_7103),.q(_w_7089));
  bfr _b_5677(.a(_w_7102),.q(_w_7103));
  bfr _b_5674(.a(_w_7099),.q(_w_7100));
  bfr _b_5673(.a(_w_7098),.q(_w_7099));
  bfr _b_5671(.a(_w_7096),.q(_w_7097));
  bfr _b_5670(.a(_w_7095),.q(_w_7096));
  bfr _b_5669(.a(_w_7094),.q(_w_7095));
  bfr _b_5668(.a(_w_7093),.q(_w_7094));
  bfr _b_5666(.a(_w_7091),.q(_w_7092));
  bfr _b_5664(.a(G176),.q(_w_7090));
  bfr _b_5663(.a(_w_7088),.q(_w_7060));
  bfr _b_5662(.a(_w_7087),.q(_w_7088));
  bfr _b_5660(.a(_w_7085),.q(_w_7086));
  bfr _b_5659(.a(_w_7084),.q(_w_7085));
  bfr _b_6724(.a(_w_8149),.q(_w_8150));
  bfr _b_5658(.a(_w_7083),.q(_w_7084));
  bfr _b_5657(.a(_w_7082),.q(_w_7083));
  bfr _b_5653(.a(_w_7078),.q(_w_7079));
  bfr _b_5650(.a(_w_7075),.q(_w_7076));
  bfr _b_7259(.a(_w_8684),.q(_w_8685));
  bfr _b_6018(.a(_w_7443),.q(_w_7444));
  bfr _b_5649(.a(_w_7074),.q(_w_7075));
  bfr _b_7109(.a(_w_8534),.q(_w_8535));
  bfr _b_5736(.a(_w_7161),.q(_w_7162));
  bfr _b_5647(.a(_w_7072),.q(_w_7073));
  bfr _b_5646(.a(_w_7071),.q(_w_7072));
  bfr _b_5644(.a(_w_7069),.q(_w_7070));
  bfr _b_5642(.a(_w_7067),.q(_w_7068));
  bfr _b_5641(.a(_w_7066),.q(_w_7067));
  bfr _b_5985(.a(_w_7410),.q(_w_7409));
  bfr _b_5640(.a(_w_7065),.q(_w_7066));
  bfr _b_5639(.a(_w_7064),.q(_w_7065));
  bfr _b_5638(.a(_w_7063),.q(_w_7064));
  bfr _b_5635(.a(G175),.q(_w_7061));
  bfr _b_5632(.a(_w_7057),.q(_w_7058));
  bfr _b_5631(.a(_w_7056),.q(_w_7057));
  bfr _b_5629(.a(_w_7054),.q(_w_7055));
  bfr _b_5628(.a(_w_7053),.q(_w_7054));
  bfr _b_5623(.a(_w_7048),.q(_w_7049));
  bfr _b_5619(.a(_w_7044),.q(_w_7045));
  bfr _b_5618(.a(_w_7043),.q(_w_7044));
  bfr _b_5617(.a(_w_7042),.q(_w_7043));
  bfr _b_5616(.a(_w_7041),.q(_w_7042));
  bfr _b_5614(.a(_w_7039),.q(_w_7040));
  bfr _b_5613(.a(_w_7038),.q(_w_7039));
  bfr _b_5612(.a(_w_7037),.q(_w_7038));
  bfr _b_7400(.a(_w_8825),.q(_w_8826));
  bfr _b_5611(.a(_w_7036),.q(_w_7037));
  bfr _b_5610(.a(_w_7035),.q(_w_7036));
  bfr _b_5607(.a(G174),.q(_w_7033));
  bfr _b_5605(.a(_w_7030),.q(_w_7031));
  bfr _b_5603(.a(_w_7028),.q(_w_7029));
  bfr _b_5602(.a(_w_7027),.q(_w_7028));
  bfr _b_6196(.a(_w_7621),.q(_w_7622));
  bfr _b_5598(.a(_w_7023),.q(_w_7024));
  bfr _b_5597(.a(_w_7022),.q(_w_7023));
  bfr _b_6057(.a(_w_7482),.q(_w_7483));
  bfr _b_5593(.a(_w_7018),.q(_w_7019));
  bfr _b_5592(.a(_w_7017),.q(_w_7018));
  bfr _b_5590(.a(_w_7015),.q(_w_7016));
  bfr _b_5585(.a(_w_7010),.q(_w_7011));
  bfr _b_5584(.a(_w_7009),.q(_w_7010));
  bfr _b_5583(.a(_w_7008),.q(_w_7009));
  bfr _b_5582(.a(_w_7007),.q(_w_7008));
  bfr _b_5580(.a(_w_7005),.q(_w_7006));
  bfr _b_5829(.a(_w_7254),.q(_w_7255));
  bfr _b_5578(.a(_w_7003),.q(_w_6975));
  bfr _b_5577(.a(_w_7002),.q(_w_7003));
  bfr _b_5837(.a(_w_7262),.q(_w_7263));
  bfr _b_5575(.a(_w_7000),.q(_w_7001));
  bfr _b_5574(.a(_w_6999),.q(_w_7000));
  bfr _b_5573(.a(_w_6998),.q(_w_6999));
  bfr _b_5572(.a(_w_6997),.q(_w_6998));
  bfr _b_5825(.a(_w_7250),.q(_w_7251));
  bfr _b_5571(.a(_w_6996),.q(_w_6997));
  bfr _b_5568(.a(_w_6993),.q(_w_6994));
  bfr _b_5566(.a(_w_6991),.q(_w_6992));
  bfr _b_5565(.a(_w_6990),.q(_w_6991));
  bfr _b_7206(.a(_w_8631),.q(_w_8632));
  bfr _b_5563(.a(_w_6988),.q(_w_6989));
  bfr _b_5560(.a(_w_6985),.q(_w_6986));
  bfr _b_5558(.a(_w_6983),.q(_w_6984));
  bfr _b_5557(.a(_w_6982),.q(_w_6983));
  bfr _b_5553(.a(_w_6978),.q(_w_6979));
  bfr _b_5552(.a(_w_6977),.q(_w_6978));
  bfr _b_5549(.a(_w_6974),.q(_w_6961));
  bfr _b_5548(.a(_w_6973),.q(_w_6974));
  bfr _b_5546(.a(_w_6971),.q(_w_6972));
  bfr _b_5545(.a(_w_6970),.q(_w_6971));
  bfr _b_5544(.a(_w_6969),.q(_w_6970));
  bfr _b_6702(.a(_w_8127),.q(_w_8128));
  bfr _b_5541(.a(_w_6966),.q(_w_6967));
  bfr _b_6552(.a(_w_7977),.q(_w_7978));
  bfr _b_5540(.a(_w_6965),.q(_w_6966));
  bfr _b_5537(.a(_w_6962),.q(_w_6963));
  bfr _b_5534(.a(_w_6959),.q(_w_6960));
  bfr _b_5532(.a(_w_6957),.q(_w_6958));
  bfr _b_5531(.a(_w_6956),.q(_w_6957));
  bfr _b_5530(.a(_w_6955),.q(_w_6956));
  bfr _b_5528(.a(_w_6953),.q(_w_6954));
  bfr _b_5526(.a(_w_6951),.q(_w_6952));
  bfr _b_5524(.a(G170),.q(_w_6950));
  bfr _b_5523(.a(_w_6948),.q(_w_6916));
  bfr _b_5515(.a(_w_6940),.q(_w_6941));
  bfr _b_5514(.a(_w_6939),.q(_w_6940));
  bfr _b_5512(.a(_w_6937),.q(_w_6938));
  bfr _b_6079(.a(_w_7504),.q(_w_7505));
  bfr _b_5511(.a(_w_6936),.q(_w_6937));
  bfr _b_5510(.a(_w_6935),.q(_w_6936));
  bfr _b_5508(.a(_w_6933),.q(_w_6934));
  bfr _b_5507(.a(_w_6932),.q(_w_6933));
  bfr _b_5505(.a(_w_6930),.q(_w_6931));
  bfr _b_6184(.a(_w_7609),.q(_w_7610));
  bfr _b_5504(.a(_w_6929),.q(_w_6930));
  bfr _b_5501(.a(_w_6926),.q(_w_6927));
  bfr _b_5500(.a(_w_6925),.q(_w_6926));
  bfr _b_5496(.a(_w_6921),.q(_w_6922));
  bfr _b_5495(.a(_w_6920),.q(_w_6921));
  bfr _b_5494(.a(_w_6919),.q(_w_6920));
  bfr _b_5492(.a(_w_6917),.q(_w_6918));
  bfr _b_5489(.a(_w_6914),.q(_w_6907));
  bfr _b_5488(.a(_w_6913),.q(_w_6914));
  bfr _b_5487(.a(_w_6912),.q(_w_6913));
  bfr _b_5485(.a(_w_6910),.q(_w_6911));
  bfr _b_5483(.a(_w_6908),.q(_w_6909));
  bfr _b_7171(.a(_w_8596),.q(_w_8597));
  bfr _b_5482(.a(G162),.q(_w_6908));
  bfr _b_5481(.a(_w_6906),.q(_w_6877));
  bfr _b_5479(.a(_w_6904),.q(_w_6905));
  bfr _b_7107(.a(_w_8532),.q(_w_8533));
  bfr _b_5478(.a(_w_6903),.q(_w_6904));
  bfr _b_5477(.a(_w_6902),.q(_w_6903));
  bfr _b_5473(.a(_w_6898),.q(_w_6899));
  bfr _b_5472(.a(_w_6897),.q(_w_6898));
  bfr _b_5471(.a(_w_6896),.q(_w_6897));
  bfr _b_5469(.a(_w_6894),.q(_w_6895));
  bfr _b_5468(.a(_w_6893),.q(_w_6894));
  bfr _b_5467(.a(_w_6892),.q(_w_6893));
  bfr _b_5466(.a(_w_6891),.q(_w_6892));
  bfr _b_5465(.a(_w_6890),.q(_w_6891));
  bfr _b_5464(.a(_w_6889),.q(_w_6890));
  bfr _b_5462(.a(_w_6887),.q(_w_6888));
  bfr _b_7522(.a(_w_8947),.q(_w_8946));
  bfr _b_5460(.a(_w_6885),.q(_w_6886));
  bfr _b_5456(.a(_w_6881),.q(_w_6882));
  bfr _b_5454(.a(_w_6879),.q(_w_6880));
  bfr _b_7127(.a(_w_8552),.q(_w_8553));
  bfr _b_5453(.a(_w_6878),.q(_w_6879));
  bfr _b_5451(.a(_w_6876),.q(_w_6848));
  bfr _b_5449(.a(_w_6874),.q(_w_6875));
  bfr _b_7354(.a(_w_8779),.q(_w_8780));
  bfr _b_5445(.a(_w_6870),.q(_w_6871));
  bfr _b_5441(.a(_w_6866),.q(_w_6867));
  bfr _b_5440(.a(_w_6865),.q(_w_6866));
  bfr _b_5437(.a(_w_6862),.q(_w_6863));
  bfr _b_5436(.a(_w_6861),.q(_w_6862));
  bfr _b_7008(.a(_w_8433),.q(_w_8400));
  bfr _b_6287(.a(_w_7712),.q(_w_7713));
  bfr _b_5434(.a(_w_6859),.q(_w_6860));
  bfr _b_5433(.a(_w_6858),.q(_w_6859));
  bfr _b_5432(.a(_w_6857),.q(_w_6858));
  bfr _b_5431(.a(_w_6856),.q(_w_6857));
  bfr _b_5430(.a(_w_6855),.q(_w_6856));
  bfr _b_5429(.a(_w_6854),.q(_w_6855));
  bfr _b_5426(.a(_w_6851),.q(_w_6852));
  bfr _b_5423(.a(G160),.q(_w_6849));
  bfr _b_5422(.a(_w_6847),.q(_w_6816));
  bfr _b_5421(.a(_w_6846),.q(_w_6847));
  bfr _b_5419(.a(_w_6844),.q(_w_6845));
  bfr _b_5418(.a(_w_6843),.q(_w_6844));
  bfr _b_5417(.a(_w_6842),.q(_w_6843));
  bfr _b_5414(.a(_w_6839),.q(_w_6840));
  bfr _b_5411(.a(_w_6836),.q(_w_6837));
  bfr _b_5408(.a(_w_6833),.q(_w_6834));
  bfr _b_5406(.a(_w_6831),.q(_w_6832));
  bfr _b_5405(.a(_w_6830),.q(_w_6831));
  bfr _b_5404(.a(_w_6829),.q(_w_6830));
  bfr _b_5402(.a(_w_6827),.q(_w_6828));
  bfr _b_5401(.a(_w_6826),.q(_w_6827));
  bfr _b_5400(.a(_w_6825),.q(_w_6826));
  bfr _b_5399(.a(_w_6824),.q(_w_6825));
  bfr _b_5397(.a(_w_6822),.q(_w_6823));
  bfr _b_5396(.a(_w_6821),.q(_w_6822));
  bfr _b_5393(.a(_w_6818),.q(_w_6819));
  bfr _b_5392(.a(_w_6817),.q(_w_6818));
  bfr _b_5391(.a(G16),.q(_w_6817));
  bfr _b_6859(.a(_w_8284),.q(_w_8285));
  bfr _b_5390(.a(_w_6815),.q(_w_6786));
  bfr _b_5387(.a(_w_6812),.q(_w_6813));
  bfr _b_5386(.a(_w_6811),.q(_w_6812));
  bfr _b_6467(.a(_w_7892),.q(_w_7893));
  bfr _b_5385(.a(_w_6810),.q(_w_6811));
  bfr _b_5384(.a(_w_6809),.q(_w_6810));
  bfr _b_5383(.a(_w_6808),.q(_w_6809));
  bfr _b_5380(.a(_w_6805),.q(_w_6806));
  bfr _b_5377(.a(_w_6802),.q(_w_6803));
  bfr _b_5376(.a(_w_6801),.q(_w_6802));
  bfr _b_5927(.a(_w_7352),.q(_w_7353));
  bfr _b_5372(.a(_w_6797),.q(_w_6798));
  bfr _b_5370(.a(_w_6795),.q(_w_6796));
  bfr _b_5369(.a(_w_6794),.q(_w_6795));
  bfr _b_5366(.a(_w_6791),.q(_w_6792));
  bfr _b_7427(.a(_w_8852),.q(_w_8853));
  bfr _b_5365(.a(_w_6790),.q(_w_6791));
  bfr _b_5364(.a(_w_6789),.q(_w_6790));
  bfr _b_5363(.a(_w_6788),.q(_w_6789));
  bfr _b_5738(.a(_w_7163),.q(_w_7164));
  bfr _b_5362(.a(_w_6787),.q(_w_6788));
  bfr _b_5361(.a(G159),.q(_w_6787));
  bfr _b_5359(.a(_w_6784),.q(_w_6785));
  bfr _b_7270(.a(_w_8695),.q(_w_8696));
  bfr _b_5358(.a(_w_6783),.q(_w_6784));
  bfr _b_5357(.a(_w_6782),.q(_w_6783));
  bfr _b_5356(.a(_w_6781),.q(_w_6782));
  bfr _b_5634(.a(_w_7059),.q(_w_7032));
  bfr _b_5354(.a(_w_6779),.q(_w_6780));
  bfr _b_5352(.a(_w_6777),.q(_w_6778));
  bfr _b_5348(.a(_w_6773),.q(_w_6774));
  bfr _b_5347(.a(_w_6772),.q(_w_6773));
  bfr _b_5863(.a(_w_7288),.q(_w_7289));
  bfr _b_5346(.a(_w_6771),.q(_w_6772));
  bfr _b_5344(.a(_w_6769),.q(_w_6770));
  bfr _b_5342(.a(_w_6767),.q(_w_6768));
  bfr _b_7363(.a(_w_8788),.q(_w_8789));
  bfr _b_5341(.a(_w_6766),.q(_w_6767));
  bfr _b_5339(.a(_w_6764),.q(_w_6765));
  bfr _b_6976(.a(_w_8401),.q(_w_8402));
  bfr _b_5338(.a(_w_6763),.q(_w_6764));
  bfr _b_5337(.a(_w_6762),.q(_w_6763));
  bfr _b_5334(.a(_w_6759),.q(_w_6760));
  bfr _b_5330(.a(_w_6755),.q(_w_6756));
  bfr _b_5329(.a(_w_6754),.q(_w_6755));
  bfr _b_5327(.a(_w_6752),.q(_w_6753));
  bfr _b_5325(.a(_w_6750),.q(_w_6751));
  bfr _b_5323(.a(_w_6748),.q(_w_6749));
  bfr _b_5321(.a(_w_6746),.q(_w_6747));
  bfr _b_5319(.a(_w_6744),.q(_w_6745));
  bfr _b_5318(.a(_w_6743),.q(_w_6744));
  bfr _b_5315(.a(_w_6740),.q(_w_6741));
  bfr _b_5314(.a(_w_6739),.q(_w_6740));
  bfr _b_5311(.a(G157),.q(_w_6737));
  bfr _b_5308(.a(_w_6733),.q(_w_6734));
  bfr _b_6200(.a(_w_7625),.q(_w_7626));
  bfr _b_5307(.a(_w_6732),.q(_w_6733));
  bfr _b_5305(.a(_w_6730),.q(_w_6731));
  bfr _b_5304(.a(_w_6729),.q(_w_6730));
  bfr _b_5303(.a(_w_6728),.q(_w_6729));
  bfr _b_5302(.a(_w_6727),.q(_w_6728));
  bfr _b_5300(.a(_w_6725),.q(_w_6726));
  bfr _b_5299(.a(_w_6724),.q(_w_6725));
  bfr _b_5298(.a(_w_6723),.q(_w_6724));
  bfr _b_5297(.a(_w_6722),.q(_w_6723));
  bfr _b_5296(.a(_w_6721),.q(_w_6722));
  bfr _b_5295(.a(_w_6720),.q(_w_6721));
  bfr _b_5291(.a(_w_6716),.q(_w_6717));
  bfr _b_6213(.a(_w_7638),.q(_w_7639));
  bfr _b_5290(.a(_w_6715),.q(_w_6716));
  bfr _b_5288(.a(_w_6713),.q(_w_6714));
  bfr _b_7208(.a(_w_8633),.q(_w_8634));
  bfr _b_5286(.a(_w_6711),.q(_w_6712));
  bfr _b_5285(.a(_w_6710),.q(_w_6711));
  bfr _b_5281(.a(_w_6706),.q(_w_6707));
  bfr _b_5279(.a(G156),.q(_w_6705));
  bfr _b_5277(.a(_w_6702),.q(_w_6703));
  bfr _b_6684(.a(_w_8109),.q(_w_8110));
  bfr _b_5274(.a(_w_6699),.q(_w_6700));
  bfr _b_5272(.a(_w_6697),.q(_w_6698));
  bfr _b_5271(.a(_w_6696),.q(_w_6697));
  bfr _b_5270(.a(_w_6695),.q(_w_6696));
  bfr _b_5269(.a(_w_6694),.q(_w_6695));
  bfr _b_5268(.a(_w_6693),.q(_w_6694));
  bfr _b_5267(.a(_w_6692),.q(_w_6693));
  bfr _b_7310(.a(_w_8735),.q(_w_8736));
  bfr _b_5265(.a(_w_6690),.q(_w_6691));
  bfr _b_5264(.a(_w_6689),.q(_w_6690));
  bfr _b_6397(.a(_w_7822),.q(_w_7823));
  bfr _b_6095(.a(_w_7520),.q(_w_7521));
  bfr _b_5263(.a(_w_6688),.q(_w_6689));
  bfr _b_5262(.a(_w_6687),.q(_w_6688));
  bfr _b_5260(.a(_w_6685),.q(_w_6686));
  bfr _b_5259(.a(_w_6684),.q(_w_6685));
  bfr _b_5258(.a(_w_6683),.q(_w_6684));
  bfr _b_5257(.a(_w_6682),.q(_w_6683));
  bfr _b_5256(.a(_w_6681),.q(_w_6682));
  bfr _b_5253(.a(_w_6678),.q(_w_6679));
  bfr _b_5250(.a(_w_6675),.q(_w_6676));
  bfr _b_5249(.a(_w_6674),.q(_w_6675));
  bfr _b_5353(.a(_w_6778),.q(_w_6779));
  bfr _b_5248(.a(_w_6673),.q(_w_6674));
  bfr _b_5247(.a(G155),.q(_w_6673));
  bfr _b_5282(.a(_w_6707),.q(_w_6708));
  bfr _b_5246(.a(_w_6671),.q(_w_6640));
  bfr _b_7352(.a(_w_8777),.q(_w_8778));
  bfr _b_5244(.a(_w_6669),.q(_w_6670));
  bfr _b_5992(.a(_w_7417),.q(_w_7418));
  bfr _b_5243(.a(_w_6668),.q(_w_6669));
  bfr _b_7193(.a(_w_8618),.q(_w_8619));
  bfr _b_6028(.a(G33),.q(_w_7454));
  bfr _b_5240(.a(_w_6665),.q(_w_6666));
  bfr _b_5239(.a(_w_6664),.q(_w_6665));
  bfr _b_5237(.a(_w_6662),.q(_w_6663));
  bfr _b_5235(.a(_w_6660),.q(_w_6661));
  bfr _b_5231(.a(_w_6656),.q(_w_6657));
  bfr _b_5230(.a(_w_6655),.q(_w_6656));
  bfr _b_6904(.a(_w_8329),.q(_w_8296));
  bfr _b_6365(.a(_w_7790),.q(_w_7791));
  bfr _b_5229(.a(_w_6654),.q(_w_6655));
  bfr _b_5224(.a(_w_6649),.q(_w_6650));
  bfr _b_5223(.a(_w_6648),.q(_w_6649));
  bfr _b_5220(.a(_w_6645),.q(_w_6646));
  bfr _b_5219(.a(_w_6644),.q(_w_6645));
  bfr _b_5217(.a(_w_6642),.q(_w_6643));
  bfr _b_5216(.a(_w_6641),.q(_w_6642));
  bfr _b_5215(.a(G153),.q(_w_6641));
  bfr _b_5214(.a(_w_6639),.q(_w_6602));
  bfr _b_5212(.a(_w_6637),.q(_w_6638));
  bfr _b_6475(.a(_w_7900),.q(_w_7901));
  bfr _b_5211(.a(_w_6636),.q(_w_6637));
  bfr _b_5210(.a(_w_6635),.q(_w_6636));
  bfr _b_5209(.a(_w_6634),.q(_w_6635));
  bfr _b_5208(.a(_w_6633),.q(_w_6634));
  bfr _b_5207(.a(_w_6632),.q(_w_6633));
  bfr _b_5205(.a(_w_6630),.q(_w_6631));
  bfr _b_5204(.a(_w_6629),.q(_w_6630));
  bfr _b_5203(.a(_w_6628),.q(_w_6629));
  bfr _b_5201(.a(_w_6626),.q(_w_6627));
  bfr _b_5199(.a(_w_6624),.q(_w_6625));
  bfr _b_5198(.a(_w_6623),.q(_w_6624));
  bfr _b_5197(.a(_w_6622),.q(_w_6623));
  bfr _b_5196(.a(_w_6621),.q(_w_6622));
  bfr _b_5194(.a(_w_6619),.q(_w_6620));
  bfr _b_5192(.a(_w_6617),.q(_w_6618));
  bfr _b_5191(.a(_w_6616),.q(_w_6617));
  bfr _b_6668(.a(_w_8093),.q(_w_8094));
  bfr _b_5190(.a(_w_6615),.q(_w_6616));
  bfr _b_5188(.a(_w_6613),.q(_w_6614));
  bfr _b_5891(.a(_w_7316),.q(_w_7317));
  bfr _b_5187(.a(_w_6612),.q(_w_6613));
  bfr _b_5184(.a(_w_6609),.q(_w_6610));
  bfr _b_5183(.a(_w_6608),.q(_w_6609));
  bfr _b_5182(.a(_w_6607),.q(_w_6608));
  bfr _b_5180(.a(_w_6605),.q(_w_6606));
  bfr _b_5179(.a(_w_6604),.q(_w_6605));
  bfr _b_5176(.a(_w_6601),.q(_w_6599));
  bfr _b_5174(.a(G150),.q(_w_6600));
  bfr _b_5173(.a(_w_6598),.q(_w_6566));
  bfr _b_5172(.a(_w_6597),.q(_w_6598));
  bfr _b_5171(.a(_w_6596),.q(_w_6597));
  bfr _b_5168(.a(_w_6593),.q(_w_6594));
  bfr _b_5167(.a(_w_6592),.q(_w_6593));
  bfr _b_5166(.a(_w_6591),.q(_w_6592));
  bfr _b_5165(.a(_w_6590),.q(_w_6591));
  bfr _b_5164(.a(_w_6589),.q(_w_6590));
  bfr _b_5163(.a(_w_6588),.q(_w_6589));
  bfr _b_5161(.a(_w_6586),.q(_w_6587));
  bfr _b_5155(.a(_w_6580),.q(_w_6581));
  bfr _b_5153(.a(_w_6578),.q(_w_6579));
  bfr _b_5152(.a(_w_6577),.q(_w_6578));
  bfr _b_5151(.a(_w_6576),.q(_w_6577));
  bfr _b_5145(.a(_w_6570),.q(_w_6571));
  bfr _b_5143(.a(_w_6568),.q(_w_6569));
  bfr _b_5142(.a(_w_6567),.q(_w_6568));
  bfr _b_5141(.a(G15),.q(_w_6567));
  bfr _b_5878(.a(_w_7303),.q(_w_7304));
  bfr _b_5137(.a(G148),.q(_w_6562));
  bfr _b_5135(.a(_w_6560),.q(_w_6561));
  bfr _b_5134(.a(G147),.q(_w_6560));
  bfr _b_5131(.a(_w_6556),.q(_w_6557));
  bfr _b_5129(.a(_w_6554),.q(_w_6555));
  bfr _b_5127(.a(_w_6552),.q(_w_6553));
  bfr _b_5125(.a(G146),.q(_w_6551));
  bfr _b_5124(.a(_w_6549),.q(_w_6541));
  bfr _b_5123(.a(_w_6548),.q(_w_6549));
  bfr _b_7558(.a(_w_8983),.q(_w_8984));
  bfr _b_5122(.a(_w_6547),.q(_w_6548));
  bfr _b_5398(.a(_w_6823),.q(_w_6824));
  bfr _b_5121(.a(_w_6546),.q(_w_6547));
  bfr _b_5120(.a(_w_6545),.q(_w_6546));
  bfr _b_5119(.a(_w_6544),.q(_w_6545));
  bfr _b_5117(.a(_w_6542),.q(_w_6543));
  bfr _b_5114(.a(_w_6539),.q(_w_6540));
  bfr _b_5113(.a(G144),.q(_w_6539));
  bfr _b_5111(.a(_w_6536),.q(_w_6537));
  bfr _b_7269(.a(_w_8694),.q(_w_8695));
  bfr _b_5110(.a(G143),.q(_w_6536));
  bfr _b_6276(.a(_w_7701),.q(_w_7702));
  bfr _b_5106(.a(G142),.q(_w_6532));
  bfr _b_6585(.a(_w_8010),.q(_w_8011));
  bfr _b_5615(.a(_w_7040),.q(_w_7041));
  bfr _b_5105(.a(_w_6530),.q(_w_6528));
  bfr _b_5104(.a(_w_6529),.q(_w_6530));
  bfr _b_5103(.a(G141),.q(_w_6529));
  bfr _b_7144(.a(G77),.q(_w_8570));
  bfr _b_5102(.a(_w_6527),.q(_w_6525));
  bfr _b_5503(.a(_w_6928),.q(_w_6929));
  bfr _b_5101(.a(_w_6526),.q(_w_6527));
  bfr _b_5100(.a(G140),.q(_w_6526));
  bfr _b_5099(.a(_w_6524),.q(_w_6493));
  bfr _b_5095(.a(_w_6520),.q(_w_6521));
  bfr _b_5094(.a(_w_6519),.q(_w_6520));
  bfr _b_5091(.a(_w_6516),.q(_w_6517));
  bfr _b_5088(.a(_w_6513),.q(_w_6514));
  bfr _b_7233(.a(_w_8658),.q(_w_8659));
  spl4L G175_s_0(.a(_w_7060),.q0(_w_3747),.q1(G175_1),.q2(_w_3749),.q3(_w_3751));
  bfr _b_2581(.a(_w_4006),.q(G5242));
  bfr _b_2352(.a(_w_3777),.q(_w_3778));
  spl2 G126_s_1(.a(G126_1),.q0(G126_4),.q1(G126_5));
  bfr _b_7010(.a(_w_8435),.q(_w_8436));
  spl4L g537_s_0(.a(n537),.q0(_w_3972),.q1(n537_1),.q2(n537_2),.q3(n537_3));
  bfr _b_5589(.a(_w_7014),.q(_w_7015));
  bfr _b_5218(.a(_w_6643),.q(_w_6644));
  and_bb g848(.a(G24_0),.b(n586_6),.q(n848));
  bfr _b_2128(.a(_w_3553),.q(_w_3554));
  bfr _b_7543(.a(_w_8968),.q(_w_8969));
  spl4L g464_s_0(.a(n464),.q0(n464_0),.q1(_w_3467),.q2(n464_2),.q3(n464_3));
  bfr _b_2339(.a(_w_3764),.q(_w_3765));
  bfr _b_2336(.a(_w_3761),.q(_w_3762));
  bfr _b_7224(.a(_w_8649),.q(_w_8650));
  bfr _b_2334(.a(_w_3759),.q(_w_3760));
  bfr _b_4493(.a(_w_5918),.q(_w_5919));
  bfr _b_2332(.a(_w_3757),.q(_w_3758));
  bfr _b_7243(.a(_w_8668),.q(_w_8669));
  inv inv_G114(.a(G114_1),.q(i_G114));
  bfr _b_5608(.a(_w_7033),.q(_w_7034));
  bfr _b_2331(.a(_w_3756),.q(_w_3757));
  bfr _b_6326(.a(_w_7751),.q(_w_7752));
  and_bi g659(.a(n658_0),.b(G176_49),.q(n659));
  bfr _b_3648(.a(_w_5073),.q(n427_2));
  or_bb g1042(.a(n1040),.b(n1041),.q(n1042));
  bfr _b_6093(.a(_w_7518),.q(_w_7519));
  bfr _b_2323(.a(_w_3748),.q(G175_0));
  bfr _b_2322(.a(_w_3747),.q(_w_3748));
  and_bi g332(.a(G139_0),.b(n331),.q(n332));
  bfr _b_5415(.a(_w_6840),.q(_w_6841));
  bfr _b_2638(.a(_w_4063),.q(_w_4064));
  bfr _b_2318(.a(_w_3743),.q(_w_3744));
  bfr _b_2310(.a(_w_3735),.q(G174_20));
  bfr _b_3430(.a(_w_4855),.q(_w_4856));
  bfr _b_2307(.a(_w_3732),.q(G173_6));
  bfr _b_2290(.a(_w_3715),.q(_w_3716));
  bfr _b_2288(.a(_w_3713),.q(_w_3714));
  bfr _b_2282(.a(_w_3707),.q(_w_3708));
  bfr _b_2280(.a(_w_3705),.q(_w_3706));
  bfr _b_2279(.a(_w_3704),.q(_w_3705));
  bfr _b_4499(.a(_w_5924),.q(n451_1));
  bfr _b_2297(.a(_w_3722),.q(_w_3723));
  bfr _b_4023(.a(_w_5448),.q(_w_5449));
  bfr _b_2277(.a(_w_3702),.q(_w_3703));
  bfr _b_6007(.a(_w_7432),.q(_w_7433));
  spl2 G27_s_0(.a(_w_7376),.q0(G27_0),.q1(G27_1));
  bfr _b_2275(.a(_w_3700),.q(_w_3701));
  and_bb g1127(.a(G64_11),.b(n1126),.q(_w_6293));
  bfr _b_2270(.a(_w_3695),.q(_w_3696));
  bfr _b_2268(.a(_w_3693),.q(_w_3694));
  bfr _b_2267(.a(_w_3692),.q(_w_3693));
  bfr _b_6060(.a(_w_7485),.q(_w_7486));
  bfr _b_2266(.a(_w_3691),.q(_w_3692));
  bfr _b_4442(.a(_w_5867),.q(n818));
  bfr _b_2265(.a(_w_3690),.q(_w_3691));
  inv inv_G155(.a(G155_1),.q(G5209));
  bfr _b_2260(.a(_w_3685),.q(_w_3686));
  bfr _b_2252(.a(_w_3677),.q(_w_3678));
  bfr _b_2736(.a(_w_4161),.q(_w_4162));
  bfr _b_2248(.a(_w_3673),.q(_w_3674));
  bfr _b_7225(.a(_w_8650),.q(_w_8651));
  bfr _b_2246(.a(_w_3671),.q(_w_3672));
  bfr _b_2245(.a(_w_3670),.q(G158_18));
  spl2 g704_s_0(.a(n704),.q0(n704_0),.q1(n704_1));
  bfr _b_6187(.a(_w_7612),.q(_w_7613));
  bfr _b_2242(.a(_w_3667),.q(G158_16));
  bfr _b_2632(.a(_w_4057),.q(_w_4058));
  bfr _b_2238(.a(_w_3663),.q(G158_24));
  bfr _b_3258(.a(_w_4683),.q(_w_4684));
  bfr _b_2236(.a(_w_3661),.q(G155_1));
  bfr _b_2233(.a(_w_3658),.q(_w_3659));
  bfr _b_2232(.a(_w_3657),.q(_w_3658));
  bfr _b_6951(.a(_w_8376),.q(_w_8377));
  bfr _b_2231(.a(_w_3656),.q(_w_3657));
  bfr _b_2228(.a(_w_3653),.q(G5219));
  spl2 g731_s_0(.a(n731),.q0(n731_0),.q1(n731_1));
  bfr _b_6937(.a(_w_8362),.q(_w_8363));
  bfr _b_2222(.a(_w_3647),.q(G141_2));
  bfr _b_5851(.a(_w_7276),.q(_w_7244));
  bfr _b_2221(.a(_w_3646),.q(_w_3647));
  bfr _b_2217(.a(_w_3642),.q(G168_0));
  bfr _b_2208(.a(_w_3633),.q(_w_3634));
  and_bi g209(.a(n208),.b(n206),.q(_w_5005));
  bfr _b_2207(.a(_w_3632),.q(_w_3633));
  bfr _b_2006(.a(_w_3431),.q(_w_3432));
  bfr _b_4572(.a(_w_5997),.q(_w_5998));
  bfr _b_6114(.a(_w_7539),.q(_w_7540));
  bfr _b_2204(.a(_w_3629),.q(_w_3630));
  bfr _b_2612(.a(_w_4037),.q(_w_4038));
  bfr _b_2192(.a(_w_3617),.q(_w_3618));
  bfr _b_6376(.a(_w_7801),.q(_w_7802));
  bfr _b_2189(.a(_w_3614),.q(_w_3615));
  bfr _b_2185(.a(_w_3610),.q(_w_3611));
  bfr _b_4228(.a(_w_5653),.q(_w_5654));
  bfr _b_2274(.a(_w_3699),.q(_w_3700));
  or_bb g541(.a(n373_1),.b(n540),.q(_w_5682));
  bfr _b_2173(.a(_w_3598),.q(_w_3599));
  bfr _b_5502(.a(_w_6927),.q(_w_6928));
  bfr _b_2922(.a(_w_4347),.q(_w_4348));
  and_bb g1100(.a(G64_14),.b(n1099),.q(_w_5701));
  bfr _b_6176(.a(_w_7601),.q(_w_7602));
  bfr _b_2313(.a(_w_3738),.q(G174_16));
  spl4L g442_s_0(.a(n442),.q0(n442_0),.q1(n442_1),.q2(n442_2),.q3(n442_3));
  spl4L g663_s_0(.a(G5258_0),.q0(_w_4018),.q1(G5258_1),.q2(G5258_2),.q3(G5258_3));
  bfr _b_2261(.a(_w_3686),.q(_w_3687));
  spl2 G109_s_1(.a(G109_1),.q0(G109_4),.q1(G109_5));
  and_bb g1141(.a(G85_1),.b(n815_8),.q(n1141));
  bfr _b_2400(.a(_w_3825),.q(_w_3826));
  bfr _b_2764(.a(_w_4189),.q(n387_2));
  bfr _b_2163(.a(_w_3588),.q(_w_3589));
  bfr _b_5252(.a(_w_6677),.q(_w_6678));
  spl3L G111_s_0(.a(_w_6406),.q0(G111_0),.q1(G111_1),.q2(G111_2));
  bfr _b_2158(.a(_w_3583),.q(_w_3584));
  bfr _b_5543(.a(_w_6968),.q(_w_6969));
  bfr _b_2154(.a(_w_3579),.q(_w_3580));
  bfr _b_3329(.a(_w_4754),.q(_w_4755));
  bfr _b_2150(.a(_w_3575),.q(_w_3576));
  bfr _b_2148(.a(_w_3573),.q(_w_3574));
  bfr _b_2147(.a(_w_3572),.q(_w_3573));
  bfr _b_2285(.a(_w_3710),.q(_w_3711));
  spl4L G126_s_2(.a(G126_2),.q0(G126_6),.q1(G126_7),.q2(G126_8),.q3(G126_9));
  and_bi g221(.a(G98_4),.b(G117_4),.q(n221));
  bfr _b_6708(.a(_w_8133),.q(_w_8113));
  bfr _b_2145(.a(_w_3570),.q(_w_3571));
  bfr _b_2144(.a(_w_3569),.q(_w_3570));
  bfr _b_2505(.a(_w_3930),.q(n249_1));
  bfr _b_2140(.a(_w_3565),.q(_w_3566));
  bfr _b_2139(.a(_w_3564),.q(_w_3565));
  bfr _b_2136(.a(_w_3561),.q(_w_3562));
  bfr _b_2109(.a(_w_3534),.q(_w_3535));
  bfr _b_5867(.a(_w_7292),.q(_w_7293));
  bfr _b_2134(.a(_w_3559),.q(G131_1));
  bfr _b_5694(.a(_w_7119),.q(_w_7104));
  bfr _b_2133(.a(_w_3558),.q(_w_3559));
  bfr _b_4535(.a(_w_5960),.q(_w_5961));
  bfr _b_2127(.a(_w_3552),.q(_w_3553));
  bfr _b_2126(.a(_w_3551),.q(_w_3552));
  bfr _b_2351(.a(_w_3776),.q(_w_3777));
  bfr _b_2545(.a(_w_3970),.q(_w_3971));
  bfr _b_3774(.a(_w_5199),.q(_w_5200));
  bfr _b_5698(.a(_w_7123),.q(_w_7124));
  bfr _b_2120(.a(_w_3545),.q(_w_3546));
  bfr _b_2113(.a(_w_3538),.q(_w_3539));
  bfr _b_2112(.a(_w_3537),.q(_w_3538));
  bfr _b_6319(.a(_w_7744),.q(_w_7745));
  bfr _b_3051(.a(_w_4476),.q(n365));
  bfr _b_2106(.a(_w_3531),.q(_w_3532));
  bfr _b_5588(.a(_w_7013),.q(_w_7014));
  bfr _b_2098(.a(_w_3523),.q(G121_3));
  bfr _b_5652(.a(_w_7077),.q(_w_7078));
  bfr _b_4170(.a(_w_5595),.q(_w_5596));
  bfr _b_5448(.a(_w_6873),.q(_w_6874));
  bfr _b_2093(.a(_w_3518),.q(G121_8));
  bfr _b_2087(.a(_w_3512),.q(G109_3));
  bfr _b_2082(.a(_w_3507),.q(_w_3508));
  bfr _b_6265(.a(_w_7690),.q(_w_7691));
  bfr _b_2825(.a(_w_4250),.q(_w_4251));
  bfr _b_3273(.a(_w_4698),.q(n1262));
  bfr _b_7241(.a(_w_8666),.q(_w_8667));
  bfr _b_2081(.a(_w_3506),.q(_w_3507));
  bfr _b_4111(.a(_w_5536),.q(_w_5537));
  bfr _b_5351(.a(_w_6776),.q(_w_6777));
  bfr _b_2079(.a(_w_3504),.q(G103_0));
  bfr _b_2076(.a(_w_3501),.q(_w_3502));
  spl4L g438_s_0(.a(n438),.q0(n438_0),.q1(n438_1),.q2(n438_2),.q3(n438_3));
  bfr _b_5990(.a(_w_7415),.q(_w_7416));
  bfr _b_2463(.a(_w_3888),.q(_w_3889));
  bfr _b_5200(.a(_w_6625),.q(_w_6626));
  spl4L G138_s_0(.a(_w_6487),.q0(G138_0),.q1(G138_1),.q2(_w_4293),.q3(G138_3));
  bfr _b_2938(.a(_w_4363),.q(G5260_0));
  bfr _b_6175(.a(_w_7600),.q(_w_7601));
  and_bb g932(.a(n929),.b(n931),.q(_w_6068));
  bfr _b_2073(.a(_w_3498),.q(n449_1));
  bfr _b_2071(.a(_w_3496),.q(_w_3497));
  bfr _b_2067(.a(_w_3492),.q(_w_3493));
  bfr _b_3002(.a(_w_4427),.q(_w_4428));
  bfr _b_3827(.a(_w_5252),.q(_w_5253));
  bfr _b_2065(.a(_w_3490),.q(n457_1));
  and_bi g1175(.a(n463_5),.b(n457_2),.q(n1175));
  bfr _b_2472(.a(_w_3897),.q(_w_3898));
  bfr _b_2061(.a(_w_3486),.q(_w_3487));
  bfr _b_5645(.a(_w_7070),.q(_w_7071));
  and_bb g669(.a(n394_4),.b(n667_1),.q(n669));
  bfr _b_2723(.a(_w_4148),.q(_w_4149));
  bfr _b_6487(.a(_w_7912),.q(_w_7913));
  bfr _b_4681(.a(_w_6106),.q(_w_6107));
  bfr _b_7125(.a(_w_8550),.q(_w_8551));
  bfr _b_6130(.a(_w_7555),.q(_w_7556));
  inv inv_G151(.a(G151),.q(_w_4477));
  bfr _b_7348(.a(G83),.q(_w_8774));
  bfr _b_2051(.a(_w_3476),.q(_w_3477));
  bfr _b_6890(.a(_w_8315),.q(_w_8316));
  bfr _b_5959(.a(_w_7384),.q(_w_7385));
  bfr _b_5107(.a(_w_6532),.q(_w_6533));
  bfr _b_2338(.a(_w_3763),.q(_w_3764));
  bfr _b_2772(.a(_w_4197),.q(_w_4198));
  bfr _b_2048(.a(_w_3473),.q(n464_1));
  bfr _b_2047(.a(_w_3472),.q(_w_3473));
  and_bi g1449(.a(G172_14),.b(n1448),.q(_w_5001));
  bfr _b_4211(.a(_w_5636),.q(_w_5637));
  bfr _b_3119(.a(_w_4544),.q(_w_4545));
  bfr _b_2043(.a(_w_3468),.q(_w_3469));
  bfr _b_6252(.a(_w_7677),.q(_w_7678));
  bfr _b_2042(.a(_w_3467),.q(_w_3468));
  bfr _b_7327(.a(_w_8752),.q(_w_8753));
  bfr _b_2040(.a(_w_3465),.q(_w_3466));
  bfr _b_2039(.a(_w_3464),.q(_w_3465));
  and_bi g656(.a(n655_0),.b(n400_2),.q(n656));
  bfr _b_2038(.a(_w_3463),.q(_w_3464));
  bfr _b_2034(.a(_w_3459),.q(_w_3460));
  bfr _b_4135(.a(_w_5560),.q(_w_5561));
  bfr _b_2072(.a(_w_3497),.q(G5260));
  spl2 g1195_s_0(.a(n1195),.q0(n1195_0),.q1(n1195_1));
  bfr _b_2029(.a(_w_3454),.q(n465_0));
  bfr _b_2028(.a(_w_3453),.q(_w_3454));
  bfr _b_2026(.a(_w_3451),.q(n469_10));
  bfr _b_5413(.a(_w_6838),.q(_w_6839));
  bfr _b_4101(.a(_w_5526),.q(_w_5527));
  bfr _b_2019(.a(_w_3444),.q(n610_1));
  bfr _b_3548(.a(_w_4973),.q(_w_4974));
  bfr _b_6542(.a(_w_7967),.q(_w_7968));
  bfr _b_2018(.a(_w_3443),.q(n779_0));
  bfr _b_3807(.a(_w_5232),.q(_w_5233));
  bfr _b_6371(.a(_w_7796),.q(_w_7797));
  bfr _b_2017(.a(_w_3442),.q(G142_3));
  bfr _b_2014(.a(_w_3439),.q(G176_0));
  bfr _b_2011(.a(_w_3436),.q(_w_3437));
  bfr _b_2601(.a(_w_4026),.q(_w_4027));
  bfr _b_5963(.a(_w_7388),.q(_w_7389));
  bfr _b_2010(.a(_w_3435),.q(_w_3436));
  bfr _b_2843(.a(_w_4268),.q(_w_4269));
  bfr _b_7341(.a(_w_8766),.q(_w_8767));
  bfr _b_6258(.a(_w_7683),.q(_w_7684));
  bfr _b_2004(.a(_w_3429),.q(G176_4));
  and_bi g1288(.a(n1286),.b(n1287),.q(_w_5615));
  bfr _b_2003(.a(_w_3428),.q(_w_3429));
  spl2 g570_s_1(.a(G5249_3),.q0(G5249_4),.q1(G5249_5));
  spl2 g1211_s_0(.a(n1211),.q0(n1211_0),.q1(n1211_1));
  bfr _b_1998(.a(_w_3423),.q(_w_3424));
  bfr _b_1997(.a(_w_3422),.q(_w_3423));
  bfr _b_5672(.a(_w_7097),.q(_w_7098));
  spl2 g1317_s_0(.a(n1317),.q0(n1317_0),.q1(n1317_1));
  bfr _b_2199(.a(_w_3624),.q(_w_3625));
  bfr _b_2226(.a(_w_3651),.q(G64_0));
  spl2 g766_s_0(.a(n766),.q0(n766_0),.q1(n766_1));
  bfr _b_6555(.a(_w_7980),.q(_w_7981));
  bfr _b_1996(.a(_w_3421),.q(_w_3422));
  and_bi g1232(.a(G98_10),.b(G128_13),.q(n1232));
  bfr _b_1992(.a(_w_3417),.q(_w_3418));
  bfr _b_4921(.a(_w_6346),.q(_w_6347));
  bfr _b_2058(.a(_w_3483),.q(_w_3484));
  bfr _b_1994(.a(_w_3419),.q(_w_3420));
  bfr _b_1993(.a(_w_3418),.q(_w_3419));
  bfr _b_3723(.a(_w_5148),.q(_w_5149));
  bfr _b_1991(.a(_w_3416),.q(_w_3417));
  bfr _b_6495(.a(_w_7920),.q(_w_7921));
  and_bi g405(.a(_w_8942),.b(G124_13),.q(n405));
  bfr _b_6163(.a(_w_7588),.q(_w_7589));
  bfr _b_1989(.a(_w_3414),.q(_w_3415));
  bfr _b_6127(.a(_w_7552),.q(_w_7553));
  bfr _b_5096(.a(_w_6521),.q(_w_6522));
  or_bb g1172(.a(n1170_1),.b(n686_3),.q(n1172));
  bfr _b_1983(.a(_w_3408),.q(G176_13));
  bfr _b_1982(.a(_w_3407),.q(_w_3408));
  bfr _b_4837(.a(_w_6262),.q(_w_6263));
  bfr _b_1978(.a(_w_3403),.q(G176_26));
  bfr _b_1977(.a(_w_3402),.q(_w_3403));
  bfr _b_5425(.a(_w_6850),.q(_w_6851));
  spl4L G172_s_0(.a(_w_6975),.q0(_w_4240),.q1(G172_1),.q2(_w_4242),.q3(_w_4244));
  bfr _b_6137(.a(G4),.q(_w_7563));
  bfr _b_1975(.a(_w_3400),.q(_w_3401));
  bfr _b_1974(.a(_w_3399),.q(_w_3400));
  bfr _b_1972(.a(_w_3397),.q(_w_3398));
  bfr _b_1970(.a(_w_3395),.q(_w_3396));
  bfr _b_1969(.a(_w_3394),.q(_w_3395));
  bfr _b_1967(.a(_w_3392),.q(_w_3393));
  bfr _b_1966(.a(_w_3391),.q(_w_3392));
  spl4L g425_s_0(.a(n425),.q0(n425_0),.q1(n425_1),.q2(_w_3690),.q3(_w_3704));
  bfr _b_3559(.a(_w_4984),.q(n594_1));
  bfr _b_4517(.a(_w_5942),.q(_w_5943));
  bfr _b_7460(.a(_w_8885),.q(_w_8886));
  bfr _b_1964(.a(_w_3389),.q(G176_30));
  bfr _b_5283(.a(_w_6708),.q(_w_6709));
  bfr _b_1960(.a(_w_3385),.q(_w_3386));
  bfr _b_1957(.a(_w_3382),.q(_w_3383));
  bfr _b_2022(.a(_w_3447),.q(G139_4));
  bfr _b_1954(.a(_w_3379),.q(_w_3380));
  bfr _b_2716(.a(_w_4141),.q(_w_4142));
  bfr _b_4607(.a(_w_6032),.q(n879));
  bfr _b_1950(.a(_w_3375),.q(_w_3376));
  bfr _b_1949(.a(_w_3374),.q(G90_3));
  and_bb g1080(.a(G39_1),.b(n630_9),.q(n1080));
  bfr _b_6804(.a(_w_8229),.q(_w_8230));
  bfr _b_1946(.a(_w_3371),.q(n959_1));
  bfr _b_1962(.a(_w_3387),.q(_w_3388));
  bfr _b_1945(.a(_w_3370),.q(n386_4));
  bfr _b_1939(.a(_w_3364),.q(G147_4));
  or_bb g1327(.a(n403_2),.b(n542_5),.q(_w_4307));
  bfr _b_6077(.a(_w_7502),.q(_w_7503));
  bfr _b_5410(.a(_w_6835),.q(_w_6836));
  spl4L G166_s_0(.a(G166),.q0(_w_5836),.q1(G166_1),.q2(G166_2),.q3(G166_3));
  spl3L G147_s_1(.a(G147_3),.q0(_w_3364),.q1(G147_5),.q2(G147_6));
  bfr _b_5744(.a(_w_7169),.q(_w_7170));
  and_bi g201(.a(_w_7445),.b(G163_9),.q(_w_4980));
  bfr _b_2954(.a(_w_4379),.q(_w_4380));
  bfr _b_3344(.a(_w_4769),.q(_w_4770));
  spl4L G147_s_0(.a(_w_6559),.q0(G147_0),.q1(G147_1),.q2(_w_3367),.q3(G147_3));
  and_bb g470(.a(G115_2),.b(G123_10),.q(n470));
  bfr _b_2311(.a(_w_3736),.q(_w_3737));
  and_bi g301(.a(n299),.b(n300),.q(n301));
  bfr _b_3879(.a(_w_5304),.q(_w_5305));
  bfr _b_4480(.a(_w_5905),.q(_w_5906));
  spl3L g959_s_0(.a(n959),.q0(n959_0),.q1(_w_3371),.q2(_w_3372));
  and_bi g770(.a(n763_0),.b(n769_0),.q(n770));
  spl4L G102_s_4(.a(G102_3),.q0(G102_15),.q1(G102_16),.q2(G102_17),.q3(G102_18));
  spl4L G176_s_12(.a(G176_18),.q0(G176_46),.q1(_w_3375),.q2(G176_48),.q3(_w_3379));
  spl4L G176_s_10(.a(G176_16),.q0(G176_38),.q1(G176_39),.q2(G176_40),.q3(_w_3381));
  bfr _b_6896(.a(_w_8321),.q(_w_8322));
  and_bi g487(.a(G119_7),.b(G117_7),.q(n487));
  spl4L G176_s_9(.a(G176_15),.q0(G176_34),.q1(G176_35),.q2(G176_36),.q3(G176_37));
  spl4L G176_s_8(.a(G176_14),.q0(_w_3384),.q1(G176_31),.q2(_w_3390),.q3(G176_33));
  bfr _b_2001(.a(_w_3426),.q(_w_3427));
  and_bi g461(.a(_w_6425),.b(G123_13),.q(_w_4677));
  bfr _b_4962(.a(_w_6387),.q(_w_6388));
  and_bi g1202(.a(n1187_0),.b(n1201_0),.q(n1202));
  spl4L G176_s_0(.a(_w_7089),.q0(_w_3439),.q1(_w_3440),.q2(G176_2),.q3(G176_3));
  bfr _b_3555(.a(_w_4980),.q(_w_4981));
  spl4L G142_s_0(.a(_w_6531),.q0(G142_0),.q1(G142_1),.q2(_w_3441),.q3(_w_3442));
  spl2 g722_s_0(.a(n722),.q0(n722_0),.q1(n722_1));
  bfr _b_2529(.a(_w_3954),.q(_w_3955));
  bfr _b_3793(.a(_w_5218),.q(_w_5219));
  bfr _b_6671(.a(_w_8096),.q(_w_8097));
  bfr _b_2314(.a(_w_3739),.q(_w_3740));
  bfr _b_2341(.a(_w_3766),.q(_w_3767));
  bfr _b_7551(.a(_w_8976),.q(_w_8977));
  bfr _b_3938(.a(_w_5363),.q(_w_5364));
  spl2 g1244_s_0(.a(n1244),.q0(n1244_0),.q1(n1244_1));
  bfr _b_6799(.a(G67),.q(_w_8225));
  spl4L g815_s_2(.a(n815_3),.q0(n815_8),.q1(n815_9),.q2(n815_10),.q3(n815_11));
  bfr _b_5140(.a(_w_6565),.q(_w_6563));
  bfr _b_2302(.a(_w_3727),.q(G173_18));
  bfr _b_2036(.a(_w_3461),.q(_w_3462));
  spl3L g224_s_0(.a(n224),.q0(n224_0),.q1(_w_5579),.q2(n224_2));
  bfr _b_4526(.a(_w_5951),.q(_w_5952));
  spl4L g804_s_1(.a(n804_2),.q0(n804_4),.q1(n804_5),.q2(n804_6),.q3(n804_7));
  bfr _b_7429(.a(_w_8854),.q(_w_8855));
  and_bi g1282(.a(n1281),.b(n1280),.q(_w_4735));
  bfr _b_4880(.a(_w_6305),.q(n1285));
  spl4L g802_s_2(.a(n802_3),.q0(n802_8),.q1(n802_9),.q2(n802_10),.q3(n802_11));
  or_bb g1099(.a(n1095),.b(n1098),.q(n1099));
  spl4L g802_s_0(.a(n802),.q0(n802_0),.q1(n802_1),.q2(n802_2),.q3(n802_3));
  bfr _b_4447(.a(_w_5872),.q(_w_5873));
  spl2 g527_s_0(.a(n527),.q0(n527_0),.q1(n527_1));
  bfr _b_2538(.a(_w_3963),.q(_w_3964));
  bfr _b_5941(.a(_w_7366),.q(_w_7367));
  bfr _b_4054(.a(_w_5479),.q(_w_5480));
  spl4L g773_s_0(.a(n773),.q0(n773_0),.q1(n773_1),.q2(n773_2),.q3(n773_3));
  bfr _b_6235(.a(_w_7660),.q(_w_7628));
  bfr _b_2580(.a(_w_4005),.q(_w_4006));
  bfr _b_5463(.a(_w_6888),.q(_w_6889));
  bfr _b_2107(.a(_w_3532),.q(_w_3533));
  spl2 g707_s_0(.a(n707),.q0(n707_0),.q1(n707_1));
  bfr _b_2514(.a(_w_3939),.q(G88_0));
  spl4L g686_s_0(.a(n686),.q0(n686_0),.q1(n686_1),.q2(n686_2),.q3(n686_3));
  or_bb g512(.a(n510),.b(n511),.q(n512));
  bfr _b_6559(.a(_w_7984),.q(_w_7985));
  spl2 g488_s_0(.a(n488),.q0(n488_0),.q1(n488_1));
  bfr _b_6543(.a(_w_7968),.q(_w_7969));
  spl4L g1015_s_0(.a(G5291_0),.q0(_w_4232),.q1(G5291_1),.q2(G5291_2),.q3(G5291_3));
  bfr _b_2904(.a(_w_4329),.q(_w_4330));
  spl2 g670_s_0(.a(n670),.q0(n670_0),.q1(n670_1));
  spl2 g617_s_0(.a(n617),.q0(n617_0),.q1(n617_1));
  bfr _b_3092(.a(_w_4517),.q(_w_4518));
  spl4L g607_s_0(.a(n607),.q0(n607_0),.q1(n607_1),.q2(n607_2),.q3(n607_3));
  and_bi g1146(.a(G160_10),.b(G5286_5),.q(_w_6301));
  bfr _b_2086(.a(_w_3511),.q(G109_0));
  bfr _b_2455(.a(_w_3880),.q(_w_3881));
  bfr _b_4463(.a(_w_5888),.q(_w_5889));
  spl4L g588_s_1(.a(n588_2),.q0(n588_4),.q1(n588_5),.q2(n588_6),.q3(n588_7));
  spl2 g665_s_0(.a(n665),.q0(n665_0),.q1(n665_1));
  bfr _b_6721(.a(_w_8146),.q(_w_8134));
  spl2 g542_s_1(.a(n542_3),.q0(n542_4),.q1(n542_5));
  bfr _b_7338(.a(_w_8763),.q(_w_8764));
  spl4L g586_s_0(.a(n586),.q0(n586_0),.q1(n586_1),.q2(n586_2),.q3(n586_3));
  spl2 g524_s_0(.a(n524),.q0(n524_0),.q1(n524_1));
  bfr _b_6139(.a(_w_7564),.q(_w_7565));
  spl2 G74_s_0(.a(_w_8468),.q0(G74_0),.q1(G74_1));
  bfr _b_7426(.a(_w_8851),.q(_w_8852));
  spl2 g518_s_0(.a(n518),.q0(n518_0),.q1(n518_1));
  and_bi g375(.a(n374_0),.b(n373_0),.q(_w_5667));
  bfr _b_3094(.a(_w_4519),.q(_w_4520));
  spl4L G94_s_2(.a(G94_2),.q0(G94_6),.q1(G94_7),.q2(G94_8),.q3(G94_9));
  bfr _b_6800(.a(_w_8225),.q(_w_8226));
  bfr _b_3327(.a(_w_4752),.q(_w_4753));
  spl4L G64_s_6(.a(G64_18),.q0(G64_22),.q1(G64_23),.q2(G64_24),.q3(G64_25));
  spl4L G64_s_3(.a(G64_2),.q0(G64_12),.q1(G64_13),.q2(G64_14),.q3(_w_3445));
  spl4L G64_s_1(.a(G64_0),.q0(G64_4),.q1(G64_5),.q2(G64_6),.q3(G64_7));
  bfr _b_2578(.a(_w_4003),.q(_w_4004));
  spl2 g625_s_1(.a(G5255_3),.q0(G5255_4),.q1(G5255_5));
  spl2 g728_s_0(.a(n728),.q0(n728_0),.q1(n728_1));
  bfr _b_4039(.a(_w_5464),.q(_w_5465));
  spl3L G139_s_1(.a(G139_3),.q0(_w_3447),.q1(G139_5),.q2(G139_6));
  bfr _b_3690(.a(_w_5115),.q(_w_5116));
  bfr _b_2174(.a(_w_3599),.q(_w_3600));
  bfr _b_5027(.a(_w_6452),.q(_w_6453));
  spl4L G139_s_0(.a(_w_6490),.q0(G139_0),.q1(G139_1),.q2(_w_3448),.q3(G139_3));
  bfr _b_3576(.a(_w_5001),.q(_w_5002));
  bfr _b_5024(.a(_w_6449),.q(_w_6450));
  bfr _b_5349(.a(_w_6774),.q(_w_6775));
  spl2 g474_s_0(.a(n474),.q0(n474_0),.q1(n474_1));
  bfr _b_2097(.a(_w_3522),.q(G121_0));
  and_bi g192(.a(_w_7456),.b(G163_6),.q(n192));
  and_bi g939(.a(G160_17),.b(G5255_5),.q(n939));
  bfr _b_5490(.a(G164),.q(_w_6915));
  spl4L G115_s_0(.a(_w_6413),.q0(_w_6188),.q1(G115_1),.q2(G115_2),.q3(G115_3));
  bfr _b_5763(.a(_w_7188),.q(_w_7189));
  bfr _b_3364(.a(_w_4789),.q(_w_4790));
  bfr _b_3936(.a(_w_5361),.q(_w_5362));
  spl2 g1334_s_0(.a(n1334),.q0(n1334_0),.q1(n1334_1));
  bfr _b_2453(.a(_w_3878),.q(_w_3879));
  bfr _b_2152(.a(_w_3577),.q(_w_3578));
  bfr _b_6647(.a(_w_8072),.q(_w_8073));
  bfr _b_4878(.a(_w_6303),.q(_w_6304));
  bfr _b_4709(.a(_w_6134),.q(_w_6135));
  bfr _b_5068(.a(G14),.q(_w_6494));
  bfr _b_5146(.a(_w_6571),.q(_w_6572));
  bfr _b_2287(.a(_w_3712),.q(_w_3713));
  spl2 g683_s_1(.a(G5260_3),.q0(G5260_4),.q1(G5260_5));
  bfr _b_4178(.a(_w_5603),.q(_w_5604));
  spl4L g683_s_0(.a(G5260_0),.q0(_w_3491),.q1(G5260_1),.q2(G5260_2),.q3(G5260_3));
  and_bi g200(.a(G66_1),.b(n199),.q(_w_5152));
  spl2 g450_s_0(.a(n450),.q0(n450_0),.q1(n450_1));
  and_bi g345(.a(n344),.b(G142_1),.q(n345));
  bfr _b_7290(.a(_w_8715),.q(_w_8716));
  bfr _b_3682(.a(_w_5107),.q(_w_5108));
  bfr _b_6420(.a(_w_7845),.q(_w_7846));
  bfr _b_4539(.a(_w_5964),.q(_w_5965));
  bfr _b_5064(.a(_w_6489),.q(_w_6487));
  bfr _b_2269(.a(_w_3694),.q(_w_3695));
  spl4L g443_s_0(.a(n443),.q0(n443_0),.q1(_w_3499),.q2(n443_2),.q3(_w_3500));
  spl4L G100_s_2(.a(G100_1),.q0(G100_8),.q1(G100_9),.q2(G100_10),.q3(G100_11));
  bfr _b_5521(.a(_w_6946),.q(_w_6947));
  spl4L g346_s_0(.a(n346),.q0(n346_0),.q1(_w_3906),.q2(n346_2),.q3(n346_3));
  bfr _b_2327(.a(_w_3752),.q(G175_3));
  bfr _b_6673(.a(_w_8098),.q(_w_8099));
  and_bi g291(.a(G90_4),.b(G168_7),.q(n291));
  bfr _b_5428(.a(_w_6853),.q(_w_6854));
  bfr _b_3518(.a(_w_4943),.q(_w_4944));
  spl4L G100_s_1(.a(G100_0),.q0(G100_4),.q1(G100_5),.q2(G100_6),.q3(G100_7));
  bfr _b_4833(.a(_w_6258),.q(_w_6259));
  spl4L G101_s_4(.a(G101_3),.q0(G101_16),.q1(G101_17),.q2(G101_18),.q3(G101_19));
  spl2 G72_s_0(.a(_w_8400),.q0(G72_0),.q1(G72_1));
  spl4L G101_s_2(.a(G101_1),.q0(G101_8),.q1(G101_9),.q2(G101_10),.q3(G101_11));
  bfr _b_4141(.a(_w_5566),.q(_w_5567));
  bfr _b_4543(.a(_w_5968),.q(_w_5969));
  spl4L G101_s_0(.a(_w_6394),.q0(G101_0),.q1(G101_1),.q2(G101_2),.q3(G101_3));
  bfr _b_5979(.a(_w_7404),.q(_w_7405));
  spl4L g435_s_0(.a(n435),.q0(_w_4225),.q1(_w_4226),.q2(_w_4229),.q3(n435_3));
  spl4L G103_s_3(.a(G103_3),.q0(G103_10),.q1(G103_11),.q2(G103_12),.q3(G103_13));
  bfr _b_6677(.a(_w_8102),.q(_w_8103));
  bfr _b_6514(.a(G53),.q(_w_7940));
  bfr _b_6256(.a(_w_7681),.q(_w_7682));
  bfr _b_3000(.a(_w_4425),.q(_w_4426));
  bfr _b_4717(.a(_w_6142),.q(_w_6143));
  bfr _b_5476(.a(_w_6901),.q(_w_6902));
  bfr _b_2012(.a(_w_3437),.q(_w_3438));
  spl2 G96_s_1(.a(G96_1),.q0(G96_4),.q1(G96_5));
  spl3L G140_s_1(.a(G140_3),.q0(G140_4),.q1(G140_5),.q2(G140_6));
  bfr _b_3489(.a(_w_4914),.q(_w_4915));
  bfr _b_6411(.a(_w_7836),.q(_w_7837));
  spl4L G140_s_0(.a(_w_6525),.q0(G140_0),.q1(G140_1),.q2(_w_3510),.q3(G140_3));
  bfr _b_3509(.a(_w_4934),.q(_w_4935));
  bfr _b_5997(.a(_w_7422),.q(_w_7423));
  bfr _b_2291(.a(_w_3716),.q(G5257));
  bfr _b_6871(.a(G69),.q(_w_8297));
  bfr _b_4284(.a(_w_5709),.q(_w_5710));
  bfr _b_6360(.a(_w_7785),.q(_w_7786));
  spl4L G105_s_3(.a(G105_3),.q0(G105_10),.q1(G105_11),.q2(G105_12),.q3(G105_13));
  and_bb g373(.a(G141_2),.b(n372_0),.q(_w_5257));
  bfr _b_4042(.a(_w_5467),.q(G174_6));
  bfr _b_6168(.a(_w_7593),.q(_w_7594));
  and_bi g1089(.a(G15_1),.b(n632_10),.q(n1089));
  bfr _b_2024(.a(_w_3449),.q(G139_2));
  spl2 g1192_s_0(.a(n1192),.q0(n1192_0),.q1(n1192_1));
  bfr _b_5072(.a(_w_6497),.q(_w_6498));
  bfr _b_2164(.a(_w_3589),.q(_w_3590));
  spl2 G78_s_0(.a(_w_8603),.q0(G78_0),.q1(G78_1));
  bfr _b_6218(.a(_w_7643),.q(_w_7644));
  bfr _b_5624(.a(_w_7049),.q(_w_7050));
  or_bb g902(.a(G158_20),.b(G5259_4),.q(n902));
  spl2 G90_s_1(.a(G90_1),.q0(G90_4),.q1(G90_5));
  spl4L G121_s_3(.a(G121_3),.q0(G121_10),.q1(G121_11),.q2(G121_12),.q3(G121_13));
  spl4L G121_s_2(.a(G121_2),.q0(G121_6),.q1(G121_7),.q2(_w_3516),.q3(_w_3519));
  or_bb g1084(.a(G174_8),.b(G5293_2),.q(_w_6276));
  bfr _b_2867(.a(_w_4292),.q(n1377));
  bfr _b_5604(.a(_w_7029),.q(_w_7030));
  bfr _b_1968(.a(_w_3393),.q(_w_3394));
  bfr _b_5656(.a(_w_7081),.q(_w_7082));
  bfr _b_2707(.a(_w_4132),.q(n408_1));
  spl4L G121_s_0(.a(G121),.q0(_w_3522),.q1(G121_1),.q2(G121_2),.q3(_w_3523));
  spl2 G16_s_0(.a(_w_6816),.q0(G16_0),.q1(G16_1));
  bfr _b_7284(.a(_w_8709),.q(_w_8710));
  bfr _b_5953(.a(_w_7378),.q(_w_7379));
  spl4L G124_s_6(.a(G124_19),.q0(G124_22),.q1(G124_23),.q2(G124_24),.q3(G124_25));
  spl4L g632_s_2(.a(n632_3),.q0(n632_8),.q1(n632_9),.q2(n632_10),.q3(n632_11));
  bfr _b_4353(.a(_w_5778),.q(_w_5779));
  and_bi g1213(.a(n253_3),.b(n1211_1),.q(n1213));
  bfr _b_7071(.a(_w_8496),.q(_w_8497));
  spl3L G125_s_0(.a(_w_6430),.q0(G125_0),.q1(G125_1),.q2(_w_3560));
  and_bb g1097(.a(G87_0),.b(n804_7),.q(n1097));
  spl4L g253_s_0(.a(n253),.q0(n253_0),.q1(_w_3595),.q2(n253_2),.q3(n253_3));
  bfr _b_6735(.a(_w_8160),.q(_w_8161));
  bfr _b_5561(.a(_w_6986),.q(_w_6987));
  and_bi g776(.a(n775),.b(n774),.q(n776));
  bfr _b_5562(.a(_w_6987),.q(_w_6988));
  spl3L g402_s_0(.a(n402),.q0(n402_0),.q1(n402_1),.q2(_w_3640));
  or_bb g398(.a(G137_2),.b(n397_0),.q(n398));
  bfr _b_4361(.a(_w_5786),.q(_w_5787));
  bfr _b_7267(.a(_w_8692),.q(_w_8693));
  spl4L G168_s_3(.a(G168_3),.q0(G168_10),.q1(G168_11),.q2(G168_12),.q3(G168_13));
  and_bi g1123(.a(G73_0),.b(n802_10),.q(n1123));
  spl4L G168_s_0(.a(G168),.q0(_w_3642),.q1(G168_1),.q2(G168_2),.q3(G168_3));
  spl4L g552_s_6(.a(n552_19),.q0(n552_22),.q1(n552_23),.q2(n552_24),.q3(n552_25));
  and_bi g427(.a(n426_0),.b(n425_0),.q(n427));
  bfr _b_3422(.a(_w_4847),.q(_w_4848));
  spl4L g552_s_4(.a(n552_3),.q0(n552_16),.q1(n552_17),.q2(n552_18),.q3(n552_19));
  bfr _b_3791(.a(_w_5216),.q(_w_5217));
  spl2 G73_s_0(.a(_w_8434),.q0(G73_0),.q1(G73_1));
  bfr _b_6316(.a(_w_7741),.q(_w_7742));
  bfr _b_3951(.a(_w_5376),.q(_w_5377));
  spl4L g552_s_2(.a(n552_1),.q0(n552_8),.q1(n552_9),.q2(n552_10),.q3(n552_11));
  spl4L g552_s_0(.a(n552),.q0(n552_0),.q1(n552_1),.q2(n552_2),.q3(n552_3));
  bfr _b_7098(.a(_w_8523),.q(_w_8524));
  spl4L g802_s_1(.a(n802_2),.q0(n802_4),.q1(n802_5),.q2(n802_6),.q3(n802_7));
  spl4L G135_s_0(.a(_w_6481),.q0(G135_0),.q1(G135_1),.q2(_w_3643),.q3(G135_3));
  bfr _b_2969(.a(_w_4394),.q(_w_4395));
  bfr _b_6672(.a(_w_8097),.q(_w_8098));
  spl2 g1332_s_0(.a(n1332),.q0(n1332_0),.q1(n1332_1));
  bfr _b_4451(.a(_w_5876),.q(_w_5877));
  bfr _b_2412(.a(_w_3837),.q(_w_3838));
  spl4L G141_s_0(.a(_w_6528),.q0(G141_0),.q1(G141_1),.q2(_w_3646),.q3(G141_3));
  bfr _b_3620(.a(_w_5045),.q(_w_5046));
  spl3L G143_s_1(.a(G143_3),.q0(G143_4),.q1(G143_5),.q2(G143_6));
  and_bi g1338(.a(n1337_0),.b(n1297_0),.q(_w_4305));
  bfr _b_2271(.a(_w_3696),.q(_w_3697));
  bfr _b_2934(.a(_w_4359),.q(_w_4360));
  bfr _b_3080(.a(_w_4505),.q(_w_4506));
  bfr _b_7156(.a(_w_8581),.q(_w_8582));
  bfr _b_2470(.a(_w_3895),.q(_w_3896));
  bfr _b_3308(.a(_w_4733),.q(n268));
  bfr _b_2119(.a(_w_3544),.q(_w_3545));
  bfr _b_5587(.a(_w_7012),.q(_w_7013));
  spl2 g512_s_0(.a(n512),.q0(n512_0),.q1(n512_1));
  spl4L G150_s_0(.a(_w_6599),.q0(G150_0),.q1(G150_1),.q2(_w_3649),.q3(G150_3));
  bfr _b_6667(.a(_w_8092),.q(_w_8093));
  bfr _b_2111(.a(_w_3536),.q(_w_3537));
  bfr _b_5087(.a(_w_6512),.q(_w_6513));
  bfr _b_2348(.a(_w_3773),.q(_w_3774));
  bfr _b_2871(.a(_w_4296),.q(n394_1));
  spl4L G159_s_3(.a(G159_3),.q0(G159_11),.q1(G159_12),.q2(G159_13),.q3(G159_14));
  bfr _b_4783(.a(_w_6208),.q(_w_6209));
  bfr _b_2201(.a(_w_3626),.q(_w_3627));
  spl3L g185_s_1(.a(G5221_2),.q0(G5221_4),.q1(G5221_5),.q2(G5221_6));
  bfr _b_6186(.a(_w_7611),.q(_w_7612));
  bfr _b_2687(.a(_w_4112),.q(n479_1));
  bfr _b_5547(.a(_w_6972),.q(_w_6973));
  spl2 G155_s_0(.a(_w_6672),.q0(G155_0),.q1(_w_3656));
  bfr _b_7549(.a(_w_8974),.q(_w_8975));
  bfr _b_2046(.a(_w_3471),.q(_w_3472));
  bfr _b_6237(.a(_w_7662),.q(_w_7663));
  spl4L G158_s_6(.a(G158_19),.q0(_w_3662),.q1(G158_25),.q2(G158_26),.q3(G158_27));
  bfr _b_2884(.a(_w_4309),.q(n1327));
  spl4L G158_s_3(.a(G158_2),.q0(G158_12),.q1(G158_13),.q2(G158_14),.q3(G158_15));
  bfr _b_2092(.a(_w_3517),.q(_w_3518));
  and_bi g870(.a(G175_8),.b(n869),.q(n870));
  bfr _b_5084(.a(_w_6509),.q(_w_6510));
  bfr _b_4996(.a(_w_6421),.q(_w_6419));
  spl2 g544_s_0(.a(n544),.q0(n544_0),.q1(_w_3677));
  and_bb g540(.a(n374_1),.b(n399_1),.q(n540));
  bfr _b_4437(.a(_w_5862),.q(_w_5863));
  bfr _b_6700(.a(_w_8125),.q(_w_8126));
  bfr _b_1976(.a(_w_3401),.q(_w_3402));
  spl2 g546_s_0(.a(n546),.q0(n546_0),.q1(n546_1));
  or_bb g806(.a(n803),.b(n805),.q(n806));
  spl2 g551_s_0(.a(G5245_0),.q0(G5245),.q1(G5247));
  bfr _b_4116(.a(_w_5541),.q(_w_5542));
  bfr _b_5222(.a(_w_6647),.q(_w_6648));
  bfr _b_2151(.a(_w_3576),.q(_w_3577));
  spl2 g990_s_1(.a(G5287_3),.q0(G5287_4),.q1(G5287_5));
  or_bb g327(.a(n322),.b(n326),.q(_w_4771));
  bfr _b_7562(.a(_w_8987),.q(_w_8956));
  bfr _b_4179(.a(_w_5604),.q(_w_5605));
  bfr _b_6776(.a(_w_8201),.q(_w_8202));
  spl2 g534_s_0(.a(n534),.q0(n534_0),.q1(n534_1));
  and_bi g1272(.a(n1271),.b(n1266),.q(n1272));
  bfr _b_3034(.a(_w_4459),.q(_w_4460));
  spl4L G117_s_1(.a(G117_3),.q0(G117_4),.q1(G117_5),.q2(G117_6),.q3(G117_7));
  spl4L g415_s_0(.a(n415),.q0(_w_4191),.q1(_w_4192),.q2(_w_4206),.q3(n415_3));
  spl2 g453_s_0(.a(n453),.q0(_w_3808),.q1(n453_1));
  bfr _b_6148(.a(_w_7573),.q(_w_7574));
  bfr _b_2701(.a(_w_4126),.q(_w_4127));
  bfr _b_2080(.a(_w_3505),.q(G103_3));
  spl4L G166_s_2(.a(G166_2),.q0(G166_7),.q1(G166_8),.q2(G166_9),.q3(G166_10));
  spl4L G167_s_0(.a(G167),.q0(_w_3717),.q1(G167_1),.q2(G167_2),.q3(G167_3));
  bfr _b_5115(.a(_w_6540),.q(_w_6538));
  or_bb g547(.a(n413_1),.b(n546_0),.q(n547));
  spl4L G177_s_3(.a(G177_2),.q0(G177_12),.q1(_w_3718),.q2(G177_14),.q3(G177_15));
  spl4L G172_s_3(.a(G172_3),.q0(G172_11),.q1(G172_12),.q2(G172_13),.q3(_w_3719));
  bfr _b_2326(.a(_w_3751),.q(_w_3752));
  spl4L G173_s_6(.a(G173_19),.q0(_w_3720),.q1(G173_25),.q2(G173_26),.q3(G173_27));
  bfr _b_5446(.a(_w_6871),.q(_w_6872));
  bfr _b_3487(.a(_w_4912),.q(_w_4913));
  bfr _b_5326(.a(_w_6751),.q(_w_6752));
  spl4L G173_s_3(.a(G173_2),.q0(G173_12),.q1(G173_13),.q2(G173_14),.q3(G173_15));
  bfr _b_7508(.a(_w_8933),.q(_w_8934));
  or_bb g290(.a(G169_8),.b(G90_0),.q(n290));
  spl4L G66_s_1(.a(G66_2),.q0(G66_3),.q1(G66_4),.q2(G66_5),.q3(G66_6));
  bfr _b_3537(.a(_w_4962),.q(_w_4963));
  spl4L G163_s_0(.a(G163),.q0(G163_0),.q1(G163_1),.q2(G163_2),.q3(G163_3));
  spl4L G173_s_2(.a(G173_1),.q0(G173_8),.q1(G173_9),.q2(G173_10),.q3(G173_11));
  spl2 G2_s_1(.a(G2_3),.q0(G2_4),.q1(G2_5));
  bfr _b_3920(.a(_w_5345),.q(_w_5346));
  bfr _b_2060(.a(_w_3485),.q(_w_3486));
  and_bi g1243(.a(n1242),.b(G149_6),.q(n1243));
  spl2 G24_s_0(.a(_w_7277),.q0(G24_0),.q1(G24_1));
  bfr _b_5606(.a(_w_7031),.q(_w_7004));
  bfr _b_2664(.a(_w_4089),.q(_w_4090));
  spl2 g421_s_1(.a(n421_3),.q0(n421_4),.q1(n421_5));
  spl2 G3_s_0(.a(_w_7413),.q0(G3_0),.q1(G3_1));
  bfr _b_3991(.a(_w_5416),.q(_w_5417));
  bfr _b_4191(.a(_w_5616),.q(_w_5617));
  bfr _b_2544(.a(_w_3969),.q(_w_3970));
  bfr _b_7277(.a(_w_8702),.q(_w_8703));
  bfr _b_6874(.a(_w_8299),.q(_w_8300));
  bfr _b_3896(.a(_w_5321),.q(_w_5322));
  spl4L G174_s_2(.a(G174_1),.q0(G174_8),.q1(G174_9),.q2(G174_10),.q3(G174_11));
  spl3L G175_s_1(.a(G175_1),.q0(G175_4),.q1(G175_5),.q2(_w_3745));
  spl2 g444_s_0(.a(n444),.q0(n444_0),.q1(n444_1));
  spl4L G94_s_0(.a(G94),.q0(_w_3488),.q1(G94_1),.q2(G94_2),.q3(_w_3489));
  spl4L G64_s_4(.a(G64_3),.q0(G64_15),.q1(G64_16),.q2(G64_17),.q3(G64_18));
  bfr _b_2095(.a(_w_3520),.q(_w_3521));
  spl2 G22_s_0(.a(_w_7212),.q0(G22_0),.q1(G22_1));
  spl4L G124_s_3(.a(G124_2),.q0(G124_12),.q1(G124_13),.q2(G124_14),.q3(G124_15));
  bfr _b_2021(.a(_w_3446),.q(G5214));
  spl2 g667_s_0(.a(n667),.q0(n667_0),.q1(n667_1));
  spl2 g194_s_0(.a(G5229_0),.q0(G5229),.q1(G5230));
  bfr _b_2474(.a(_w_3899),.q(_w_3900));
  bfr _b_4649(.a(_w_6074),.q(_w_6075));
  bfr _b_6392(.a(_w_7817),.q(_w_7818));
  spl2 g550_s_0(.a(G5244_0),.q0(G5244),.q1(G5246));
  bfr _b_2746(.a(_w_4171),.q(_w_4172));
  bfr _b_4123(.a(_w_5548),.q(_w_5549));
  spl2 g400_s_1(.a(n400_3),.q0(_w_3788),.q1(n400_5));
  bfr _b_5665(.a(_w_7090),.q(_w_7091));
  bfr _b_2347(.a(_w_3772),.q(_w_3773));
  bfr _b_2377(.a(_w_3802),.q(_w_3803));
  spl4L g1027_s_0(.a(G5293_0),.q0(_w_3794),.q1(G5293_1),.q2(G5293_2),.q3(G5293_3));
  bfr _b_3245(.a(_w_4670),.q(_w_4671));
  spl3L g375_s_1(.a(n375_3),.q0(_w_3802),.q1(n375_5),.q2(n375_6));
  or_bb g591(.a(n585),.b(n590),.q(_w_5451));
  bfr _b_6980(.a(_w_8405),.q(_w_8406));
  spl4L g375_s_0(.a(n375),.q0(_w_3804),.q1(n375_1),.q2(_w_3805),.q3(n375_3));
  and_bi g1081(.a(G40_1),.b(n632_9),.q(n1081));
  bfr _b_4559(.a(_w_5984),.q(_w_5985));
  or_bb g986(.a(G176_9),.b(n779_1),.q(n986));
  bfr _b_4392(.a(_w_5817),.q(_w_5818));
  spl4L g630_s_2(.a(n630_3),.q0(n630_8),.q1(n630_9),.q2(n630_10),.q3(n630_11));
  bfr _b_2759(.a(_w_4184),.q(_w_4185));
  bfr _b_3005(.a(_w_4430),.q(_w_4431));
  bfr _b_3883(.a(_w_5308),.q(_w_5309));
  spl4L G98_s_4(.a(G98_3),.q0(G98_16),.q1(G98_17),.q2(G98_18),.q3(G98_19));
  bfr _b_6215(.a(_w_7640),.q(_w_7641));
  bfr _b_2304(.a(_w_3729),.q(_w_3730));
  spl3L G114_s_0(.a(_w_6411),.q0(_w_3816),.q1(G114_0),.q2(_w_3853));
  spl4L g421_s_0(.a(n421),.q0(n421_0),.q1(_w_3607),.q2(_w_3622),.q3(_w_3637));
  spl2 G40_s_0(.a(_w_7595),.q0(G40_0),.q1(G40_1));
  spl2 G54_s_0(.a(_w_7961),.q0(G54_0),.q1(_w_3897));
  bfr _b_2730(.a(_w_4155),.q(_w_4156));
  bfr _b_5261(.a(_w_6686),.q(_w_6687));
  bfr _b_3543(.a(_w_4968),.q(_w_4969));
  bfr _b_4310(.a(_w_5735),.q(_w_5736));
  spl4L G64_s_0(.a(_w_8148),.q0(_w_3651),.q1(G64_1),.q2(G64_2),.q3(G64_3));
  spl3L g469_s_1(.a(n469_2),.q0(n469_4),.q1(n469_5),.q2(n469_6));
  bfr _b_3890(.a(_w_5315),.q(_w_5316));
  bfr _b_3458(.a(_w_4883),.q(_w_4884));
  bfr _b_3769(.a(_w_5194),.q(_w_5195));
  bfr _b_2909(.a(_w_4334),.q(_w_4335));
  bfr _b_1948(.a(_w_3373),.q(G90_0));
  spl2 g463_s_1(.a(n463_3),.q0(n463_4),.q1(n463_5));
  bfr _b_1953(.a(_w_3378),.q(G176_47));
  spl2 g234_s_0(.a(n234),.q0(_w_3923),.q1(n234_1));
  bfr _b_2123(.a(_w_3548),.q(_w_3549));
  or_bb g488(.a(n486),.b(n487),.q(n488));
  spl3L g249_s_0(.a(n249),.q0(n249_0),.q1(_w_3926),.q2(n249_2));
  and_bb g279(.a(n259),.b(n278),.q(n279));
  bfr _b_2822(.a(_w_4247),.q(_w_4248));
  bfr _b_2099(.a(_w_3524),.q(_w_3525));
  bfr _b_2103(.a(_w_3528),.q(_w_3529));
  bfr _b_2689(.a(_w_4114),.q(_w_4115));
  spl4L G123_s_2(.a(G123_1),.q0(G123_8),.q1(G123_9),.q2(_w_3931),.q3(_w_3932));
  and_bi g1096(.a(G77_0),.b(n802_7),.q(n1096));
  bfr _b_6088(.a(_w_7513),.q(_w_7514));
  spl4L G123_s_1(.a(G123_0),.q0(_w_3933),.q1(G123_5),.q2(G123_6),.q3(G123_7));
  spl4L G123_s_0(.a(G123),.q0(G123_0),.q1(G123_1),.q2(_w_3935),.q3(G123_3));
  bfr _b_6970(.a(_w_8395),.q(_w_8396));
  spl2 g373_s_0(.a(n373),.q0(n373_0),.q1(n373_1));
  bfr _b_2130(.a(_w_3555),.q(_w_3556));
  bfr _b_3721(.a(_w_5146),.q(_w_5147));
  bfr _b_1973(.a(_w_3398),.q(G176_32));
  bfr _b_4551(.a(_w_5976),.q(_w_5977));
  bfr _b_6956(.a(_w_8381),.q(_w_8382));
  bfr _b_6010(.a(_w_7435),.q(_w_7436));
  bfr _b_4794(.a(_w_6219),.q(_w_6220));
  bfr _b_4332(.a(_w_5757),.q(n233_1));
  spl2 g1187_s_0(.a(n1187),.q0(n1187_0),.q1(n1187_1));
  bfr _b_6765(.a(_w_8190),.q(_w_8191));
  bfr _b_3683(.a(_w_5108),.q(_w_5109));
  bfr _b_6635(.a(_w_8060),.q(_w_8061));
  bfr _b_2198(.a(_w_3623),.q(_w_3624));
  spl2 G87_s_0(.a(_w_8908),.q0(G87_0),.q1(G87_1));
  bfr _b_4986(.a(G114),.q(_w_6412));
  spl4L G88_s_0(.a(G88),.q0(_w_3938),.q1(_w_3940),.q2(_w_3942),.q3(G88_3));
  and_bi g1104(.a(n1103),.b(n1101),.q(_w_6286));
  spl4L G92_s_3(.a(G92_3),.q0(G92_10),.q1(G92_11),.q2(G92_12),.q3(G92_13));
  and_bi g552(.a(G176_44),.b(G177_16),.q(n552));
  spl3L g744_s_1(.a(n744_3),.q0(n744_4),.q1(n744_5),.q2(n744_6));
  bfr _b_5506(.a(_w_6931),.q(_w_6932));
  bfr _b_4004(.a(_w_5429),.q(_w_5430));
  bfr _b_4433(.a(_w_5858),.q(_w_5859));
  spl2 G25_s_0(.a(_w_7310),.q0(G25_0),.q1(G25_1));
  spl4L G96_s_2(.a(G96_2),.q0(G96_6),.q1(G96_7),.q2(G96_8),.q3(G96_9));
  spl3L g399_s_0(.a(n399),.q0(n399_0),.q1(n399_1),.q2(_w_3946));
  bfr _b_7474(.a(_w_8899),.q(_w_8900));
  spl2 g184_s_0(.a(G5213_0),.q0(_w_3952),.q1(G5213_1));
  spl4L G169_s_3(.a(G169_3),.q0(G169_11),.q1(G169_12),.q2(G169_13),.q3(G169_14));
  or_bb g617(.a(n443_3),.b(n445_2),.q(n617));
  and_bi g1014(.a(n1013),.b(n1011),.q(n1014));
  bfr _b_3988(.a(_w_5413),.q(_w_5414));
  spl3L G169_s_1(.a(G169_1),.q0(G169_4),.q1(G169_5),.q2(G169_6));
  spl2 g494_s_0(.a(n494),.q0(n494_0),.q1(n494_1));
  and_bi g263(.a(G147_0),.b(n262),.q(n263));
  spl2 g179_s_0(.a(G5199_0),.q0(_w_3958),.q1(G5199_1));
  bfr _b_4153(.a(_w_5578),.q(n679));
  bfr _b_6633(.a(G59),.q(_w_8059));
  spl4L G167_s_2(.a(G167_2),.q0(G167_6),.q1(G167_7),.q2(G167_8),.q3(G167_9));
  bfr _b_3649(.a(_w_5074),.q(_w_5075));
  spl2 g1377_s_0(.a(n1377),.q0(n1377_0),.q1(n1377_1));
  spl2 g392_s_0(.a(n392),.q0(n392_0),.q1(n392_1));
  spl4L G103_s_0(.a(G103),.q0(_w_3504),.q1(G103_1),.q2(G103_2),.q3(_w_3505));
  bfr _b_2227(.a(_w_3652),.q(G5217));
  bfr _b_4788(.a(_w_6213),.q(_w_6214));
  spl4L G158_s_2(.a(G158_1),.q0(G158_8),.q1(G158_9),.q2(G158_10),.q3(G158_11));
  bfr _b_2900(.a(_w_4325),.q(_w_4326));
  spl2 g743_s_0(.a(G5262_0),.q0(_w_3973),.q1(G5262_1));
  bfr _b_6948(.a(_w_8373),.q(_w_8374));
  bfr _b_2105(.a(_w_3530),.q(_w_3531));
  bfr _b_3783(.a(_w_5208),.q(_w_5209));
  bfr _b_2519(.a(_w_3944),.q(G92_0));
  spl2 g394_s_1(.a(n394_3),.q0(_w_3974),.q1(n394_5));
  and_bb g1022(.a(_w_7715),.b(n552_7),.q(_w_6199));
  bfr _b_4113(.a(_w_5538),.q(_w_5539));
  spl4L g442_s_1(.a(n442_3),.q0(_w_4002),.q1(n442_5),.q2(n442_6),.q3(n442_7));
  bfr _b_2811(.a(_w_4236),.q(_w_4237));
  spl2 g1204_s_0(.a(n1204),.q0(n1204_0),.q1(n1204_1));
  spl2 g506_s_0(.a(G5242_0),.q0(_w_4003),.q1(G5242_1));
  spl2 g533_s_0(.a(G5243_0),.q0(_w_4007),.q1(G5243_1));
  spl4L G109_s_3(.a(G109_3),.q0(G109_10),.q1(G109_11),.q2(G109_12),.q3(G109_13));
  bfr _b_2743(.a(_w_4168),.q(_w_4169));
  bfr _b_2053(.a(_w_3478),.q(_w_3479));
  bfr _b_5459(.a(_w_6884),.q(_w_6885));
  spl2 g615_s_1(.a(G5254_3),.q0(G5254_4),.q1(G5254_5));
  bfr _b_4965(.a(_w_6390),.q(_w_6354));
  spl4L g439_s_0(.a(n439),.q0(_w_4782),.q1(n439_1),.q2(_w_4783),.q3(n439_3));
  bfr _b_5788(.a(_w_7213),.q(_w_7214));
  bfr _b_2239(.a(_w_3664),.q(G158_20));
  spl4L G176_s_1(.a(G176_0),.q0(_w_3421),.q1(G176_5),.q2(G176_6),.q3(_w_3430));
  spl4L G149_s_0(.a(_w_6563),.q0(G149_0),.q1(G149_1),.q2(_w_4063),.q3(G149_3));
  bfr _b_4627(.a(_w_6052),.q(n1047));
  spl2 g978_s_1(.a(G5285_3),.q0(G5285_4),.q1(G5285_5));
  bfr _b_3582(.a(_w_5007),.q(_w_5008));
  spl2 g996_s_1(.a(G5288_3),.q0(G5288_4),.q1(G5288_5));
  bfr _b_5626(.a(_w_7051),.q(_w_7052));
  bfr _b_3820(.a(_w_5245),.q(_w_5246));
  spl4L g246_s_0(.a(n246),.q0(n246_0),.q1(n246_1),.q2(_w_4101),.q3(n246_3));
  spl2 g521_s_0(.a(n521),.q0(n521_0),.q1(n521_1));
  spl2 g451_s_1(.a(n451_3),.q0(n451_4),.q1(n451_5));
  bfr _b_7214(.a(_w_8639),.q(_w_8640));
  spl3L g653_s_0(.a(n653),.q0(n653_0),.q1(n653_1),.q2(n653_2));
  bfr _b_7547(.a(_w_8972),.q(_w_8973));
  bfr _b_2337(.a(_w_3762),.q(_w_3763));
  bfr _b_4345(.a(_w_5770),.q(_w_5771));
  spl2 g256_s_0(.a(n256),.q0(n256_0),.q1(_w_4081));
  bfr _b_7285(.a(_w_8710),.q(_w_8711));
  or_bb g1107(.a(n1105),.b(n1106),.q(n1107));
  spl2 G71_s_0(.a(_w_8366),.q0(G71_0),.q1(G71_1));
  bfr _b_4095(.a(_w_5520),.q(_w_5521));
  spl4L g378_s_0(.a(n378),.q0(n378_0),.q1(n378_1),.q2(n378_2),.q3(n378_3));
  spl4L g1021_s_0(.a(G5292_0),.q0(_w_4093),.q1(G5292_1),.q2(G5292_2),.q3(G5292_3));
  or_bb g947(.a(G160_16),.b(G5258_5),.q(_w_6275));
  bfr _b_3540(.a(_w_4965),.q(_w_4966));
  bfr _b_6942(.a(_w_8367),.q(_w_8368));
  bfr _b_1940(.a(_w_3365),.q(_w_3366));
  bfr _b_3898(.a(_w_5323),.q(_w_5324));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(n250_1));
  spl2 g479_s_1(.a(n479_3),.q0(n479_4),.q1(n479_5));
  bfr _b_2862(.a(_w_4287),.q(G176_20));
  bfr _b_7159(.a(_w_8584),.q(_w_8585));
  bfr _b_3569(.a(_w_4994),.q(_w_4995));
  bfr _b_2070(.a(_w_3495),.q(_w_3496));
  bfr _b_6004(.a(_w_7429),.q(_w_7430));
  spl2 g408_s_0(.a(n408),.q0(n408_0),.q1(_w_4126));
  and_bi g1446(.a(_w_7491),.b(G177_5),.q(_w_4831));
  bfr _b_2368(.a(_w_3793),.q(n400_4));
  bfr _b_2955(.a(_w_4380),.q(_w_4381));
  bfr _b_7272(.a(_w_8697),.q(_w_8698));
  bfr _b_6754(.a(_w_8179),.q(_w_8180));
  or_bb g715(.a(n391_3),.b(n397_3),.q(n715));
  bfr _b_2166(.a(_w_3591),.q(_w_3592));
  bfr _b_2015(.a(_w_3440),.q(G176_1));
  and_bi g1115(.a(G74_0),.b(n802_9),.q(n1115));
  spl3L g414_s_0(.a(n414),.q0(n414_0),.q1(_w_4134),.q2(_w_4137));
  spl4L G160_s_5(.a(G160_18),.q0(_w_4143),.q1(G160_21),.q2(_w_4144),.q3(G160_23));
  spl4L G160_s_3(.a(G160_2),.q0(G160_12),.q1(G160_13),.q2(G160_14),.q3(G160_15));
  spl4L G160_s_1(.a(G160_0),.q0(G160_4),.q1(G160_5),.q2(_w_4145),.q3(G160_7));
  bfr _b_2325(.a(_w_3750),.q(G175_2));
  or_bb g707(.a(n705),.b(n706),.q(n707));
  spl2 G105_s_1(.a(G105_1),.q0(G105_4),.q1(G105_5));
  spl4L g581_s_0(.a(G5251_0),.q0(_w_4148),.q1(G5251_1),.q2(G5251_2),.q3(G5251_3));
  spl2 g307_s_0(.a(n307),.q0(n307_0),.q1(_w_4171));
  and_bi g1451(.a(G23_0),.b(n588_11),.q(n1451));
  and_bi g1203(.a(n1201_1),.b(n1187_1),.q(n1203));
  bfr _b_3542(.a(_w_4967),.q(_w_4968));
  or_bb g1076(.a(G174_10),.b(G5292_2),.q(_w_5898));
  bfr _b_3295(.a(_w_4720),.q(_w_4721));
  bfr _b_6164(.a(_w_7589),.q(_w_7590));
  spl3L g434_s_0(.a(n434),.q0(n434_0),.q1(_w_4175),.q2(_w_4176));
  spl3L g380_s_0(.a(n380),.q0(n380_0),.q1(n380_1),.q2(_w_4181));
  bfr _b_3362(.a(_w_4787),.q(_w_4788));
  spl4L g387_s_0(.a(n387),.q0(n387_0),.q1(_w_4182),.q2(_w_4186),.q3(_w_4190));
  bfr _b_5189(.a(_w_6614),.q(_w_6615));
  spl3L g388_s_0(.a(n388),.q0(n388_0),.q1(n388_1),.q2(n388_2));
  spl4L g412_s_0(.a(n412),.q0(n412_0),.q1(n412_1),.q2(n412_2),.q3(n412_3));
  spl2 g701_s_0(.a(n701),.q0(n701_0),.q1(n701_1));
  spl2 g435_s_1(.a(n435_3),.q0(n435_4),.q1(n435_5));
  spl2 g1176_s_0(.a(n1176),.q0(n1176_0),.q1(n1176_1));
  bfr _b_5004(.a(_w_6429),.q(_w_6428));
  spl2 g1223_s_0(.a(n1223),.q0(n1223_0),.q1(n1223_1));
  bfr _b_3790(.a(_w_5215),.q(_w_5216));
  spl2 g1275_s_0(.a(n1275),.q0(n1275_0),.q1(n1275_1));
  bfr _b_3192(.a(_w_4617),.q(G5256));
  bfr _b_4875(.a(_w_6300),.q(n1140));
  bfr _b_5379(.a(_w_6804),.q(_w_6805));
  spl2 G5_s_0(.a(_w_7842),.q0(G5_0),.q1(G5_1));
  bfr _b_6983(.a(_w_8408),.q(_w_8409));
  spl2 g1292_s_0(.a(n1292),.q0(n1292_0),.q1(n1292_1));
  spl2 g1300_s_0(.a(n1300),.q0(n1300_0),.q1(n1300_1));
  spl2 g1305_s_0(.a(n1305),.q0(n1305_0),.q1(n1305_1));
  and_bi g182(.a(_w_8147),.b(G165_0),.q(_w_5540));
  bfr _b_2589(.a(_w_4014),.q(_w_4015));
  bfr _b_3719(.a(_w_5144),.q(_w_5145));
  spl2 g1359_s_0(.a(n1359),.q0(n1359_0),.q1(n1359_1));
  spl3L G138_s_1(.a(G138_3),.q0(_w_4246),.q1(G138_5),.q2(G138_6));
  bfr _b_2705(.a(_w_4130),.q(_w_4131));
  bfr _b_7030(.a(_w_8455),.q(_w_8456));
  bfr _b_6525(.a(_w_7950),.q(_w_7951));
  bfr _b_3965(.a(_w_5390),.q(_w_5391));
  spl4L G161_s_2(.a(G161_2),.q0(G161_7),.q1(G161_8),.q2(G161_9),.q3(G161_10));
  bfr _b_2294(.a(_w_3719),.q(G172_14));
  spl2 g1374_s_0(.a(n1374),.q0(n1374_0),.q1(n1374_1));
  and_bi g218(.a(n216),.b(n217),.q(_w_5477));
  spl2 g1386_s_0(.a(n1386),.q0(n1386_0),.q1(n1386_1));
  spl2 g1398_s_0(.a(n1398),.q0(n1398_0),.q1(n1398_1));
  bfr _b_5010(.a(_w_6435),.q(_w_6434));
  spl2 g547_s_0(.a(n547),.q0(n547_0),.q1(_w_4247));
  bfr _b_2159(.a(_w_3584),.q(_w_3585));
  spl3L G152_s_0(.a(_w_6602),.q0(_w_3652),.q1(_w_3653),.q2(G152_0));
  spl2 g1428_s_0(.a(n1428),.q0(n1428_0),.q1(n1428_1));
  bfr _b_4383(.a(_w_5808),.q(_w_5809));
  spl4L inv_G1_s_0(.a(i_G1),.q0(G5222),.q1(G5223),.q2(G5224),.q3(G5225));
  spl4L g1444_s_0(.a(n1444),.q0(n1444_0),.q1(n1444_1),.q2(n1444_2),.q3(n1444_3));
  and_bb g1071(.a(n1068),.b(n1070),.q(_w_5920));
  bfr _b_6523(.a(_w_7948),.q(_w_7949));
  spl2 inv_G114_s_0(.a(i_G114),.q0(G5226),.q1(G5227));
  bfr _b_6662(.a(_w_8087),.q(_w_8088));
  bfr _b_4523(.a(_w_5948),.q(n807));
  bfr _b_2059(.a(_w_3484),.q(_w_3485));
  spl3L inv_G151_s_0(.a(i_G151),.q0(G5196),.q1(G5201),.q2(G5202));
  bfr _b_2196(.a(_w_3621),.q(n421_1));
  bfr _b_2037(.a(_w_3462),.q(_w_3463));
  bfr _b_7346(.a(_w_8771),.q(_w_8772));
  bfr _b_4659(.a(_w_6084),.q(_w_6085));
  inv inv_G156(.a(G156_1),.q(G5208));
  spl2 G107_s_1(.a(G107_1),.q0(G107_4),.q1(G107_5));
  inv inv_G129(.a(G129_1),.q(G5204));
  bfr _b_2808(.a(_w_4233),.q(_w_4234));
  inv inv_G125(.a(G125_2),.q(G5203));
  bfr _b_2062(.a(_w_3487),.q(n459_2));
  and_bb g687(.a(n462_2),.b(n472_4),.q(n687));
  spl4L g773_s_1(.a(n773_3),.q0(n773_4),.q1(n773_5),.q2(n773_6),.q3(n773_7));
  spl2 g1314_s_0(.a(n1314),.q0(n1314_0),.q1(n1314_1));
  or_ii g1480(.a(G64_5),.b(n1479),.q(G5315));
  bfr _b_1961(.a(_w_3386),.q(_w_3387));
  and_bb g973(.a(G54_1),.b(n552_4),.q(n973));
  spl2 g695_s_0(.a(n695),.q0(n695_0),.q1(n695_1));
  bfr _b_3716(.a(_w_5141),.q(_w_5142));
  bfr _b_3550(.a(_w_4975),.q(n900));
  and_bb g1475(.a(n1472),.b(n1474),.q(n1475));
  bfr _b_2293(.a(_w_3718),.q(G177_13));
  bfr _b_5826(.a(_w_7251),.q(_w_7252));
  bfr _b_2167(.a(_w_3592),.q(_w_3593));
  and_bi g1474(.a(G161_14),.b(n1473),.q(_w_4253));
  or_bb g1472(.a(G160_6),.b(n1444_3),.q(n1472));
  bfr _b_4040(.a(_w_5465),.q(_w_5466));
  bfr _b_4031(.a(_w_5456),.q(_w_5457));
  or_bb g781(.a(n457_1),.b(n780),.q(_w_4621));
  bfr _b_6210(.a(_w_7635),.q(_w_7636));
  bfr _b_3815(.a(_w_5240),.q(_w_5241));
  bfr _b_2237(.a(_w_3662),.q(_w_3663));
  bfr _b_4475(.a(_w_5900),.q(_w_5901));
  bfr _b_2328(.a(_w_3753),.q(_w_3754));
  and_bi g1467(.a(G79_0),.b(n802_11),.q(n1467));
  bfr _b_7052(.a(_w_8477),.q(_w_8478));
  bfr _b_3720(.a(_w_5145),.q(n477_1));
  or_bb g1463(.a(G158_6),.b(n1444_2),.q(n1463));
  spl4L g451_s_0(.a(n451),.q0(n451_0),.q1(_w_5923),.q2(_w_5925),.q3(_w_5927));
  bfr _b_4779(.a(_w_6204),.q(_w_6205));
  and_bi g1459(.a(G23_1),.b(n632_11),.q(n1459));
  and_bb g1458(.a(n1455),.b(n1457),.q(n1458));
  bfr _b_6049(.a(_w_7474),.q(_w_7475));
  bfr _b_3824(.a(_w_5249),.q(G130_0));
  or_bb g1454(.a(n1450),.b(n1453),.q(_w_4256));
  spl4L G105_s_0(.a(G105),.q0(_w_4257),.q1(G105_1),.q2(G105_2),.q3(_w_4258));
  spl4L G161_s_0(.a(_w_6877),.q0(_w_4259),.q1(G161_1),.q2(_w_4261),.q3(_w_4263));
  bfr _b_5690(.a(_w_7115),.q(_w_7116));
  bfr _b_3861(.a(_w_5286),.q(_w_5287));
  and_bi g1448(.a(G173_5),.b(n1447_0),.q(n1448));
  bfr _b_6665(.a(_w_8090),.q(_w_8091));
  bfr _b_5862(.a(_w_7287),.q(_w_7288));
  bfr _b_4547(.a(_w_5972),.q(_w_5973));
  or_bb g1444(.a(n1440_1),.b(n1443),.q(n1444));
  bfr _b_6337(.a(_w_7762),.q(_w_7763));
  bfr _b_2160(.a(_w_3585),.q(_w_3586));
  bfr _b_6454(.a(_w_7879),.q(_w_7880));
  spl2 g429_s_0(.a(n429),.q0(n429_0),.q1(_w_4265));
  bfr _b_6755(.a(_w_8180),.q(_w_8181));
  and_bi g415(.a(n414_0),.b(n413_0),.q(n415));
  bfr _b_3231(.a(_w_4656),.q(_w_4657));
  bfr _b_3666(.a(_w_5091),.q(_w_5092));
  spl4L g418_s_0(.a(n418),.q0(n418_0),.q1(n418_1),.q2(n418_2),.q3(n418_3));
  bfr _b_4351(.a(_w_5776),.q(_w_5777));
  bfr _b_2250(.a(_w_3675),.q(_w_3676));
  and_bi g1437(.a(G176_33),.b(n1436),.q(n1437));
  and_bi g1435(.a(n1434_0),.b(n1377_0),.q(_w_4278));
  spl2 g1298_s_0(.a(n1298),.q0(n1298_0),.q1(n1298_1));
  bfr _b_6912(.a(_w_8337),.q(_w_8338));
  bfr _b_6465(.a(_w_7890),.q(_w_7891));
  or_bb g654(.a(G2_5),.b(n537_4),.q(n654));
  bfr _b_4422(.a(_w_5847),.q(_w_5848));
  or_bb g1431(.a(n1429),.b(n1430),.q(n1431));
  spl2 g466_s_0(.a(n466),.q0(n466_0),.q1(n466_1));
  and_bi g1430(.a(n1428_1),.b(n1407_1),.q(n1430));
  bfr _b_7512(.a(_w_8937),.q(_w_8938));
  bfr _b_2427(.a(_w_3852),.q(G5218));
  and_bi g1428(.a(n1427),.b(n1426),.q(n1428));
  and_bi g563(.a(n439_1),.b(n443_1),.q(n563));
  and_bi g1176(.a(n458_2),.b(n1175),.q(n1176));
  bfr _b_4760(.a(_w_6185),.q(_w_6186));
  or_bb g1427(.a(n1416_1),.b(n1425_1),.q(n1427));
  and_bi g270(.a(G126_4),.b(G168_5),.q(n270));
  bfr _b_4734(.a(_w_6159),.q(_w_6160));
  spl2 G176_s_5(.a(G176_11),.q0(_w_4282),.q1(G176_21));
  and_bi g1424(.a(n1423),.b(G137_6),.q(n1424));
  bfr _b_4052(.a(_w_5477),.q(_w_5478));
  spl4L G169_s_2(.a(G169_2),.q0(G169_7),.q1(G169_8),.q2(G169_9),.q3(G169_10));
  and_bb g1421(.a(G102_18),.b(G103_12),.q(n1421));
  bfr _b_4312(.a(_w_5737),.q(_w_5738));
  bfr _b_3415(.a(_w_4840),.q(_w_4841));
  spl2 g1288_s_0(.a(n1288),.q0(n1288_0),.q1(n1288_1));
  bfr _b_3061(.a(_w_4486),.q(_w_4487));
  bfr _b_2353(.a(_w_3778),.q(_w_3779));
  bfr _b_6538(.a(_w_7963),.q(_w_7964));
  bfr _b_3514(.a(_w_4939),.q(_w_4940));
  and_bi g1418(.a(G103_11),.b(G101_19),.q(n1418));
  spl2 g327_s_0(.a(n327),.q0(n327_0),.q1(n327_1));
  and_bi g881(.a(G25_1),.b(n632_6),.q(n881));
  or_bb g1417(.a(G100_5),.b(G103_10),.q(n1417));
  or_bb g1416(.a(n1411),.b(n1415),.q(n1416));
  spl2 g783_s_0(.a(n783),.q0(n783_0),.q1(n783_1));
  and_bi g1413(.a(G98_18),.b(G109_13),.q(n1413));
  and_bb g1412(.a(G102_17),.b(G109_12),.q(n1412));
  bfr _b_7499(.a(_w_8924),.q(_w_8925));
  spl4L g552_s_1(.a(n552_0),.q0(n552_4),.q1(n552_5),.q2(n552_6),.q3(n552_7));
  bfr _b_3341(.a(_w_4766),.q(_w_4767));
  bfr _b_6106(.a(_w_7531),.q(_w_7532));
  bfr _b_2660(.a(_w_4085),.q(_w_4086));
  bfr _b_4580(.a(_w_6005),.q(_w_6006));
  and_bi g1410(.a(n1408),.b(n1409),.q(n1410));
  bfr _b_6062(.a(_w_7487),.q(_w_7488));
  and_bi g577(.a(G177_27),.b(n576),.q(n577));
  and_bi g1402(.a(G141_5),.b(n1401),.q(n1402));
  spl3L G145_s_1(.a(G145_3),.q0(G145_4),.q1(G145_5),.q2(G145_6));
  bfr _b_2761(.a(_w_4186),.q(_w_4187));
  spl4L g588_s_0(.a(n588),.q0(n588_0),.q1(n588_1),.q2(n588_2),.q3(n588_3));
  and_bi g1401(.a(n1399),.b(n1400),.q(n1401));
  bfr _b_3428(.a(_w_4853),.q(n1441));
  bfr _b_2292(.a(_w_3717),.q(G167_0));
  bfr _b_7145(.a(_w_8570),.q(_w_8571));
  spl2 g1027_s_1(.a(G5293_3),.q0(G5293_4),.q1(G5293_5));
  and_bi g1330(.a(G157_3),.b(n1329),.q(n1330));
  bfr _b_3414(.a(_w_4839),.q(_w_4840));
  or_bb g1397(.a(n1386_1),.b(n1395_1),.q(n1397));
  or_bb g1393(.a(n1391),.b(n1392),.q(n1393));
  bfr _b_2439(.a(_w_3864),.q(_w_3865));
  bfr _b_2780(.a(_w_4205),.q(n415_1));
  spl2 g1297_s_0(.a(n1297),.q0(n1297_0),.q1(n1297_1));
  bfr _b_7232(.a(_w_8657),.q(_w_8658));
  and_bi g1388(.a(G105_11),.b(G101_16),.q(n1388));
  or_bb g1386(.a(n1381),.b(n1385),.q(n1386));
  spl2 g485_s_0(.a(n485),.q0(n485_0),.q1(n485_1));
  bfr _b_4985(.a(_w_6410),.q(_w_6409));
  spl2 g503_s_0(.a(n503),.q0(n503_0),.q1(n503_1));
  bfr _b_7410(.a(_w_8835),.q(_w_8836));
  bfr _b_3948(.a(_w_5373),.q(_w_5374));
  and_bi g1383(.a(G98_15),.b(G107_13),.q(n1383));
  bfr _b_2305(.a(_w_3730),.q(_w_3731));
  and_bb g187(.a(G163_0),.b(_w_7455),.q(_w_6227));
  bfr _b_4136(.a(_w_5561),.q(_w_5562));
  and_bi g1380(.a(n1378),.b(n1379),.q(n1380));
  bfr _b_7021(.a(_w_8446),.q(_w_8447));
  or_bb g1378(.a(G100_9),.b(G107_10),.q(n1378));
  or_bb g1377(.a(n1375),.b(n1376),.q(_w_4290));
  spl2 g737_s_0(.a(n737),.q0(n737_0),.q1(n737_1));
  bfr _b_2526(.a(_w_3951),.q(n399_2));
  spl4L g625_s_0(.a(G5255_0),.q0(_w_3682),.q1(G5255_1),.q2(G5255_2),.q3(G5255_3));
  and_bi g1376(.a(n1362_1),.b(n1374_1),.q(n1376));
  bfr _b_2312(.a(_w_3737),.q(_w_3738));
  bfr _b_5793(.a(_w_7218),.q(_w_7219));
  bfr _b_3475(.a(_w_4900),.q(_w_4901));
  spl2 g763_s_0(.a(n763),.q0(n763_0),.q1(n763_1));
  bfr _b_6728(.a(_w_8153),.q(_w_8154));
  and_bi g1374(.a(n1373),.b(n1372),.q(n1374));
  or_bb g1373(.a(n1371_1),.b(n346_3),.q(n1373));
  bfr _b_2206(.a(_w_3631),.q(_w_3632));
  and_bi g1370(.a(n1369),.b(G140_6),.q(n1370));
  bfr _b_3894(.a(_w_5319),.q(_w_5320));
  bfr _b_6935(.a(_w_8360),.q(_w_8361));
  bfr _b_5046(.a(_w_6471),.q(_w_6472));
  bfr _b_2102(.a(_w_3527),.q(_w_3528));
  bfr _b_1958(.a(_w_3383),.q(G176_41));
  bfr _b_3254(.a(_w_4679),.q(_w_4680));
  bfr _b_3399(.a(_w_4824),.q(_w_4825));
  bfr _b_6046(.a(_w_7471),.q(_w_7472));
  or_bb g1369(.a(n1367),.b(n1368),.q(n1369));
  and_bi g353(.a(G166_13),.b(G103_6),.q(n353));
  and_bi g1368(.a(G98_14),.b(G94_13),.q(n1368));
  bfr _b_2202(.a(_w_3627),.q(_w_3628));
  bfr _b_3464(.a(_w_4889),.q(_w_4890));
  bfr _b_7496(.a(_w_8921),.q(_w_8922));
  spl2 g698_s_0(.a(n698),.q0(n698_0),.q1(n698_1));
  bfr _b_4626(.a(_w_6051),.q(G5308));
  and_bb g1367(.a(G102_13),.b(G94_12),.q(n1367));
  bfr _b_2458(.a(_w_3883),.q(_w_3884));
  bfr _b_3618(.a(_w_5043),.q(_w_5044));
  spl4L g406_s_0(.a(n406),.q0(n406_0),.q1(n406_1),.q2(n406_2),.q3(n406_3));
  inv inv_G1(.a(G1_1),.q(i_G1));
  bfr _b_6382(.a(_w_7807),.q(_w_7808));
  bfr _b_4010(.a(_w_5435),.q(G176_51));
  spl2 g574_s_0(.a(n574),.q0(n574_0),.q1(n574_1));
  or_bb g1362(.a(n1360),.b(n1361),.q(n1362));
  bfr _b_5538(.a(_w_6963),.q(_w_6964));
  bfr _b_2171(.a(_w_3596),.q(_w_3597));
  spl2 g482_s_0(.a(G5239_0),.q0(G5239),.q1(G5240));
  bfr _b_6198(.a(_w_7623),.q(_w_7624));
  and_bb g347(.a(n337_0),.b(n346_0),.q(_w_4889));
  bfr _b_7179(.a(_w_8604),.q(_w_8605));
  bfr _b_6969(.a(_w_8394),.q(_w_8395));
  or_bb g1043(.a(n1039),.b(n1042),.q(_w_6100));
  bfr _b_3303(.a(_w_4728),.q(_w_4729));
  bfr _b_3434(.a(_w_4859),.q(G145_3));
  or_bb g1359(.a(n1354),.b(n1358),.q(n1359));
  and_bi g1358(.a(n1357),.b(G144_6),.q(n1358));
  bfr _b_4008(.a(_w_5433),.q(_w_5434));
  bfr _b_6657(.a(_w_8082),.q(_w_8083));
  bfr _b_5814(.a(_w_7239),.q(_w_7240));
  or_bb g1357(.a(n1355),.b(n1356),.q(n1357));
  bfr _b_2574(.a(_w_3999),.q(_w_4000));
  bfr _b_6149(.a(_w_7574),.q(_w_7575));
  spl2 G177_s_5(.a(G177_17),.q0(G177_20),.q1(G177_21));
  and_bi g1354(.a(G144_5),.b(n1353),.q(n1354));
  and_bi g1353(.a(n1351),.b(n1352),.q(n1353));
  bfr _b_3999(.a(_w_5424),.q(_w_5425));
  and_bi g1352(.a(G92_11),.b(G101_13),.q(n1352));
  or_bb g1351(.a(G100_11),.b(G92_10),.q(n1351));
  and_ii g984(.a(n979),.b(n983),.q(_w_6069));
  bfr _b_2023(.a(_w_3448),.q(_w_3449));
  or_bb g1348(.a(n1346),.b(n1347),.q(n1348));
  bfr _b_2090(.a(_w_3515),.q(n393_1));
  bfr _b_3862(.a(_w_5287),.q(_w_5288));
  and_bi g1347(.a(G98_12),.b(G90_13),.q(n1347));
  or_bb g802(.a(G158_26),.b(G159_4),.q(n802));
  bfr _b_5655(.a(_w_7080),.q(_w_7081));
  spl2 g620_s_0(.a(n620),.q0(n620_0),.q1(n620_1));
  and_bb g1346(.a(G102_11),.b(G90_12),.q(n1346));
  and_bi g1345(.a(G143_5),.b(n1344),.q(n1345));
  spl4L G102_s_0(.a(_w_6395),.q0(G102_0),.q1(G102_1),.q2(G102_2),.q3(G102_3));
  bfr _b_5525(.a(_w_6950),.q(_w_6951));
  bfr _b_2182(.a(_w_3607),.q(_w_3608));
  spl4L G64_s_2(.a(G64_1),.q0(G64_8),.q1(G64_9),.q2(G64_10),.q3(G64_11));
  or_bb g1074(.a(n1072),.b(n1073),.q(n1074));
  or_bb g1342(.a(G100_12),.b(G90_10),.q(n1342));
  or_bb g1341(.a(n1338),.b(n1340),.q(n1341));
  and_bb g1295(.a(G157_1),.b(n1294),.q(n1295));
  and_bi g1339(.a(n1297_1),.b(n1337_1),.q(n1339));
  bfr _b_6375(.a(_w_7800),.q(_w_7801));
  spl4L g394_s_0(.a(n394),.q0(n394_0),.q1(_w_4295),.q2(_w_4297),.q3(n394_3));
  bfr _b_7488(.a(_w_8913),.q(_w_8914));
  bfr _b_6921(.a(_w_8346),.q(_w_8347));
  spl4L G103_s_2(.a(G103_2),.q0(G103_6),.q1(G103_7),.q2(G103_8),.q3(G103_9));
  bfr _b_4066(.a(_w_5491),.q(_w_5492));
  and_bi g1335(.a(n1332_0),.b(n1334_0),.q(n1335));
  bfr _b_3605(.a(_w_5030),.q(_w_5031));
  bfr _b_5368(.a(_w_6793),.q(_w_6794));
  bfr _b_3291(.a(_w_4716),.q(G5253));
  bfr _b_4214(.a(_w_5639),.q(_w_5640));
  and_bi g1329(.a(n1324_1),.b(n403_3),.q(n1329));
  or_bb g1325(.a(G157_2),.b(n1324_0),.q(n1325));
  bfr _b_7138(.a(_w_8563),.q(_w_8564));
  and_bi g717(.a(n384_2),.b(n378_2),.q(n717));
  bfr _b_2002(.a(_w_3427),.q(_w_3428));
  or_bb g1323(.a(n1322),.b(n542_4),.q(n1323));
  or_bb g1321(.a(n1314_0),.b(n1320_0),.q(_w_4310));
  or_bb g731(.a(n729),.b(n730),.q(_w_5296));
  or_bb g1320(.a(n1318),.b(n1319),.q(n1320));
  bfr _b_7065(.a(_w_8490),.q(_w_8491));
  bfr _b_2438(.a(_w_3863),.q(_w_3864));
  spl2 g1015_s_1(.a(G5291_3),.q0(G5291_4),.q1(G5291_5));
  or_bb g305(.a(n303),.b(n304),.q(n305));
  or_bb g1340(.a(G176_32),.b(n1339),.q(n1340));
  bfr _b_2554(.a(_w_3979),.q(_w_3980));
  and_bi g1319(.a(n1317_1),.b(n1303_3),.q(n1319));
  bfr _b_4072(.a(_w_5497),.q(_w_5498));
  bfr _b_3857(.a(_w_5282),.q(_w_5283));
  bfr _b_4907(.a(_w_6332),.q(_w_6333));
  bfr _b_5332(.a(G158),.q(_w_6758));
  and_bi g1315(.a(n426_2),.b(n415_4),.q(n1315));
  bfr _b_5743(.a(_w_7168),.q(_w_7169));
  and_bi g1314(.a(n1313),.b(n546_1),.q(_w_4311));
  or_bb g1423(.a(n1421),.b(n1422),.q(n1423));
  and_bi g554(.a(n442_1),.b(G21_0),.q(n554));
  bfr _b_7537(.a(_w_8962),.q(_w_8963));
  and_bi g1311(.a(n1310),.b(n1309),.q(n1311));
  bfr _b_2110(.a(_w_3535),.q(_w_3536));
  bfr _b_3603(.a(_w_5028),.q(_w_5029));
  bfr _b_7207(.a(_w_8632),.q(_w_8633));
  spl3L G161_s_1(.a(G161_1),.q0(G161_4),.q1(G161_5),.q2(_w_4288));
  spl2 G77_s_0(.a(_w_8569),.q0(G77_0),.q1(G77_1));
  and_bi g417(.a(_w_8948),.b(G124_9),.q(n417));
  bfr _b_7356(.a(_w_8781),.q(_w_8782));
  bfr _b_6071(.a(_w_7496),.q(_w_7497));
  bfr _b_3552(.a(_w_4977),.q(G98_4));
  and_bb g1306(.a(n1303_0),.b(n1305_0),.q(n1306));
  and_bi g1422(.a(G98_19),.b(G103_13),.q(n1422));
  spl2 g600_s_0(.a(n600),.q0(n600_0),.q1(n600_1));
  or_bb g1135(.a(n1131),.b(n1134),.q(n1135));
  and_bi g1457(.a(G175_14),.b(n1456),.q(_w_4319));
  and_bi g1296(.a(n1295),.b(n1293),.q(n1296));
  spl4L g472_s_0(.a(n472),.q0(n472_0),.q1(n472_1),.q2(_w_4321),.q3(n472_3));
  bfr _b_6125(.a(_w_7550),.q(_w_7551));
  spl3L G1_s_0(.a(_w_6354),.q0(_w_4322),.q1(G1_0),.q2(G1_1));
  or_bb g1292(.a(n1290),.b(n1291),.q(n1292));
  spl2 g337_s_0(.a(n337),.q0(n337_0),.q1(_w_4324));
  bfr _b_7380(.a(_w_8805),.q(_w_8806));
  and_bi g1291(.a(n1289_1),.b(n1288_1),.q(n1291));
  bfr _b_4238(.a(_w_5663),.q(_w_5664));
  and_bi g1290(.a(n1288_0),.b(n1289_0),.q(n1290));
  or_bb g618(.a(n451_1),.b(n617_0),.q(n618));
  bfr _b_4478(.a(_w_5903),.q(_w_5904));
  bfr _b_7294(.a(_w_8719),.q(_w_8720));
  and_bb g714(.a(n391_2),.b(n397_2),.q(n714));
  and_bb g572(.a(G2_0),.b(n381_1),.q(n572));
  bfr _b_6416(.a(_w_7841),.q(_w_7821));
  bfr _b_3391(.a(_w_4816),.q(_w_4817));
  and_bi g705(.a(n704_0),.b(n442_5),.q(n705));
  bfr _b_3032(.a(_w_4457),.q(n426_1));
  bfr _b_4347(.a(_w_5772),.q(_w_5773));
  bfr _b_4204(.a(_w_5629),.q(_w_5630));
  or_bb g695(.a(n693),.b(n694),.q(_w_4340));
  and_bi g994(.a(G177_13),.b(n993),.q(_w_4898));
  bfr _b_4148(.a(_w_5573),.q(_w_5574));
  or_bb g1205(.a(n1184_0),.b(n1204_0),.q(_w_4344));
  spl2 g1289_s_0(.a(n1289),.q0(n1289_0),.q1(n1289_1));
  spl4L g469_s_0(.a(n469),.q0(n469_0),.q1(n469_1),.q2(n469_2),.q3(n469_3));
  and_bi g297(.a(n296),.b(G143_1),.q(n297));
  bfr _b_4603(.a(_w_6028),.q(_w_6029));
  and_bi g681(.a(G177_20),.b(n680),.q(n681));
  bfr _b_3486(.a(_w_4911),.q(_w_4912));
  spl4L g978_s_0(.a(G5285_0),.q0(_w_4345),.q1(G5285_1),.q2(G5285_2),.q3(G5285_3));
  and_bi g690(.a(n689_0),.b(n686_0),.q(n690));
  bfr _b_5293(.a(_w_6718),.q(_w_6719));
  bfr _b_2817(.a(_w_4242),.q(_w_4243));
  bfr _b_5317(.a(_w_6742),.q(_w_6743));
  bfr _b_3929(.a(_w_5354),.q(_w_5355));
  or_bb g1425(.a(n1420),.b(n1424),.q(n1425));
  bfr _b_7218(.a(_w_8643),.q(_w_8644));
  bfr _b_7044(.a(_w_8469),.q(_w_8470));
  and_bb g925(.a(G86_1),.b(n815_1),.q(n925));
  and_bi g888(.a(G76_0),.b(n802_1),.q(n888));
  and_bi g238(.a(G150_0),.b(n237),.q(n238));
  bfr _b_4260(.a(_w_5685),.q(_w_5686));
  bfr _b_5750(.a(G2),.q(_w_7176));
  bfr _b_2303(.a(_w_3728),.q(G173_5));
  bfr _b_4860(.a(_w_6285),.q(n220));
  bfr _b_4939(.a(_w_6364),.q(_w_6365));
  bfr _b_7292(.a(_w_8717),.q(_w_8718));
  bfr _b_2031(.a(_w_3456),.q(_w_3457));
  bfr _b_5092(.a(_w_6517),.q(_w_6518));
  and_bb g863(.a(n860),.b(n862),.q(_w_4353));
  spl4L g456_s_0(.a(n456),.q0(n456_0),.q1(_w_3936),.q2(_w_3937),.q3(n456_3));
  and_ii g683(.a(n676),.b(n682),.q(_w_4355));
  spl2 G86_s_0(.a(_w_8875),.q0(G86_0),.q1(G86_1));
  or_bb g1075(.a(n1071),.b(n1074),.q(_w_4364));
  bfr _b_5760(.a(_w_7185),.q(_w_7186));
  or_bb g767(.a(n421_1),.b(n766_0),.q(n767));
  bfr _b_5324(.a(_w_6749),.q(_w_6750));
  and_bi g1166(.a(G145_6),.b(n464_2),.q(_w_4367));
  bfr _b_2712(.a(_w_4137),.q(_w_4138));
  or_bb g773(.a(n477_1),.b(n772),.q(n773));
  and_bb g672(.a(G176_52),.b(n365_1),.q(n672));
  or_bb g222(.a(n220),.b(n221),.q(_w_4368));
  and_bb g873(.a(G26_1),.b(n630_5),.q(n873));
  bfr _b_2187(.a(_w_3612),.q(_w_3613));
  bfr _b_3926(.a(_w_5351),.q(_w_5352));
  or_bb g1091(.a(n1087),.b(n1090),.q(_w_6280));
  or_bb g893(.a(G158_22),.b(G5260_4),.q(n893));
  bfr _b_5280(.a(_w_6705),.q(_w_6706));
  bfr _b_2308(.a(_w_3733),.q(_w_3734));
  bfr _b_2613(.a(_w_4038),.q(_w_4039));
  bfr _b_7513(.a(_w_8938),.q(_w_8939));
  bfr _b_3390(.a(_w_4815),.q(_w_4816));
  or_bb g667(.a(n386_2),.b(n666_0),.q(n667));
  and_bi g1138(.a(G160_11),.b(G5287_5),.q(n1138));
  and_ii g663(.a(n651),.b(n662),.q(_w_4374));
  bfr _b_2115(.a(_w_3540),.q(_w_3541));
  bfr _b_4817(.a(_w_6242),.q(_w_6243));
  and_bb g684(.a(n456_2),.b(n469_5),.q(n684));
  bfr _b_2812(.a(_w_4237),.q(_w_4238));
  bfr _b_2965(.a(_w_4390),.q(_w_4391));
  or_bb g448(.a(n446),.b(n447),.q(_w_4382));
  and_bb g693(.a(G123_6),.b(G132_2),.q(n693));
  and_bb g647(.a(G176_48),.b(n327_1),.q(n647));
  bfr _b_5971(.a(_w_7396),.q(_w_7397));
  and_bi g1212(.a(n1211_0),.b(n253_2),.q(n1212));
  bfr _b_3111(.a(_w_4536),.q(_w_4537));
  spl2 G92_s_1(.a(G92_1),.q0(G92_4),.q1(G92_5));
  or_bb g643(.a(n641),.b(n642),.q(n643));
  bfr _b_3596(.a(_w_5021),.q(_w_5022));
  and_bi g1222(.a(n1221),.b(G147_6),.q(n1222));
  bfr _b_2175(.a(_w_3600),.q(_w_3601));
  and_bb g449(.a(G149_2),.b(n448_0),.q(n449));
  bfr _b_2760(.a(_w_4185),.q(n387_1));
  and_bb g637(.a(G2_2),.b(n403_1),.q(n637));
  bfr _b_3455(.a(_w_4880),.q(n249));
  and_bb g952(.a(G69_1),.b(n815_6),.q(n952));
  bfr _b_6489(.a(_w_7914),.q(_w_7915));
  bfr _b_4046(.a(_w_5471),.q(_w_5472));
  or_bb g1447(.a(n1263_1),.b(n1446),.q(n1447));
  bfr _b_6564(.a(_w_7989),.q(_w_7990));
  spl4L G170_s_0(.a(_w_6949),.q0(_w_4544),.q1(_w_4548),.q2(G170_2),.q3(G170_3));
  and_bi g633(.a(G22_1),.b(n632_0),.q(n633));
  spl2 g243_s_0(.a(n243),.q0(n243_0),.q1(_w_6233));
  bfr _b_6438(.a(_w_7863),.q(_w_7864));
  and_bb g1148(.a(G161_12),.b(n1147),.q(n1148));
  bfr _b_3756(.a(_w_5181),.q(_w_5182));
  and_bb g631(.a(G3_1),.b(n630_0),.q(n631));
  or_bb g696(.a(n438_2),.b(n448_2),.q(n696));
  or_bb g1269(.a(n379_3),.b(n386_5),.q(n1269));
  bfr _b_5932(.a(_w_7357),.q(_w_7358));
  spl3L g581_s_1(.a(G5251_3),.q0(G5251_4),.q1(G5251_5),.q2(G5251_6));
  spl2 g407_s_0(.a(n407),.q0(n407_0),.q1(_w_4118));
  and_bb g1312(.a(n1311_0),.b(n542_2),.q(n1312));
  and_bb g629(.a(n626),.b(n628),.q(_w_4399));
  bfr _b_3694(.a(_w_5119),.q(_w_5120));
  bfr _b_7058(.a(_w_8483),.q(_w_8484));
  bfr _b_6497(.a(_w_7922),.q(_w_7923));
  and_bi g957(.a(n469_7),.b(G61_0),.q(n957));
  bfr _b_4106(.a(_w_5531),.q(_w_5532));
  bfr _b_6966(.a(_w_8391),.q(_w_8392));
  and_bi g628(.a(G175_0),.b(n627),.q(n628));
  bfr _b_6259(.a(_w_7684),.q(_w_7685));
  bfr _b_3435(.a(_w_4860),.q(_w_4861));
  bfr _b_4720(.a(_w_6145),.q(_w_6146));
  spl4L G168_s_2(.a(G168_2),.q0(G168_6),.q1(G168_7),.q2(G168_8),.q3(G168_9));
  and_bi g627(.a(G174_27),.b(G5248_2),.q(n627));
  bfr _b_5389(.a(_w_6814),.q(_w_6815));
  bfr _b_2512(.a(_w_3937),.q(n456_2));
  bfr _b_2935(.a(_w_4360),.q(_w_4361));
  bfr _b_6567(.a(_w_7992),.q(_w_7993));
  bfr _b_4479(.a(_w_5904),.q(G173_0));
  bfr _b_5951(.a(G27),.q(_w_7377));
  and_bb g723(.a(n412_2),.b(n418_2),.q(n723));
  bfr _b_6860(.a(_w_8285),.q(_w_8286));
  spl2 g398_s_0(.a(n398),.q0(n398_0),.q1(_w_4400));
  and_bi g829(.a(G173_21),.b(G5254_1),.q(n829));
  bfr _b_4703(.a(_w_6128),.q(n968));
  or_bb g658(.a(n656),.b(n657),.q(n658));
  bfr _b_4672(.a(_w_6097),.q(_w_6098));
  bfr _b_6507(.a(_w_7932),.q(_w_7933));
  and_bi g620(.a(n618),.b(n619),.q(_w_4408));
  bfr _b_7451(.a(_w_8876),.q(_w_8877));
  bfr _b_1990(.a(_w_3415),.q(_w_3416));
  bfr _b_2551(.a(_w_3976),.q(_w_3977));
  spl2 g1350_s_0(.a(n1350),.q0(n1350_0),.q1(n1350_1));
  bfr _b_3884(.a(_w_5309),.q(_w_5310));
  or_bb g746(.a(n547_1),.b(n745),.q(n746));
  and_ii g615(.a(n606),.b(n614),.q(_w_4410));
  spl3L g428_s_0(.a(n428),.q0(n428_0),.q1(_w_4417),.q2(n428_2));
  bfr _b_3348(.a(_w_4773),.q(_w_4774));
  bfr _b_2615(.a(_w_4040),.q(_w_4041));
  and_bi g1085(.a(G174_7),.b(G5288_2),.q(n1085));
  bfr _b_6347(.a(_w_7772),.q(_w_7773));
  bfr _b_3188(.a(_w_4613),.q(G158_6));
  bfr _b_6824(.a(_w_8249),.q(_w_8250));
  spl2 G36_s_0(.a(_w_7458),.q0(G36_0),.q1(G36_1));
  bfr _b_6587(.a(_w_8012),.q(_w_8013));
  bfr _b_2209(.a(_w_3634),.q(_w_3635));
  and_bi g589(.a(G22_0),.b(n588_0),.q(n589));
  or_bb g426(.a(G140_4),.b(n424_1),.q(n426));
  bfr _b_6898(.a(_w_8323),.q(_w_8324));
  or_bb g588(.a(G172_5),.b(G173_25),.q(n588));
  and_bi g421(.a(n420_0),.b(n419_0),.q(n421));
  and_bi g1303(.a(n1301),.b(n1302),.q(n1303));
  bfr _b_5972(.a(_w_7397),.q(_w_7398));
  and_bb g823(.a(n820),.b(n822),.q(n823));
  bfr _b_3490(.a(_w_4915),.q(_w_4916));
  and_bi g586(.a(G173_26),.b(G172_4),.q(n586));
  and_bi g1394(.a(n1393),.b(G138_6),.q(n1394));
  and_bb g382(.a(G107_7),.b(G124_22),.q(n382));
  bfr _b_4513(.a(_w_5938),.q(_w_5939));
  bfr _b_7181(.a(_w_8606),.q(_w_8607));
  bfr _b_4578(.a(_w_6003),.q(_w_6004));
  bfr _b_4624(.a(_w_6049),.q(n909));
  bfr _b_6995(.a(_w_8420),.q(_w_8421));
  or_bb g385(.a(G139_2),.b(n384_0),.q(n385));
  and_bb g571(.a(_w_7799),.b(n552_24),.q(n571));
  and_bb g592(.a(_w_7153),.b(n552_23),.q(n592));
  and_bi g894(.a(G158_21),.b(G5249_4),.q(n894));
  bfr _b_2361(.a(_w_3786),.q(_w_3787));
  bfr _b_3707(.a(_w_5132),.q(_w_5133));
  spl2 g1308_s_0(.a(n1308),.q0(n1308_0),.q1(n1308_1));
  and_ii g570(.a(n562),.b(n569),.q(_w_4429));
  bfr _b_2088(.a(_w_3513),.q(_w_3514));
  bfr _b_5022(.a(_w_6447),.q(_w_6448));
  bfr _b_5233(.a(_w_6658),.q(_w_6659));
  bfr _b_2350(.a(_w_3775),.q(_w_3776));
  bfr _b_7115(.a(_w_8540),.q(_w_8541));
  and_bi g1086(.a(G175_13),.b(n1085),.q(n1086));
  and_bb g871(.a(n868),.b(n870),.q(_w_6031));
  spl2 g1320_s_0(.a(n1320),.q0(n1320_0),.q1(n1320_1));
  bfr _b_5015(.a(G132),.q(_w_6440));
  and_bb g569(.a(n566),.b(n568),.q(_w_4436));
  and_bi g501(.a(n497_0),.b(n500_0),.q(n501));
  or_bb g909(.a(n905),.b(n908),.q(_w_6049));
  spl4L g426_s_0(.a(n426),.q0(n426_0),.q1(_w_4444),.q2(_w_4458),.q3(_w_4462));
  and_bi g492(.a(G130_4),.b(G132_0),.q(n492));
  and_bi g560(.a(n559),.b(n557),.q(_w_4466));
  or_bb g365(.a(n360),.b(n364),.q(_w_4467));
  bfr _b_6739(.a(_w_8164),.q(_w_8165));
  bfr _b_3635(.a(_w_5060),.q(_w_5061));
  and_bi g645(.a(n644),.b(n637_0),.q(n645));
  and_bi g559(.a(G177_29),.b(n558),.q(n559));
  bfr _b_6051(.a(_w_7476),.q(_w_7477));
  or_bb g876(.a(G174_16),.b(G5260_2),.q(n876));
  and_bi g903(.a(G158_17),.b(G5255_4),.q(n903));
  spl2 g1226_s_0(.a(n1226),.q0(n1226_0),.q1(n1226_1));
  bfr _b_4951(.a(_w_6376),.q(_w_6377));
  and_bb g553(.a(_w_8113),.b(n552_14),.q(n553));
  bfr _b_4697(.a(_w_6122),.q(_w_6123));
  bfr _b_2654(.a(_w_4079),.q(_w_4080));
  and_bi g341(.a(G142_0),.b(n340),.q(n341));
  spl4L G176_s_6(.a(G176_12),.q0(_w_4515),.q1(G176_23),.q2(G176_24),.q3(G176_25));
  bfr _b_2656(.a(_w_4081),.q(_w_4082));
  bfr _b_6435(.a(_w_7860),.q(_w_7861));
  or_bb g550(.a(n543),.b(n549),.q(_w_4523));
  or_bb g549(.a(n407_1),.b(n548),.q(_w_4543));
  bfr _b_3657(.a(_w_5082),.q(_w_5083));
  and_bi g630(.a(G174_26),.b(G175_4),.q(n630));
  bfr _b_7405(.a(_w_8830),.q(_w_8831));
  and_bi g1008(.a(n1007),.b(n1005),.q(n1008));
  bfr _b_5567(.a(_w_6992),.q(_w_6993));
  spl2 g473_s_0(.a(n473),.q0(n473_0),.q1(n473_1));
  bfr _b_7106(.a(_w_8531),.q(_w_8532));
  bfr _b_6308(.a(_w_7733),.q(_w_7734));
  bfr _b_2673(.a(_w_4098),.q(_w_4099));
  or_bb g595(.a(n433_1),.b(n594_0),.q(n595));
  and_bb g537(.a(n393_1),.b(n536),.q(n537));
  and_bi g1273(.a(n537_5),.b(n1272_0),.q(n1273));
  spl4L G174_s_0(.a(_w_7032),.q0(_w_4552),.q1(_w_4554),.q2(_w_4556),.q3(G174_3));
  or_bb g536(.a(n534_0),.b(n535),.q(n536));
  and_bi g284(.a(G140_0),.b(n283),.q(n284));
  spl2 g430_s_0(.a(n430),.q0(n430_0),.q1(n430_1));
  or_bb g535(.a(n386_1),.b(n392_1),.q(_w_4558));
  bfr _b_3197(.a(_w_4622),.q(_w_4623));
  spl2 g1198_s_0(.a(n1198),.q0(n1198_0),.q1(n1198_1));
  bfr _b_4927(.a(_w_6352),.q(n689));
  bfr _b_5774(.a(_w_7199),.q(_w_7200));
  bfr _b_5034(.a(_w_6459),.q(_w_6460));
  and_bb g1460(.a(G4_1),.b(n630_11),.q(n1460));
  bfr _b_5777(.a(_w_7202),.q(_w_7203));
  and_bb g596(.a(n434_1),.b(n595),.q(_w_4559));
  bfr _b_4453(.a(_w_5878),.q(n463_3));
  bfr _b_4518(.a(_w_5943),.q(_w_5944));
  or_bi g533(.a(n531),.b(n532),.q(_w_4562));
  bfr _b_3312(.a(_w_4737),.q(n1282));
  bfr _b_4207(.a(_w_5632),.q(_w_5633));
  bfr _b_5887(.a(_w_7312),.q(_w_7313));
  or_bb g724(.a(n412_3),.b(n418_3),.q(n724));
  and_ii g713(.a(n711),.b(n712),.q(_w_4585));
  bfr _b_6426(.a(_w_7851),.q(_w_7852));
  bfr _b_5930(.a(_w_7355),.q(_w_7356));
  bfr _b_4663(.a(_w_6088),.q(_w_6089));
  or_bb g532(.a(n515_1),.b(n530_1),.q(n532));
  and_bb g531(.a(n515_0),.b(n530_0),.q(n531));
  bfr _b_7445(.a(_w_8870),.q(_w_8871));
  bfr _b_4711(.a(_w_6136),.q(_w_6137));
  and_bb g429(.a(n415_0),.b(n428_0),.q(_w_4606));
  and_bi g528(.a(n524_0),.b(n527_0),.q(n528));
  bfr _b_6313(.a(_w_7738),.q(_w_7739));
  bfr _b_4803(.a(_w_6228),.q(n1063));
  bfr _b_6844(.a(_w_8269),.q(_w_8270));
  bfr _b_5322(.a(_w_6747),.q(_w_6748));
  bfr _b_4839(.a(_w_6264),.q(_w_6265));
  and_bi g942(.a(G70_1),.b(n813_5),.q(n942));
  bfr _b_7455(.a(_w_8880),.q(_w_8881));
  and_bb g664(.a(_w_7994),.b(n552_16),.q(_w_5751));
  bfr _b_4566(.a(_w_5991),.q(_w_5992));
  spl2 g298_s_0(.a(n298),.q0(n298_0),.q1(n298_1));
  and_bi g526(.a(G107_9),.b(G105_9),.q(n526));
  and_bb g523(.a(n518_1),.b(n521_1),.q(n523));
  bfr _b_2604(.a(_w_4029),.q(_w_4030));
  or_bb g522(.a(n518_0),.b(n521_0),.q(n522));
  bfr _b_4488(.a(_w_5913),.q(_w_5914));
  bfr _b_3147(.a(_w_4572),.q(_w_4573));
  or_bb g668(.a(n394_2),.b(n667_0),.q(n668));
  or_bb g634(.a(n631),.b(n633),.q(n634));
  or_ii g185(.a(G11_1),.b(_w_6424),.q(G5221_0));
  and_bb g768(.a(n421_2),.b(n766_1),.q(n768));
  bfr _b_2603(.a(_w_4028),.q(_w_4029));
  bfr _b_2594(.a(_w_4019),.q(_w_4020));
  bfr _b_6408(.a(_w_7833),.q(_w_7834));
  bfr _b_4546(.a(_w_5971),.q(_w_5972));
  bfr _b_6512(.a(_w_7937),.q(_w_7938));
  bfr _b_3653(.a(_w_5078),.q(_w_5079));
  bfr _b_7117(.a(_w_8542),.q(_w_8543));
  and_bi g736(.a(n731_1),.b(n734_1),.q(n736));
  bfr _b_3449(.a(_w_4874),.q(n1122));
  bfr _b_4025(.a(_w_5450),.q(G5259_0));
  bfr _b_4296(.a(_w_5721),.q(_w_5722));
  bfr _b_2215(.a(_w_3640),.q(_w_3641));
  or_bb g515(.a(n513),.b(n514),.q(_w_4608));
  bfr _b_2263(.a(_w_3688),.q(_w_3689));
  bfr _b_3660(.a(_w_5085),.q(_w_5086));
  bfr _b_2013(.a(_w_3438),.q(G176_7));
  bfr _b_6155(.a(_w_7580),.q(_w_7581));
  bfr _b_4747(.a(_w_6172),.q(G150_4));
  and_bi g510(.a(G92_8),.b(G94_8),.q(n510));
  spl4L G158_s_1(.a(G158_0),.q0(G158_4),.q1(G158_5),.q2(_w_4611),.q3(G158_7));
  and_bi g509(.a(n507),.b(n508),.q(n509));
  spl3L g458_s_0(.a(n458),.q0(n458_0),.q1(n458_1),.q2(_w_4704));
  bfr _b_5029(.a(_w_6454),.q(_w_6455));
  and_bb g508(.a(G88_7),.b(G90_9),.q(n508));
  bfr _b_2731(.a(_w_4156),.q(_w_4157));
  bfr _b_7252(.a(_w_8677),.q(_w_8678));
  bfr _b_4620(.a(_w_6045),.q(_w_6046));
  bfr _b_5043(.a(_w_6468),.q(_w_6469));
  and_bi g1279(.a(n1276),.b(n1278),.q(n1279));
  bfr _b_5836(.a(_w_7261),.q(_w_7262));
  and_bb g702(.a(n432_2),.b(n476_2),.q(n702));
  bfr _b_7359(.a(_w_8784),.q(_w_8785));
  bfr _b_7101(.a(_w_8526),.q(_w_8527));
  bfr _b_6118(.a(_w_7543),.q(_w_7544));
  or_bb g626(.a(G174_15),.b(G5250_2),.q(n626));
  bfr _b_6181(.a(_w_7606),.q(_w_7607));
  or_bb g858(.a(n856),.b(n857),.q(n858));
  or_bb g760(.a(n545_1),.b(n759),.q(n760));
  or_bb g319(.a(G169_11),.b(G96_0),.q(n319));
  bfr _b_3448(.a(_w_4873),.q(n318));
  and_bb g928(.a(G64_19),.b(n927),.q(G5279));
  bfr _b_2300(.a(_w_3725),.q(_w_3726));
  or_bb g503(.a(n501),.b(n502),.q(n503));
  or_bb g813(.a(G160_26),.b(G161_4),.q(n813));
  and_bb g1054(.a(G172_12),.b(n1053),.q(n1054));
  bfr _b_2585(.a(_w_4010),.q(_w_4011));
  bfr _b_5098(.a(_w_6523),.q(_w_6524));
  spl2 g509_s_0(.a(n509),.q0(n509_0),.q1(n509_1));
  and_bi g1299(.a(n1298_0),.b(n413_2),.q(n1299));
  bfr _b_5846(.a(_w_7271),.q(_w_7272));
  bfr _b_5378(.a(_w_6803),.q(_w_6804));
  and_bi g1177(.a(n469_9),.b(n464_4),.q(n1177));
  bfr _b_2887(.a(_w_4312),.q(n1314));
  bfr _b_4609(.a(_w_6034),.q(_w_6035));
  bfr _b_4766(.a(_w_6191),.q(_w_6192));
  and_bi g495(.a(G121_8),.b(n494_0),.q(n495));
  bfr _b_6510(.a(_w_7935),.q(_w_7936));
  bfr _b_2807(.a(_w_4232),.q(_w_4233));
  spl4L G101_s_1(.a(G101_0),.q0(G101_4),.q1(G101_5),.q2(G101_6),.q3(G101_7));
  bfr _b_4229(.a(_w_5654),.q(_w_5655));
  spl4L G126_s_3(.a(G126_3),.q0(G126_10),.q1(G126_11),.q2(G126_12),.q3(G126_13));
  or_bb g378(.a(n376),.b(n377),.q(n378));
  bfr _b_3066(.a(_w_4491),.q(_w_4492));
  and_bb g481(.a(n466_0),.b(n480),.q(n481));
  bfr _b_4782(.a(_w_6207),.q(n1031));
  and_bi g493(.a(G132_1),.b(G130_5),.q(n493));
  bfr _b_5144(.a(_w_6569),.q(_w_6570));
  and_bi g480(.a(n479_0),.b(n473_0),.q(_w_4637));
  spl4L G124_s_4(.a(G124_3),.q0(G124_16),.q1(G124_17),.q2(G124_18),.q3(G124_19));
  bfr _b_4682(.a(_w_6107),.q(_w_6108));
  bfr _b_6914(.a(_w_8339),.q(_w_8340));
  and_bb g181(.a(G1_0),.b(_w_6443),.q(_w_4642));
  spl4L G137_s_0(.a(_w_6484),.q0(G137_0),.q1(G137_1),.q2(_w_4643),.q3(G137_3));
  bfr _b_3062(.a(_w_4487),.q(_w_4488));
  bfr _b_5914(.a(_w_7339),.q(_w_7340));
  bfr _b_5570(.a(_w_6995),.q(_w_6996));
  spl2 g776_s_0(.a(n776),.q0(n776_0),.q1(n776_1));
  and_bi g1198(.a(n1197),.b(n1196),.q(n1198));
  bfr _b_6944(.a(_w_8369),.q(_w_8370));
  bfr _b_2146(.a(_w_3571),.q(_w_3572));
  bfr _b_4286(.a(_w_5711),.q(_w_5712));
  spl2 g1263_s_0(.a(n1263),.q0(n1263_0),.q1(n1263_1));
  or_bb g474(.a(_w_6428),.b(G123_8),.q(n474));
  bfr _b_2349(.a(_w_3774),.q(_w_3775));
  bfr _b_3167(.a(_w_4592),.q(_w_4593));
  bfr _b_6029(.a(_w_7454),.q(_w_7453));
  bfr _b_2861(.a(_w_4286),.q(_w_4287));
  bfr _b_4646(.a(_w_6071),.q(_w_6072));
  bfr _b_5741(.a(_w_7166),.q(_w_7167));
  bfr _b_3219(.a(_w_4644),.q(G137_2));
  bfr _b_2210(.a(_w_3635),.q(_w_3636));
  bfr _b_4692(.a(_w_6117),.q(_w_6118));
  or_bb g472(.a(n470),.b(n471),.q(_w_4648));
  and_bi g409(.a(n408_0),.b(n407_0),.q(n409));
  and_bi g1120(.a(G158_7),.b(G5285_4),.q(n1120));
  bfr _b_2814(.a(_w_4239),.q(G5291));
  bfr _b_7245(.a(_w_8670),.q(_w_8637));
  bfr _b_2025(.a(_w_3450),.q(n469_9));
  and_bi g230(.a(G98_5),.b(G119_4),.q(n230));
  bfr _b_5284(.a(_w_6709),.q(_w_6710));
  and_bb g970(.a(G5251_4),.b(n959_1),.q(n970));
  bfr _b_4217(.a(_w_5642),.q(_w_5643));
  and_bb g467(.a(G113_2),.b(G123_12),.q(n467));
  spl2 G80_s_0(.a(_w_8673),.q0(G80_0),.q1(G80_1));
  bfr _b_2005(.a(_w_3430),.q(_w_3431));
  bfr _b_4007(.a(_w_5432),.q(G5245_0));
  bfr _b_2264(.a(_w_3689),.q(G5255));
  and_bi g1057(.a(G40_0),.b(n588_9),.q(n1057));
  bfr _b_7506(.a(_w_8931),.q(_w_8932));
  and_bb g771(.a(n758),.b(n770),.q(_w_6054));
  or_bb g926(.a(n924),.b(n925),.q(n926));
  bfr _b_3869(.a(_w_5294),.q(_w_5295));
  spl2 g689_s_0(.a(n689),.q0(n689_0),.q1(n689_1));
  spl3L G149_s_1(.a(G149_3),.q0(_w_6114),.q1(G149_5),.q2(G149_6));
  bfr _b_3805(.a(_w_5230),.q(_w_5231));
  or_bb g1143(.a(n1141),.b(n1142),.q(n1143));
  bfr _b_2575(.a(_w_4000),.q(_w_4001));
  bfr _b_5394(.a(_w_6819),.q(_w_6820));
  bfr _b_4098(.a(_w_5523),.q(_w_5524));
  bfr _b_5292(.a(_w_6717),.q(_w_6718));
  and_bi g245(.a(G113_1),.b(G102_6),.q(n245));
  bfr _b_3567(.a(_w_4992),.q(_w_4993));
  bfr _b_4216(.a(_w_5641),.q(_w_5642));
  spl4L G144_s_0(.a(_w_6538),.q0(G144_0),.q1(G144_1),.q2(_w_3916),.q3(G144_3));
  and_bb g463(.a(G146_2),.b(n462_0),.q(n463));
  and_bb g979(.a(_w_7918),.b(n552_13),.q(_w_4656));
  and_bi g708(.a(n701_0),.b(n707_0),.q(n708));
  bfr _b_3460(.a(_w_4885),.q(_w_4886));
  and_bi g1208(.a(n1205),.b(n1207),.q(n1208));
  bfr _b_7382(.a(G84),.q(_w_8808));
  bfr _b_2366(.a(_w_3791),.q(_w_3792));
  and_bi g465(.a(n464_0),.b(n463_0),.q(n465));
  bfr _b_4745(.a(_w_6170),.q(_w_6171));
  spl3L G135_s_1(.a(G135_3),.q0(_w_4667),.q1(G135_5),.q2(G135_6));
  and_bi g519(.a(G109_8),.b(G111_0),.q(n519));
  bfr _b_4509(.a(_w_5934),.q(_w_5935));
  and_bi g1156(.a(G160_7),.b(G5285_5),.q(n1156));
  bfr _b_3934(.a(_w_5359),.q(_w_5360));
  bfr _b_4402(.a(_w_5827),.q(G5313));
  and_bi g330(.a(G107_4),.b(G168_11),.q(n330));
  spl2 g277_s_0(.a(n277),.q0(n277_0),.q1(_w_4675));
  bfr _b_3485(.a(_w_4910),.q(_w_4911));
  bfr _b_6580(.a(_w_8005),.q(_w_8006));
  bfr _b_4418(.a(_w_5843),.q(_w_5844));
  bfr _b_7265(.a(_w_8690),.q(_w_8691));
  and_bb g824(.a(G16_0),.b(n586_1),.q(n824));
  bfr _b_4017(.a(_w_5442),.q(n905));
  bfr _b_2255(.a(_w_3680),.q(_w_3681));
  bfr _b_7246(.a(G8),.q(_w_8672));
  bfr _b_3269(.a(_w_4694),.q(_w_4695));
  bfr _b_2230(.a(_w_3655),.q(G159_6));
  bfr _b_6758(.a(_w_8183),.q(_w_8148));
  bfr _b_5556(.a(_w_6981),.q(_w_6982));
  spl2 g1371_s_0(.a(n1371),.q0(n1371_0),.q1(n1371_1));
  bfr _b_3006(.a(_w_4431),.q(_w_4432));
  bfr _b_3960(.a(_w_5385),.q(_w_5386));
  and_bb g180(.a(G66_0),.b(_w_8224),.q(_w_4678));
  or_bb g1134(.a(n1132),.b(n1133),.q(n1134));
  bfr _b_4073(.a(_w_5498),.q(_w_5499));
  and_bi g451(.a(n450_0),.b(n449_0),.q(_w_4679));
  bfr _b_3876(.a(_w_5301),.q(_w_5302));
  or_bb g450(.a(G149_4),.b(n448_1),.q(n450));
  bfr _b_7444(.a(_w_8869),.q(_w_8870));
  bfr _b_4181(.a(_w_5606),.q(_w_5607));
  bfr _b_4611(.a(_w_6036),.q(_w_6037));
  bfr _b_5749(.a(_w_7174),.q(_w_7153));
  spl2 G18_s_0(.a(_w_7120),.q0(G18_0),.q1(G18_1));
  and_bi g1324(.a(n1321),.b(n1323),.q(n1324));
  and_bi g853(.a(G174_23),.b(G5253_2),.q(n853));
  bfr _b_5885(.a(G25),.q(_w_7311));
  or_bb g444(.a(n442_0),.b(n443_0),.q(n444));
  bfr _b_2621(.a(_w_4046),.q(_w_4047));
  and_bi g300(.a(G92_4),.b(G168_8),.q(n300));
  bfr _b_4719(.a(_w_6144),.q(_w_6145));
  and_bi g240(.a(G166_0),.b(G128_6),.q(n240));
  spl4L G161_s_3(.a(G161_3),.q0(G161_11),.q1(G161_12),.q2(G161_13),.q3(G161_14));
  bfr _b_4006(.a(_w_5431),.q(_w_5432));
  bfr _b_3042(.a(_w_4467),.q(_w_4468));
  or_bb g971(.a(G5251_5),.b(n959_2),.q(n971));
  and_bi g321(.a(n319),.b(n320),.q(n321));
  bfr _b_6996(.a(_w_8421),.q(_w_8422));
  bfr _b_1999(.a(_w_3424),.q(_w_3425));
  bfr _b_6972(.a(_w_8397),.q(_w_8398));
  bfr _b_4328(.a(_w_5753),.q(_w_5754));
  bfr _b_4892(.a(_w_6317),.q(n1184));
  and_bi g762(.a(n415_2),.b(n760_1),.q(n762));
  and_bi g358(.a(G105_4),.b(G168_13),.q(n358));
  or_bb g438(.a(n436),.b(n437),.q(n438));
  and_bi g302(.a(G144_0),.b(n301),.q(n302));
  bfr _b_4628(.a(_w_6053),.q(n914));
  bfr _b_7536(.a(_w_8961),.q(_w_8962));
  and_bi g437(.a(G129_0),.b(G123_22),.q(n437));
  or_bb g1363(.a(G100_10),.b(G94_10),.q(n1363));
  and_bi g811(.a(G161_0),.b(n810),.q(n811));
  bfr _b_2212(.a(_w_3637),.q(n421_3));
  bfr _b_4009(.a(_w_5434),.q(_w_5435));
  bfr _b_4708(.a(_w_6133),.q(n991));
  and_bi g272(.a(G149_0),.b(n271),.q(n272));
  bfr _b_2668(.a(_w_4093),.q(_w_4094));
  bfr _b_2137(.a(_w_3562),.q(_w_3563));
  or_bb g1221(.a(n1219),.b(n1220),.q(n1221));
  bfr _b_6691(.a(_w_8116),.q(_w_8117));
  or_bb g296(.a(n294),.b(n295),.q(n296));
  spl4L g804_s_2(.a(n804_3),.q0(n804_8),.q1(n804_9),.q2(n804_10),.q3(n804_11));
  spl2 g1285_s_0(.a(n1285),.q0(n1285_0),.q1(n1285_1));
  bfr _b_2534(.a(_w_3959),.q(_w_3960));
  and_bi g1019(.a(G177_10),.b(n1018),.q(_w_5624));
  and_bb g808(.a(G64_25),.b(n807),.q(G5265));
  bfr _b_5870(.a(_w_7295),.q(_w_7296));
  or_bb g610(.a(n608),.b(n609),.q(n610));
  or_bb g241(.a(n239),.b(n240),.q(n241));
  bfr _b_5116(.a(G145),.q(_w_6542));
  bfr _b_3216(.a(_w_4641),.q(n480));
  bfr _b_3662(.a(_w_5087),.q(_w_5088));
  bfr _b_2186(.a(_w_3611),.q(_w_3612));
  spl4L G102_s_2(.a(G102_1),.q0(G102_7),.q1(G102_8),.q2(G102_9),.q3(G102_10));
  and_bb g1477(.a(G78_1),.b(n815_11),.q(n1477));
  spl2 g491_s_0(.a(n491),.q0(n491_0),.q1(n491_1));
  bfr _b_3321(.a(_w_4746),.q(_w_4747));
  or_bb g289(.a(n284),.b(n288),.q(_w_4682));
  and_bi g288(.a(n287),.b(G140_1),.q(n288));
  bfr _b_2317(.a(_w_3742),.q(_w_3743));
  bfr _b_2342(.a(_w_3767),.q(_w_3768));
  and_bi g206(.a(_w_8330),.b(G163_11),.q(_w_4699));
  bfr _b_6952(.a(_w_8377),.q(_w_8378));
  and_bi g761(.a(n760_0),.b(n415_1),.q(n761));
  bfr _b_3059(.a(_w_4484),.q(_w_4485));
  or_bb g1067(.a(n1063),.b(n1066),.q(_w_6230));
  spl2 g1311_s_0(.a(n1311),.q0(n1311_0),.q1(n1311_1));
  and_bi g282(.a(G94_4),.b(G168_6),.q(n282));
  bfr _b_5600(.a(_w_7025),.q(_w_7026));
  bfr _b_3467(.a(_w_4892),.q(_w_4893));
  bfr _b_6572(.a(_w_7997),.q(_w_7998));
  bfr _b_4500(.a(_w_5925),.q(_w_5926));
  bfr _b_5054(.a(_w_6479),.q(_w_6480));
  and_bi g236(.a(G128_4),.b(G168_0),.q(n236));
  bfr _b_2258(.a(_w_3683),.q(_w_3684));
  bfr _b_2970(.a(_w_4395),.q(_w_4396));
  or_bb g281(.a(G169_7),.b(G94_0),.q(n281));
  and_bb g993(.a(G176_21),.b(n233_1),.q(n993));
  spl4L G100_s_3(.a(G100_2),.q0(G100_12),.q1(G100_13),.q2(G100_14),.q3(G100_15));
  spl4L G107_s_0(.a(G107),.q0(_w_4701),.q1(G107_1),.q2(G107_2),.q3(_w_4702));
  and_bi g584(.a(G172_0),.b(n583),.q(n584));
  bfr _b_2894(.a(_w_4319),.q(_w_4320));
  and_bb g1231(.a(G102_9),.b(G128_12),.q(n1231));
  spl4L g397_s_0(.a(n397),.q0(n397_0),.q1(n397_1),.q2(n397_2),.q3(n397_3));
  bfr _b_5480(.a(_w_6905),.q(_w_6906));
  and_bi g520(.a(G111_1),.b(G109_9),.q(n520));
  spl4L G126_s_0(.a(G126),.q0(_w_3638),.q1(G126_1),.q2(G126_2),.q3(_w_3639));
  and_bi g1001(.a(n1000),.b(G5243_1),.q(n1001));
  bfr _b_3726(.a(_w_5151),.q(G160_2));
  and_bb g517(.a(G103_9),.b(G96_9),.q(n517));
  and_bi g1332(.a(n1326),.b(n1331),.q(n1332));
  and_bb g638(.a(G2_4),.b(n402_1),.q(_w_4738));
  bfr _b_7472(.a(_w_8897),.q(_w_8898));
  or_bb g834(.a(n832),.b(n833),.q(n834));
  spl4L G174_s_3(.a(G174_2),.q0(G174_12),.q1(G174_13),.q2(G174_14),.q3(G174_15));
  and_bb g207(.a(G163_12),.b(_w_7409),.q(_w_4703));
  and_bi g265(.a(G166_5),.b(G121_6),.q(n265));
  bfr _b_4018(.a(_w_5443),.q(_w_5444));
  spl2 G84_s_0(.a(_w_8807),.q0(G84_0),.q1(G84_1));
  bfr _b_5439(.a(_w_6864),.q(_w_6865));
  and_bi g1092(.a(G158_14),.b(G5288_4),.q(_w_6284));
  bfr _b_3400(.a(_w_4825),.q(_w_4826));
  and_bb g278(.a(n268_0),.b(n277_0),.q(n278));
  bfr _b_5090(.a(_w_6515),.q(_w_6516));
  spl4L G174_s_1(.a(G174_0),.q0(G174_4),.q1(_w_5463),.q2(_w_5464),.q3(G174_7));
  bfr _b_7521(.a(G91),.q(_w_8947));
  spl4L g381_s_0(.a(n381),.q0(n381_0),.q1(n381_1),.q2(n381_2),.q3(n381_3));
  bfr _b_2309(.a(_w_3734),.q(G174_24));
  bfr _b_3427(.a(_w_4852),.q(_w_4853));
  bfr _b_6652(.a(_w_8077),.q(_w_8078));
  and_bi g276(.a(n275),.b(G149_1),.q(n276));
  bfr _b_2298(.a(_w_3723),.q(_w_3724));
  and_bb g1056(.a(G39_0),.b(n586_9),.q(n1056));
  bfr _b_7085(.a(_w_8510),.q(_w_8511));
  bfr _b_2751(.a(_w_4176),.q(_w_4177));
  and_bi g557(.a(n556_0),.b(G176_35),.q(_w_4705));
  and_bb g636(.a(_w_7939),.b(n552_20),.q(_w_4706));
  or_bb g1034(.a(n1032),.b(n1033),.q(n1034));
  bfr _b_5294(.a(_w_6719),.q(_w_6720));
  and_bb g655(.a(n653_0),.b(n654),.q(n655));
  bfr _b_2122(.a(_w_3547),.q(_w_3548));
  bfr _b_3493(.a(_w_4918),.q(_w_4919));
  or_bb g225(.a(G100_21),.b(G119_0),.q(n225));
  bfr _b_3357(.a(_w_4782),.q(n439_0));
  and_bi g1003(.a(n1002),.b(G5262_1),.q(G5289));
  bfr _b_5591(.a(_w_7016),.q(_w_7017));
  spl2 G41_s_0(.a(_w_7628),.q0(G41_0),.q1(G41_1));
  bfr _b_2651(.a(_w_4076),.q(_w_4077));
  bfr _b_7141(.a(_w_8566),.q(_w_8567));
  and_bi g1101(.a(G158_12),.b(G5287_4),.q(_w_4707));
  bfr _b_2321(.a(_w_3746),.q(G175_6));
  and_bi g261(.a(G121_4),.b(G168_4),.q(n261));
  bfr _b_5739(.a(_w_7164),.q(_w_7165));
  and_bb g273(.a(G126_5),.b(G167_5),.q(n273));
  spl4L g630_s_1(.a(n630_2),.q0(n630_4),.q1(n630_5),.q2(n630_6),.q3(n630_7));
  bfr _b_4584(.a(_w_6009),.q(_w_6010));
  bfr _b_5126(.a(_w_6551),.q(_w_6552));
  bfr _b_3035(.a(_w_4460),.q(_w_4461));
  bfr _b_3989(.a(_w_5414),.q(_w_5415));
  and_bb g1163(.a(G64_7),.b(n1162),.q(G5309));
  and_bb g676(.a(_w_7973),.b(n552_15),.q(n676));
  bfr _b_6801(.a(_w_8226),.q(_w_8227));
  and_bi g601(.a(n600_0),.b(G176_41),.q(n601));
  bfr _b_7385(.a(_w_8810),.q(_w_8811));
  bfr _b_5722(.a(_w_7147),.q(_w_7148));
  and_bi g729(.a(n424_2),.b(n728_0),.q(n729));
  and_bi g1443(.a(_w_7510),.b(G177_6),.q(_w_6070));
  bfr _b_3286(.a(_w_4711),.q(_w_4712));
  bfr _b_6253(.a(_w_7678),.q(_w_7679));
  and_bi g271(.a(n269),.b(n270),.q(n271));
  spl4L g605_s_0(.a(G5253_0),.q0(_w_4709),.q1(G5253_1),.q2(G5253_2),.q3(G5253_3));
  or_bb g1215(.a(G100_15),.b(G121_10),.q(n1215));
  bfr _b_3309(.a(_w_4734),.q(n459));
  bfr _b_5475(.a(_w_6900),.q(_w_6901));
  bfr _b_4486(.a(_w_5911),.q(_w_5912));
  spl4L g990_s_0(.a(G5287_0),.q0(_w_4717),.q1(G5287_1),.q2(G5287_2),.q3(G5287_3));
  and_bb g379(.a(G135_2),.b(n378_0),.q(n379));
  bfr _b_5599(.a(_w_7024),.q(_w_7025));
  spl2 g786_s_0(.a(n786),.q0(n786_0),.q1(n786_1));
  bfr _b_3104(.a(_w_4529),.q(_w_4530));
  bfr _b_5407(.a(_w_6832),.q(_w_6833));
  and_bi g1404(.a(G98_17),.b(G96_13),.q(n1404));
  spl2 g1201_s_0(.a(n1201),.q0(n1201_0),.q1(n1201_1));
  bfr _b_2546(.a(_w_3971),.q(G5248));
  or_bb g703(.a(G125_1),.b(n474_1),.q(_w_4372));
  bfr _b_3164(.a(_w_4589),.q(_w_4590));
  spl2 g365_s_0(.a(n365),.q0(n365_0),.q1(_w_4133));
  or_bb g268(.a(n263),.b(n267),.q(_w_4725));
  and_bi g459(.a(n458_0),.b(n457_0),.q(_w_4734));
  and_bb g1020(.a(n1017),.b(n1019),.q(n1020));
  bfr _b_3375(.a(_w_4800),.q(_w_4801));
  and_bi g1360(.a(n1350_0),.b(n1359_0),.q(n1360));
  bfr _b_3115(.a(_w_4540),.q(_w_4541));
  bfr _b_6211(.a(_w_7636),.q(_w_7637));
  and_bi g196(.a(_w_8944),.b(G163_7),.q(_w_4742));
  bfr _b_7137(.a(_w_8562),.q(_w_8563));
  spl2 g1431_s_0(.a(n1431),.q0(n1431_0),.q1(n1431_1));
  bfr _b_4915(.a(_w_6340),.q(_w_6341));
  and_bb g1112(.a(G159_12),.b(n1111),.q(n1112));
  or_bb g310(.a(G109_0),.b(G169_10),.q(n310));
  bfr _b_2655(.a(_w_4080),.q(n403_3));
  bfr _b_7047(.a(_w_8472),.q(_w_8473));
  bfr _b_2734(.a(_w_4159),.q(_w_4160));
  bfr _b_3307(.a(_w_4732),.q(_w_4733));
  spl2 G15_s_0(.a(_w_6566),.q0(G15_0),.q1(G15_1));
  and_bb g366(.a(n356_0),.b(n365_0),.q(n366));
  and_bi g394(.a(n393_0),.b(n392_0),.q(n394));
  bfr _b_4180(.a(_w_5605),.q(_w_5606));
  and_bi g205(.a(G66_3),.b(n204),.q(G5233));
  bfr _b_7443(.a(_w_8868),.q(_w_8869));
  bfr _b_2778(.a(_w_4203),.q(_w_4204));
  bfr _b_7018(.a(_w_8443),.q(_w_8444));
  or_bb g462(.a(n460),.b(n461),.q(_w_4745));
  bfr _b_2296(.a(_w_3721),.q(G173_24));
  and_bi g609(.a(n435_2),.b(n607_1),.q(n609));
  and_bi g976(.a(G177_4),.b(n975),.q(n976));
  bfr _b_3456(.a(_w_4881),.q(n197));
  bfr _b_5320(.a(_w_6745),.q(_w_6746));
  and_bb g294(.a(G167_7),.b(G90_5),.q(n294));
  or_bb g307(.a(n302),.b(n306),.q(_w_4750));
  spl2 g645_s_0(.a(n645),.q0(n645_0),.q1(n645_1));
  bfr _b_7416(.a(G85),.q(_w_8842));
  and_bb g389(.a(G105_7),.b(G124_20),.q(n389));
  bfr _b_3480(.a(_w_4905),.q(_w_4906));
  and_bb g1004(.a(_w_7757),.b(n552_10),.q(_w_4438));
  or_bb g1281(.a(n380_2),.b(n386_6),.q(n1281));
  bfr _b_3290(.a(_w_4715),.q(_w_4716));
  spl2 G162_s_0(.a(_w_6907),.q0(G162_0),.q1(G162_1));
  and_bi g568(.a(G177_28),.b(n567),.q(n568));
  or_bb g251(.a(G100_18),.b(G130_0),.q(n251));
  and_bb g1259(.a(n1250_1),.b(n1257_1),.q(n1259));
  and_bi g704(.a(n703),.b(n702),.q(n704));
  spl2 G21_s_0(.a(_w_7205),.q0(G21_0),.q1(G21_1));
  spl2 G128_s_1(.a(G128_1),.q0(G128_4),.q1(G128_5));
  and_bi g791(.a(n790),.b(n565_1),.q(n791));
  or_bb g325(.a(n323),.b(n324),.q(n325));
  bfr _b_7516(.a(_w_8941),.q(_w_8908));
  and_bi g738(.a(n737_0),.b(n725_0),.q(n738));
  bfr _b_2251(.a(_w_3676),.q(G158_2));
  bfr _b_7388(.a(_w_8813),.q(_w_8814));
  bfr _b_2854(.a(_w_4279),.q(_w_4280));
  bfr _b_1943(.a(_w_3368),.q(G147_2));
  spl4L G175_s_2(.a(G175_2),.q0(G175_7),.q1(G175_8),.q2(G175_9),.q3(G175_10));
  and_bi g411(.a(_w_8946),.b(G124_11),.q(n411));
  or_bb g346(.a(n341),.b(n345),.q(n346));
  bfr _b_5817(.a(_w_7242),.q(_w_7243));
  bfr _b_2117(.a(_w_3542),.q(_w_3543));
  bfr _b_4124(.a(_w_5549),.q(_w_5550));
  bfr _b_1951(.a(_w_3376),.q(_w_3377));
  bfr _b_1981(.a(_w_3406),.q(_w_3407));
  spl4L G160_s_6(.a(G160_19),.q0(_w_4769),.q1(G160_25),.q2(G160_26),.q3(G160_27));
  bfr _b_5162(.a(_w_6587),.q(_w_6588));
  or_bb g1155(.a(G160_8),.b(G5290_5),.q(_w_6302));
  and_bb g919(.a(G64_20),.b(n918),.q(G5278));
  bfr _b_3692(.a(_w_5117),.q(_w_5118));
  or_bb g504(.a(n491_0),.b(n503_0),.q(n504));
  bfr _b_4465(.a(_w_5890),.q(_w_5891));
  bfr _b_4781(.a(_w_6206),.q(G5293_0));
  and_bb g1072(.a(G17_1),.b(n630_8),.q(n1072));
  or_bb g566(.a(G176_37),.b(n565_0),.q(_w_4784));
  or_bb g954(.a(n950),.b(n953),.q(_w_4785));
  or_ii g195(.a(_w_7449),.b(G5221_6),.q(_w_4786));
  or_bb g469(.a(n467),.b(n468),.q(_w_4823));
  bfr _b_3737(.a(_w_5162),.q(_w_5163));
  and_bi g253(.a(n251),.b(n252),.q(n253));
  or_bb g640(.a(n399_2),.b(n639),.q(n640));
  bfr _b_5014(.a(_w_6439),.q(_w_6438));
  and_bi g210(.a(G66_4),.b(n209),.q(G5234));
  and_ii g978(.a(n973),.b(n977),.q(_w_5616));
  and_bb g1018(.a(G176_27),.b(n307_1),.q(n1018));
  and_bi g581(.a(n473_1),.b(n580),.q(G5251_0));
  bfr _b_3696(.a(_w_5121),.q(_w_5122));
  bfr _b_4999(.a(G12),.q(_w_6424));
  bfr _b_7104(.a(_w_8529),.q(_w_8530));
  bfr _b_2244(.a(_w_3669),.q(G158_17));
  and_bi g1441(.a(n552_5),.b(_w_7821),.q(_w_4842));
  bfr _b_6865(.a(_w_8290),.q(_w_8291));
  bfr _b_4718(.a(_w_6143),.q(_w_6144));
  bfr _b_6843(.a(_w_8268),.q(_w_8269));
  bfr _b_3964(.a(_w_5389),.q(_w_5390));
  spl4L G145_s_0(.a(_w_6541),.q0(G145_0),.q1(G145_1),.q2(_w_4854),.q3(_w_4857));
  and_bb g425(.a(G140_2),.b(n424_0),.q(n425));
  and_bi g1356(.a(G98_13),.b(G92_13),.q(n1356));
  or_bb g354(.a(n352),.b(n353),.q(n354));
  bfr _b_3124(.a(_w_4549),.q(_w_4550));
  and_bi g1199(.a(n1198_0),.b(n451_4),.q(n1199));
  and_bb g258(.a(n250_0),.b(n257),.q(n258));
  bfr _b_3123(.a(_w_4548),.q(_w_4549));
  bfr _b_1941(.a(_w_3366),.q(G5261));
  and_bb g446(.a(G123_18),.b(G126_7),.q(n446));
  or_bb g456(.a(n454),.b(n455),.q(_w_4668));
  and_bi g479(.a(n478_0),.b(n477_0),.q(n479));
  and_bi g1400(.a(G96_11),.b(G101_17),.q(n1400));
  bfr _b_6899(.a(_w_8324),.q(_w_8325));
  and_bb g995(.a(n992),.b(n994),.q(n995));
  spl3L G144_s_1(.a(G144_3),.q0(G144_4),.q1(G144_5),.q2(G144_6));
  bfr _b_3655(.a(_w_5080),.q(_w_5081));
  bfr _b_2306(.a(_w_3731),.q(_w_3732));
  bfr _b_2820(.a(_w_4245),.q(G172_3));
  bfr _b_6856(.a(_w_8281),.q(_w_8282));
  spl4L G176_s_4(.a(G176_3),.q0(G176_16),.q1(G176_17),.q2(G176_18),.q3(G176_19));
  and_bi g249(.a(n247),.b(n248),.q(_w_4875));
  or_bb g266(.a(n264),.b(n265),.q(n266));
  bfr _b_2740(.a(_w_4165),.q(_w_4166));
  bfr _b_7505(.a(_w_8930),.q(_w_8931));
  and_bb g197(.a(G163_8),.b(_w_8671),.q(_w_4881));
  and_bi g246(.a(n244),.b(n245),.q(_w_4882));
  bfr _b_7080(.a(_w_8505),.q(_w_8506));
  spl2 g1009_s_1(.a(G5290_3),.q0(G5290_4),.q1(G5290_5));
  and_bi g486(.a(G117_6),.b(G119_6),.q(n486));
  bfr _b_4657(.a(_w_6082),.q(_w_6083));
  bfr _b_6140(.a(_w_7565),.q(_w_7566));
  or_bb g938(.a(G160_20),.b(G5259_5),.q(n938));
  and_bb g1382(.a(G102_14),.b(G107_12),.q(n1382));
  bfr _b_4544(.a(_w_5969),.q(_w_5970));
  spl4L g815_s_1(.a(n815_2),.q0(n815_4),.q1(n815_5),.q2(n815_6),.q3(n815_7));
  and_bi g315(.a(G166_10),.b(G109_6),.q(n315));
  or_bb g530(.a(n528),.b(n529),.q(n530));
  spl4L G98_s_1(.a(G98_0),.q0(_w_4977),.q1(_w_4978),.q2(G98_6),.q3(G98_7));
  bfr _b_3339(.a(_w_4764),.q(_w_4765));
  and_bi g286(.a(G166_7),.b(G94_6),.q(n286));
  bfr _b_6953(.a(_w_8378),.q(_w_8379));
  and_bi g711(.a(n710_0),.b(n692_0),.q(n711));
  or_bb g1445(.a(G173_6),.b(n1444_0),.q(n1445));
  and_bi g350(.a(n348),.b(n349),.q(n350));
  bfr _b_3229(.a(_w_4654),.q(n472));
  or_bb g521(.a(n519),.b(n520),.q(n521));
  bfr _b_2213(.a(_w_3638),.q(G126_0));
  spl3L G102_s_1(.a(G102_0),.q0(G102_4),.q1(G102_5),.q2(G102_6));
  bfr _b_5636(.a(_w_7061),.q(_w_7062));
  and_bb g239(.a(G128_5),.b(G167_0),.q(n239));
  bfr _b_3764(.a(_w_5189),.q(_w_5190));
  bfr _b_2289(.a(_w_3714),.q(_w_3715));
  bfr _b_2802(.a(_w_4227),.q(_w_4228));
  spl3L g537_s_1(.a(n537_3),.q0(n537_4),.q1(_w_4631),.q2(_w_4634));
  spl2 g500_s_0(.a(n500),.q0(n500_0),.q1(n500_1));
  bfr _b_2229(.a(_w_3654),.q(_w_3655));
  and_bi g485(.a(n483),.b(n484),.q(n485));
  and_ii g1009(.a(n1004),.b(n1008),.q(_w_6149));
  or_bb g1337(.a(n1335),.b(n1336),.q(n1337));
  bfr _b_2608(.a(_w_4033),.q(_w_4034));
  and_bi g608(.a(n607_0),.b(n435_1),.q(n608));
  spl3L g445_s_0(.a(n445),.q0(n445_0),.q1(n445_1),.q2(n445_2));
  and_bi g1268(.a(n1267),.b(n388_2),.q(n1268));
  or_bb g497(.a(n495),.b(n496),.q(n497));
  and_bb g1079(.a(n1076),.b(n1078),.q(_w_6271));
  and_bi g1159(.a(G73_1),.b(n813_10),.q(n1159));
  spl4L G160_s_2(.a(G160_1),.q0(G160_8),.q1(G160_9),.q2(G160_10),.q3(G160_11));
  and_bi g496(.a(n494_1),.b(G121_9),.q(n496));
  or_bb g882(.a(n880),.b(n881),.q(n882));
  bfr _b_2333(.a(_w_3758),.q(_w_3759));
  bfr _b_5037(.a(_w_6462),.q(_w_6463));
  or_bb g269(.a(G126_0),.b(G169_6),.q(n269));
  bfr _b_2527(.a(_w_3952),.q(_w_3953));
  spl2 g1184_s_0(.a(n1184),.q0(n1184_0),.q1(n1184_1));
  bfr _b_2770(.a(_w_4195),.q(_w_4196));
  bfr _b_3705(.a(_w_5130),.q(_w_5131));
  bfr _b_5732(.a(_w_7157),.q(_w_7158));
  and_bb g756(.a(n645_1),.b(n755),.q(n756));
  bfr _b_2118(.a(_w_3543),.q(_w_3544));
  spl4L g469_s_2(.a(n469_3),.q0(n469_7),.q1(n469_8),.q2(_w_3450),.q3(_w_3451));
  or_bb g287(.a(n285),.b(n286),.q(n287));
  spl3L G172_s_1(.a(G172_1),.q0(G172_4),.q1(G172_5),.q2(_w_4943));
  bfr _b_4824(.a(_w_6249),.q(_w_6250));
  bfr _b_7221(.a(_w_8646),.q(_w_8647));
  or_bb g1478(.a(n1476),.b(n1477),.q(_w_4945));
  and_bi g396(.a(_w_6396),.b(G124_15),.q(n396));
  bfr _b_5960(.a(_w_7385),.q(_w_7386));
  bfr _b_3198(.a(_w_4623),.q(_w_4624));
  bfr _b_6306(.a(_w_7731),.q(_w_7732));
  or_bb g393(.a(G138_4),.b(n391_1),.q(n393));
  and_bi g741(.a(n740_0),.b(n722_0),.q(n741));
  and_bb g889(.a(G86_0),.b(n804_1),.q(n889));
  spl2 g381_s_1(.a(n381_3),.q0(n381_4),.q1(n381_5));
  bfr _b_6113(.a(_w_7538),.q(_w_7539));
  and_bb g567(.a(G176_38),.b(n243_1),.q(n567));
  bfr _b_4771(.a(_w_6196),.q(_w_6197));
  and_ii g605(.a(n592),.b(n604),.q(_w_4946));
  spl4L G176_s_2(.a(G176_1),.q0(G176_8),.q1(_w_3412),.q2(G176_10),.q3(G176_11));
  bfr _b_4110(.a(_w_5535),.q(_w_5536));
  or_bb g737(.a(n735),.b(n736),.q(n737));
  and_bi g623(.a(G177_24),.b(n622),.q(n623));
  or_bb g1276(.a(n1275_0),.b(n643_1),.q(_w_6166));
  bfr _b_5761(.a(_w_7186),.q(_w_7187));
  bfr _b_3247(.a(_w_4672),.q(_w_4673));
  bfr _b_4126(.a(_w_5551),.q(_w_5552));
  bfr _b_2064(.a(_w_3489),.q(G94_3));
  and_bi g226(.a(G119_1),.b(G101_5),.q(_w_5331));
  or_bi g506(.a(n505),.b(n504),.q(_w_4953));
  bfr _b_3656(.a(_w_5081),.q(_w_5082));
  bfr _b_5108(.a(_w_6533),.q(_w_6534));
  or_bb g900(.a(n896),.b(n899),.q(_w_4975));
  and_bi g447(.a(G127_0),.b(G123_17),.q(n447));
  and_bb g1094(.a(G159_10),.b(n1093),.q(n1094));
  and_bb g1016(.a(_w_7184),.b(n552_8),.q(_w_6181));
  and_bi g1095(.a(n1094),.b(n1092),.q(_w_4976));
  spl2 g1257_s_0(.a(n1257),.q0(n1257_0),.q1(n1257_1));
  bfr _b_2735(.a(_w_4160),.q(_w_4161));
  or_bb g189(.a(n187),.b(n188),.q(n189));
  bfr _b_5529(.a(_w_6954),.q(_w_6955));
  and_bb g1151(.a(G84_1),.b(n815_9),.q(n1151));
  spl2 G42_s_0(.a(_w_7661),.q0(G42_0),.q1(G42_1));
  bfr _b_2917(.a(_w_4342),.q(_w_4343));
  and_bb g539(.a(n537_0),.b(n538),.q(n539));
  bfr _b_6809(.a(_w_8234),.q(_w_8235));
  bfr _b_3392(.a(_w_4817),.q(_w_4818));
  spl4L g650_s_0(.a(G5257_0),.q0(_w_3710),.q1(G5257_1),.q2(G5257_2),.q3(G5257_3));
  bfr _b_4997(.a(G119),.q(_w_6423));
  bfr _b_7412(.a(_w_8837),.q(_w_8838));
  bfr _b_5559(.a(_w_6984),.q(_w_6985));
  and_bb g454(.a(G117_5),.b(G123_16),.q(n454));
  bfr _b_5621(.a(_w_7046),.q(_w_7047));
  or_bb g233(.a(n228),.b(n232),.q(n233));
  and_bb g457(.a(G145_2),.b(n456_0),.q(_w_4979));
  bfr _b_4872(.a(_w_6297),.q(G123_14));
  bfr _b_2161(.a(_w_3586),.q(_w_3587));
  bfr _b_4560(.a(_w_5985),.q(_w_5986));
  bfr _b_5139(.a(_w_6564),.q(_w_6565));
  and_bi g682(.a(n681),.b(n679),.q(_w_5628));
  spl2 g594_s_0(.a(n594),.q0(n594_0),.q1(_w_4982));
  and_bi g213(.a(G5221_10),.b(n212),.q(n213));
  spl2 g420_s_0(.a(n420),.q0(n420_0),.q1(n420_1));
  or_bb g653(.a(n537_2),.b(n652),.q(n653));
  bfr _b_3724(.a(_w_5149),.q(G160_1));
  spl4L G166_s_3(.a(G166_3),.q0(G166_11),.q1(G166_12),.q2(G166_13),.q3(G166_14));
  or_bb g277(.a(n272),.b(n276),.q(_w_4992));
  bfr _b_2256(.a(_w_3681),.q(n544_1));
  bfr _b_4189(.a(_w_5614),.q(n370));
  and_bi g223(.a(n222),.b(G145_1),.q(n223));
  spl2 G6_s_0(.a(_w_8080),.q0(G6_0),.q1(G6_1));
  and_bb g1145(.a(G64_9),.b(n1144),.q(_w_5003));
  and_bi g564(.a(n442_4),.b(n563),.q(_w_5004));
  bfr _b_6978(.a(_w_8403),.q(_w_8404));
  bfr _b_4912(.a(_w_6337),.q(_w_6338));
  and_bb g308(.a(n298_0),.b(n307_0),.q(n308));
  bfr _b_7442(.a(_w_8867),.q(_w_8868));
  spl2 G85_s_0(.a(_w_8841),.q0(G85_0),.q1(G85_1));
  or_bb g442(.a(n440),.b(n441),.q(_w_5473));
  bfr _b_1986(.a(_w_3411),.q(G176_14));
  and_bb g404(.a(G124_4),.b(G88_5),.q(n404));
  bfr _b_5518(.a(_w_6943),.q(_w_6944));
  or_bb g1017(.a(G176_26),.b(n769_1),.q(n1017));
  bfr _b_4474(.a(_w_5899),.q(_w_5900));
  and_bi g621(.a(n620_0),.b(G176_45),.q(n621));
  and_bi g293(.a(G143_0),.b(n292),.q(n293));
  bfr _b_6146(.a(_w_7571),.q(_w_7572));
  or_bb g380(.a(G135_4),.b(n378_1),.q(n380));
  or_bb g1195(.a(n1193),.b(n1194),.q(n1195));
  bfr _b_5373(.a(_w_6798),.q(_w_6799));
  bfr _b_3405(.a(_w_4830),.q(n896));
  and_bi g678(.a(n677),.b(n666_1),.q(n678));
  and_bi g217(.a(G117_1),.b(G101_4),.q(n217));
  and_bi g1316(.a(n415_5),.b(n426_3),.q(n1316));
  spl3L g476_s_0(.a(n476),.q0(n476_0),.q1(n476_1),.q2(n476_2));
  and_bi g339(.a(G88_1),.b(G100_17),.q(n339));
  spl4L G160_s_4(.a(G160_3),.q0(_w_5038),.q1(_w_5040),.q2(_w_5042),.q3(G160_19));
  or_bb g750(.a(n427_1),.b(n744_1),.q(n750));
  spl3L G141_s_1(.a(G141_3),.q0(_w_3645),.q1(G141_5),.q2(G141_6));
  and_bi g257(.a(n256_0),.b(n253_0),.q(_w_5043));
  or_bb g575(.a(G176_39),.b(n574_0),.q(_w_5051));
  bfr _b_3457(.a(_w_4882),.q(_w_4883));
  bfr _b_5854(.a(_w_7279),.q(_w_7280));
  and_bb g793(.a(n610_1),.b(n792),.q(n793));
  bfr _b_3411(.a(_w_4836),.q(_w_4837));
  spl3L g427_s_0(.a(n427),.q0(n427_0),.q1(_w_5052),.q2(_w_5063));
  bfr _b_6091(.a(_w_7516),.q(_w_7517));
  or_bb g1267(.a(n381_5),.b(n387_3),.q(n1267));
  bfr _b_3943(.a(_w_5368),.q(_w_5369));
  and_bb g1041(.a(G42_1),.b(n586_7),.q(n1041));
  bfr _b_4327(.a(_w_5752),.q(_w_5753));
  or_ii g186(.a(G5221_1),.b(_w_8184),.q(_w_5074));
  bfr _b_7438(.a(_w_8863),.q(_w_8864));
  and_bb g433(.a(G148_2),.b(n432_0),.q(_w_5110));
  and_bi g922(.a(G161_6),.b(n921),.q(n922));
  bfr _b_2315(.a(_w_3740),.q(G174_17));
  or_bb g565(.a(n445_1),.b(n564),.q(_w_5113));
  and_bb g751(.a(n427_2),.b(n744_2),.q(n751));
  and_bi g188(.a(_w_7453),.b(G163_4),.q(n188));
  or_bb g1116(.a(n1114),.b(n1115),.q(n1116));
  bfr _b_4273(.a(_w_5698),.q(G99_1));
  bfr _b_2262(.a(_w_3687),.q(_w_3688));
  bfr _b_2828(.a(_w_4253),.q(_w_4254));
  bfr _b_2995(.a(_w_4420),.q(_w_4421));
  bfr _b_7268(.a(_w_8693),.q(_w_8694));
  spl4L g542_s_0(.a(n542),.q0(n542_0),.q1(_w_4625),.q2(_w_4626),.q3(n542_3));
  and_bi g1234(.a(n1233),.b(G150_6),.q(n1234));
  and_bb g280(.a(n234_0),.b(n279),.q(_w_5117));
  or_bb g632(.a(G174_25),.b(G175_5),.q(n632));
  bfr _b_5897(.a(_w_7322),.q(_w_7323));
  bfr _b_4840(.a(_w_6265),.q(_w_6266));
  bfr _b_4675(.a(_w_6100),.q(_w_6101));
  or_bb g335(.a(n333),.b(n334),.q(n335));
  bfr _b_6220(.a(_w_7645),.q(_w_7646));
  bfr _b_6131(.a(_w_7556),.q(_w_7557));
  bfr _b_3797(.a(_w_5222),.q(_w_5223));
  and_bi g242(.a(n241),.b(G150_1),.q(n242));
  bfr _b_6915(.a(_w_8340),.q(_w_8341));
  and_bi g371(.a(_w_8952),.b(G124_25),.q(n371));
  spl2 g477_s_0(.a(n477),.q0(n477_0),.q1(_w_5138));
  bfr _b_2598(.a(_w_4023),.q(_w_4024));
  and_bi g727(.a(_w_6407),.b(G124_5),.q(n727));
  spl4L G160_s_0(.a(_w_6848),.q0(_w_5146),.q1(_w_5148),.q2(_w_5150),.q3(G160_3));
  spl2 g692_s_0(.a(n692),.q0(n692_0),.q1(n692_1));
  and_bi g524(.a(n522),.b(n523),.q(n524));
  bfr _b_3133(.a(_w_4558),.q(n535));
  bfr _b_5375(.a(_w_6800),.q(_w_6801));
  bfr _b_2178(.a(_w_3603),.q(_w_3604));
  and_bb g1219(.a(G102_8),.b(G121_12),.q(n1219));
  or_bb g1301(.a(n409_4),.b(n421_4),.q(n1301));
  and_bb g367(.a(n347),.b(n366),.q(n367));
  bfr _b_7323(.a(_w_8748),.q(_w_8749));
  spl4L g561_s_0(.a(G5248_0),.q0(_w_3963),.q1(G5248_1),.q2(G5248_2),.q3(G5248_3));
  bfr _b_4215(.a(_w_5640),.q(_w_5641));
  bfr _b_5178(.a(_w_6603),.q(_w_6604));
  bfr _b_4699(.a(_w_6124),.q(_w_6125));
  and_bb g538(.a(n375_1),.b(n400_1),.q(n538));
  and_bi g1392(.a(G98_16),.b(G105_13),.q(n1392));
  bfr _b_4330(.a(_w_5755),.q(_w_5756));
  and_bi g862(.a(G175_7),.b(n861),.q(n862));
  bfr _b_6368(.a(_w_7793),.q(_w_7794));
  and_bi g1038(.a(G172_10),.b(n1037),.q(n1038));
  bfr _b_2610(.a(_w_4035),.q(_w_4036));
  or_bb g235(.a(G128_0),.b(G169_0),.q(_w_5153));
  and_bb g562(.a(_w_8036),.b(n552_25),.q(n562));
  or_bb g688(.a(n462_3),.b(n472_5),.q(n688));
  bfr _b_2769(.a(_w_4194),.q(_w_4195));
  bfr _b_4366(.a(_w_5791),.q(_w_5792));
  bfr _b_4923(.a(_w_6348),.q(n1247));
  bfr _b_5800(.a(_w_7225),.q(_w_7226));
  or_bb g918(.a(n914),.b(n917),.q(_w_5154));
  bfr _b_5630(.a(_w_7055),.q(_w_7056));
  or_bb g1126(.a(n1122),.b(n1125),.q(n1126));
  bfr _b_6394(.a(_w_7819),.q(_w_7820));
  bfr _b_6138(.a(_w_7563),.q(_w_7564));
  bfr _b_3888(.a(_w_5313),.q(_w_5314));
  and_bb g212(.a(G163_14),.b(_w_7447),.q(_w_5155));
  spl2 g268_s_0(.a(n268),.q0(n268_0),.q1(_w_5254));
  bfr _b_2203(.a(_w_3628),.q(_w_3629));
  and_bb g368(.a(n328),.b(n367),.q(n368));
  and_bb g1246(.a(n1235_1),.b(n1244_1),.q(n1246));
  bfr _b_3978(.a(_w_5403),.q(_w_5404));
  bfr _b_6179(.a(_w_7604),.q(_w_7605));
  or_bb g719(.a(n717),.b(n718),.q(n719));
  bfr _b_6429(.a(_w_7854),.q(_w_7855));
  and_bi g214(.a(n213),.b(n211),.q(_w_5196));
  bfr _b_4707(.a(_w_6132),.q(_w_6133));
  bfr _b_7432(.a(_w_8857),.q(_w_8858));
  bfr _b_2320(.a(_w_3745),.q(_w_3746));
  and_bi g1361(.a(n1359_1),.b(n1350_1),.q(n1361));
  or_bb g406(.a(n404),.b(n405),.q(_w_5256));
  and_bi g215(.a(G66_5),.b(n214),.q(G5235));
  bfr _b_7321(.a(_w_8746),.q(_w_8747));
  bfr _b_5519(.a(_w_6944),.q(_w_6945));
  or_bi g183(.a(_w_6915),.b(G11_0),.q(_w_5258));
  bfr _b_3961(.a(_w_5386),.q(_w_5387));
  bfr _b_3994(.a(_w_5419),.q(_w_5420));
  bfr _b_3539(.a(_w_4964),.q(_w_4965));
  bfr _b_4520(.a(_w_5945),.q(_w_5946));
  bfr _b_2989(.a(_w_4414),.q(_w_4415));
  bfr _b_2219(.a(_w_3644),.q(G135_2));
  or_bb g243(.a(n238),.b(n242),.q(_w_4597));
  bfr _b_2564(.a(_w_3989),.q(_w_3990));
  bfr _b_5748(.a(_w_7173),.q(_w_7174));
  and_bi g262(.a(n260),.b(n261),.q(n262));
  bfr _b_2284(.a(_w_3709),.q(n425_3));
  or_bb g852(.a(G174_24),.b(G5257_2),.q(n852));
  bfr _b_7172(.a(_w_8597),.q(_w_8598));
  and_bi g360(.a(G138_0),.b(n359),.q(n360));
  and_bb g323(.a(G167_10),.b(G96_5),.q(n323));
  bfr _b_3203(.a(_w_4628),.q(_w_4629));
  and_bb g1277(.a(n1275_1),.b(n643_2),.q(_w_5330));
  or_bb g1286(.a(n1268_1),.b(n375_5),.q(n1286));
  and_bb g1328(.a(n1311_1),.b(n1327),.q(n1328));
  and_bb g666(.a(n387_1),.b(n665_0),.q(n666));
  or_bb g1125(.a(n1123),.b(n1124),.q(n1125));
  bfr _b_6405(.a(_w_7830),.q(_w_7831));
  or_bb g439(.a(G150_2),.b(n438_0),.q(_w_4681));
  spl2 g289_s_0(.a(n289),.q0(n289_0),.q1(_w_5332));
  and_bb g892(.a(G64_23),.b(n891),.q(G5275));
  and_bi g435(.a(n434_0),.b(n433_0),.q(n435));
  bfr _b_2523(.a(_w_3948),.q(_w_3949));
  bfr _b_5934(.a(_w_7359),.q(_w_7360));
  or_bb g594(.a(n449_1),.b(n593),.q(n594));
  and_bi g1375(.a(n1374_0),.b(n1362_0),.q(n1375));
  bfr _b_2898(.a(_w_4323),.q(G5216));
  and_bb g410(.a(G124_12),.b(G90_7),.q(n410));
  and_bi g1284(.a(n1282_1),.b(n653_2),.q(n1284));
  bfr _b_4230(.a(_w_5655),.q(_w_5656));
  bfr _b_6455(.a(_w_7880),.q(_w_7881));
  bfr _b_6280(.a(_w_7705),.q(_w_7706));
  bfr _b_5720(.a(_w_7145),.q(_w_7146));
  bfr _b_2609(.a(_w_4034),.q(_w_4035));
  and_bi g673(.a(G177_21),.b(n672),.q(_w_5335));
  and_bb g413(.a(G143_2),.b(n412_0),.q(_w_5337));
  bfr _b_7314(.a(G82),.q(_w_8740));
  and_bi g336(.a(n335),.b(G139_1),.q(n336));
  and_bi g856(.a(G14_1),.b(n632_1),.q(n856));
  bfr _b_2876(.a(_w_4301),.q(_w_4302));
  bfr _b_6105(.a(_w_7530),.q(_w_7531));
  bfr _b_1944(.a(_w_3369),.q(_w_3370));
  bfr _b_2530(.a(_w_3955),.q(_w_3956));
  spl4L G107_s_3(.a(G107_3),.q0(G107_10),.q1(G107_11),.q2(G107_12),.q3(G107_13));
  bfr _b_2847(.a(_w_4272),.q(_w_4273));
  spl4L G96_s_0(.a(G96),.q0(_w_5338),.q1(G96_1),.q2(G96_2),.q3(_w_5339));
  bfr _b_3684(.a(_w_5109),.q(G5220));
  and_bi g1336(.a(n1334_1),.b(n1332_1),.q(n1336));
  and_bb g639(.a(n398_1),.b(n537_1),.q(n639));
  bfr _b_6104(.a(G39),.q(_w_7530));
  bfr _b_5620(.a(_w_7045),.q(_w_7046));
  bfr _b_3916(.a(_w_5341),.q(_w_5342));
  bfr _b_2211(.a(_w_3636),.q(n421_2));
  spl2 G129_s_0(.a(_w_6434),.q0(G129_0),.q1(_w_5340));
  bfr _b_7011(.a(_w_8436),.q(_w_8437));
  bfr _b_6478(.a(_w_7903),.q(_w_7904));
  or_bb g859(.a(n855),.b(n858),.q(_w_5376));
  bfr _b_5328(.a(_w_6753),.q(_w_6754));
  and_bi g694(.a(_w_6441),.b(G123_5),.q(n694));
  bfr _b_5712(.a(_w_7137),.q(_w_7138));
  and_bi g306(.a(n305),.b(G144_1),.q(n306));
  bfr _b_5554(.a(_w_6979),.q(_w_6980));
  and_bi g706(.a(n442_6),.b(n704_1),.q(n706));
  and_bb g651(.a(_w_8015),.b(n552_17),.q(n651));
  bfr _b_6749(.a(_w_8174),.q(_w_8175));
  or_bb g356(.a(n351),.b(n355),.q(_w_4933));
  bfr _b_3368(.a(_w_4793),.q(_w_4794));
  or_bb g710(.a(n708),.b(n709),.q(_w_5388));
  bfr _b_4854(.a(_w_6279),.q(G5274));
  spl2 G79_s_0(.a(_w_8637),.q0(G79_0),.q1(G79_1));
  and_ii g561(.a(n553),.b(n560),.q(_w_5396));
  or_bb g929(.a(G160_22),.b(G5260_5),.q(n929));
  bfr _b_3117(.a(_w_4542),.q(G5244_0));
  or_bb g424(.a(n422),.b(n423),.q(n424));
  bfr _b_2218(.a(_w_3643),.q(_w_3644));
  and_bi g513(.a(n512_0),.b(n509_0),.q(n513));
  and_bi g815(.a(G160_25),.b(G161_5),.q(n815));
  spl2 G39_s_0(.a(_w_7529),.q0(G39_0),.q1(G39_1));
  bfr _b_6664(.a(_w_8089),.q(_w_8090));
  or_bb g1307(.a(n1303_1),.b(n1305_1),.q(n1307));
  and_bi g1229(.a(n1227),.b(n1228),.q(n1229));
  and_bb g748(.a(n409_2),.b(n746_1),.q(n748));
  and_bb g700(.a(n695_1),.b(n698_1),.q(n700));
  bfr _b_3634(.a(_w_5059),.q(_w_5060));
  bfr _b_2155(.a(_w_3580),.q(_w_3581));
  bfr _b_3570(.a(_w_4995),.q(_w_4996));
  spl4L G100_s_4(.a(G100_3),.q0(G100_16),.q1(G100_17),.q2(G100_18),.q3(G100_19));
  bfr _b_2362(.a(_w_3787),.q(G113_6));
  bfr _b_4887(.a(_w_6312),.q(_w_6313));
  bfr _b_7485(.a(_w_8910),.q(_w_8911));
  bfr _b_2193(.a(_w_3618),.q(_w_3619));
  and_bi g800(.a(G159_0),.b(n799),.q(n800));
  bfr _b_5676(.a(_w_7101),.q(_w_7102));
  bfr _b_4069(.a(_w_5494),.q(G176_45));
  and_bb g619(.a(n451_2),.b(n617_1),.q(n619));
  and_bb g1180(.a(n1176_0),.b(n1179_0),.q(n1180));
  bfr _b_4092(.a(_w_5517),.q(_w_5518));
  or_bi g551(.a(n469_1),.b(n472_1),.q(_w_5408));
  bfr _b_6605(.a(_w_8030),.q(_w_8031));
  bfr _b_4410(.a(_w_5835),.q(n725));
  bfr _b_5999(.a(_w_7424),.q(_w_7425));
  bfr _b_4897(.a(_w_6322),.q(_w_6323));
  or_bb g1289(.a(n402_2),.b(n640_2),.q(n1289));
  spl4L G176_s_13(.a(G176_19),.q0(G176_50),.q1(_w_5433),.q2(G176_52),.q3(G176_53));
  bfr _b_7399(.a(_w_8824),.q(_w_8825));
  bfr _b_6692(.a(_w_8117),.q(_w_8118));
  bfr _b_2513(.a(_w_3938),.q(_w_3939));
  bfr _b_6790(.a(_w_8215),.q(_w_8216));
  spl4L g1303_s_0(.a(n1303),.q0(_w_5436),.q1(_w_5438),.q2(n1303_2),.q3(n1303_3));
  bfr _b_4532(.a(_w_5957),.q(_w_5958));
  bfr _b_6334(.a(_w_7759),.q(_w_7760));
  and_bi g1334(.a(n1333),.b(n401_1),.q(_w_4921));
  and_bi g614(.a(n613),.b(n611),.q(_w_5440));
  bfr _b_6020(.a(G30),.q(_w_7446));
  bfr _b_2441(.a(_w_3866),.q(_w_3867));
  bfr _b_3191(.a(_w_4616),.q(_w_4617));
  or_bb g507(.a(G88_6),.b(G90_8),.q(n507));
  bfr _b_7227(.a(_w_8652),.q(_w_8653));
  bfr _b_3904(.a(_w_5329),.q(n204));
  and_bi g362(.a(G166_14),.b(G105_6),.q(n362));
  bfr _b_3355(.a(_w_4780),.q(_w_4781));
  bfr _b_4992(.a(G117),.q(_w_6418));
  spl4L G113_s_0(.a(_w_6409),.q0(G113_0),.q1(G113_1),.q2(G113_2),.q3(G113_3));
  spl2 G130_s_1(.a(G130_3),.q0(G130_4),.q1(G130_5));
  spl2 G165_s_0(.a(G165),.q0(G165_0),.q1(G165_1));
  or_bb g1399(.a(G100_7),.b(G96_10),.q(n1399));
  bfr _b_5333(.a(_w_6758),.q(_w_6759));
  bfr _b_3141(.a(_w_4566),.q(_w_4567));
  and_bi g312(.a(n310),.b(n311),.q(n312));
  and_bb g905(.a(n902),.b(n904),.q(_w_5442));
  bfr _b_3803(.a(_w_5228),.q(n214));
  bfr _b_6601(.a(_w_8026),.q(_w_8027));
  and_bi g1218(.a(G147_5),.b(n1217),.q(n1218));
  bfr _b_6679(.a(_w_8104),.q(_w_8105));
  bfr _b_4115(.a(_w_5540),.q(_w_5541));
  and_bi g313(.a(G135_0),.b(n312),.q(n313));
  spl4L G176_s_11(.a(G176_17),.q0(G176_42),.q1(_w_5493),.q2(G176_44),.q3(_w_5494));
  and_bi g1283(.a(n653_1),.b(n1282_0),.q(n1283));
  bfr _b_2839(.a(_w_4264),.q(G161_3));
  spl2 g675_s_1(.a(G5259_3),.q0(G5259_4),.q1(G5259_5));
  bfr _b_6399(.a(_w_7824),.q(_w_7825));
  bfr _b_2779(.a(_w_4204),.q(_w_4205));
  and_bb g576(.a(G176_40),.b(n318_1),.q(n576));
  bfr _b_7220(.a(_w_8645),.q(_w_8646));
  bfr _b_5513(.a(_w_6938),.q(_w_6939));
  bfr _b_2346(.a(_w_3771),.q(_w_3772));
  bfr _b_3332(.a(_w_4757),.q(_w_4758));
  inv inv_G113(.a(G113_6),.q(G5194));
  bfr _b_1995(.a(_w_3420),.q(G176_9));
  bfr _b_2129(.a(_w_3554),.q(_w_3555));
  and_bi g390(.a(_w_6398),.b(G124_17),.q(_w_5455));
  bfr _b_2528(.a(_w_3953),.q(_w_3954));
  or_bb g827(.a(n823),.b(n826),.q(_w_5456));
  or_bb g316(.a(n314),.b(n315),.q(n316));
  and_bi g489(.a(n488_0),.b(n485_0),.q(n489));
  or_bb g478(.a(G147_4),.b(n476_1),.q(_w_5460));
  spl2 g1235_s_0(.a(n1235),.q0(n1235_0),.q1(n1235_1));
  and_bi g948(.a(G160_4),.b(G5254_5),.q(n948));
  bfr _b_4374(.a(_w_5799),.q(_w_5800));
  or_bb g391(.a(n389),.b(n390),.q(n391));
  or_bb g1271(.a(n1268_0),.b(n1270),.q(n1271));
  bfr _b_7060(.a(_w_8485),.q(_w_8486));
  bfr _b_4455(.a(_w_5880),.q(n753));
  bfr _b_7150(.a(_w_8575),.q(_w_8576));
  spl4L G92_s_2(.a(G92_2),.q0(G92_6),.q1(G92_7),.q2(G92_8),.q3(G92_9));
  or_bb g357(.a(G105_0),.b(G169_14),.q(n357));
  bfr _b_4647(.a(_w_6072),.q(_w_6073));
  bfr _b_3554(.a(_w_4979),.q(n457));
  bfr _b_6698(.a(_w_8123),.q(_w_8124));
  bfr _b_4503(.a(_w_5928),.q(_w_5929));
  and_bi g1364(.a(G94_11),.b(G101_14),.q(n1364));
  and_bi g558(.a(G176_36),.b(n253_1),.q(n558));
  or_bb g1211(.a(n1209),.b(n1210),.q(n1211));
  or_bb g434(.a(G148_4),.b(n432_1),.q(_w_5470));
  bfr _b_2927(.a(_w_4352),.q(G5285));
  bfr _b_4947(.a(_w_6372),.q(_w_6373));
  or_bb g1304(.a(n1298_1),.b(n425_3),.q(n1304));
  bfr _b_5869(.a(_w_7294),.q(_w_7295));
  bfr _b_5136(.a(_w_6561),.q(_w_6559));
  bfr _b_3718(.a(_w_5143),.q(_w_5144));
  and_bb g328(.a(n318_0),.b(n327_0),.q(n328));
  bfr _b_4648(.a(_w_6073),.q(_w_6074));
  or_bb g329(.a(G107_0),.b(G169_12),.q(n329));
  spl4L G90_s_0(.a(G90),.q0(_w_3373),.q1(G90_1),.q2(G90_2),.q3(_w_3374));
  bfr _b_2008(.a(_w_3433),.q(_w_3434));
  bfr _b_6878(.a(_w_8303),.q(_w_8304));
  bfr _b_4266(.a(_w_5691),.q(_w_5692));
  bfr _b_4958(.a(_w_6383),.q(_w_6384));
  inv inv_G66(.a(G66_6),.q(G5193));
  spl2 G68_s_0(.a(_w_8262),.q0(G68_0),.q1(G68_1));
  bfr _b_7398(.a(_w_8823),.q(_w_8824));
  bfr _b_7351(.a(_w_8776),.q(_w_8777));
  bfr _b_6117(.a(_w_7542),.q(_w_7543));
  bfr _b_4835(.a(_w_6260),.q(_w_6261));
  bfr _b_5017(.a(_w_6442),.q(_w_6441));
  and_bi g1379(.a(G107_11),.b(G101_15),.q(n1379));
  bfr _b_3452(.a(_w_4877),.q(_w_4878));
  bfr _b_5684(.a(_w_7109),.q(_w_7110));
  bfr _b_4490(.a(_w_5915),.q(_w_5916));
  and_bi g331(.a(n329),.b(n330),.q(n331));
  and_bb g616(.a(_w_7875),.b(n552_21),.q(n616));
  and_ii g1027(.a(n1022),.b(n1026),.q(_w_6202));
  bfr _b_4556(.a(_w_5981),.q(n202));
  bfr _b_6479(.a(_w_7904),.q(_w_7905));
  inv inv_G127(.a(G127_1),.q(G5197));
  and_bi g603(.a(G177_26),.b(n602),.q(_w_5482));
  and_bb g376(.a(G109_7),.b(G124_24),.q(n376));
  and_bi g583(.a(G173_27),.b(G5248_1),.q(n583));
  bfr _b_2420(.a(_w_3845),.q(_w_3846));
  bfr _b_2069(.a(_w_3494),.q(_w_3495));
  bfr _b_7051(.a(_w_8476),.q(_w_8477));
  bfr _b_3678(.a(_w_5103),.q(_w_5104));
  bfr _b_5030(.a(_w_6455),.q(_w_6456));
  spl4L G109_s_2(.a(G109_2),.q0(G109_6),.q1(_w_5484),.q2(G109_8),.q3(G109_9));
  bfr _b_4146(.a(_w_5571),.q(_w_5572));
  and_bi g343(.a(G102_7),.b(G88_4),.q(n343));
  bfr _b_5395(.a(_w_6820),.q(_w_6821));
  bfr _b_3757(.a(_w_5182),.q(_w_5183));
  bfr _b_4764(.a(_w_6189),.q(n1028));
  bfr _b_5726(.a(_w_7151),.q(_w_7152));
  and_bi g906(.a(G70_0),.b(n802_5),.q(n906));
  and_bi g1263(.a(n1262),.b(n1208),.q(n1263));
  or_bb g911(.a(G158_16),.b(G5258_4),.q(_w_5485));
  bfr _b_3860(.a(_w_5285),.q(_w_5286));
  and_bi g1007(.a(G177_12),.b(n1006),.q(_w_5486));
  bfr _b_4777(.a(_w_6202),.q(_w_6203));
  bfr _b_3418(.a(_w_4843),.q(_w_4844));
  spl4L G177_s_0(.a(_w_7104),.q0(_w_5495),.q1(_w_5496),.q2(_w_5501),.q3(G177_3));
  bfr _b_3146(.a(_w_4571),.q(_w_4572));
  spl4L G98_s_0(.a(_w_8955),.q0(G98_0),.q1(G98_1),.q2(G98_2),.q3(G98_3));
  bfr _b_5499(.a(_w_6924),.q(_w_6925));
  inv inv_G165(.a(G165_1),.q(_w_5502));
  bfr _b_5740(.a(_w_7165),.q(_w_7166));
  bfr _b_3646(.a(_w_5071),.q(_w_5072));
  bfr _b_5050(.a(_w_6475),.q(_w_6476));
  spl4L g552_s_3(.a(n552_2),.q0(n552_12),.q1(n552_13),.q2(n552_14),.q3(n552_15));
  or_bb g1371(.a(n1366),.b(n1370),.q(n1371));
  bfr _b_3680(.a(_w_5105),.q(_w_5106));
  and_bb g191(.a(_w_6436),.b(G163_5),.q(n191));
  bfr _b_6991(.a(_w_8416),.q(_w_8417));
  spl3L G159_s_1(.a(G159_1),.q0(G159_4),.q1(G159_5),.q2(_w_3654));
  and_bi g877(.a(G174_4),.b(G5249_2),.q(n877));
  bfr _b_3808(.a(_w_5233),.q(_w_5234));
  or_bb g728(.a(n726),.b(n727),.q(n728));
  bfr _b_2517(.a(_w_3942),.q(_w_3943));
  and_bi g679(.a(n678_0),.b(G176_53),.q(_w_5578));
  bfr _b_5794(.a(_w_7219),.q(_w_7220));
  bfr _b_5751(.a(_w_7176),.q(_w_7177));
  spl4L G128_s_3(.a(G128_3),.q0(G128_10),.q1(G128_11),.q2(G128_12),.q3(G128_13));
  or_bb g1214(.a(n1212),.b(n1213),.q(n1214));
  and_bi g739(.a(n725_1),.b(n737_1),.q(n739));
  bfr _b_5938(.a(_w_7363),.q(_w_7364));
  bfr _b_3436(.a(_w_4861),.q(_w_4862));
  or_bb g275(.a(n273),.b(n274),.q(n275));
  and_bi g502(.a(n500_1),.b(n497_1),.q(n502));
  bfr _b_7446(.a(_w_8871),.q(_w_8872));
  bfr _b_2214(.a(_w_3639),.q(G126_3));
  bfr _b_2641(.a(_w_4066),.q(_w_4067));
  and_bi g351(.a(G137_0),.b(n350),.q(n351));
  bfr _b_4571(.a(_w_5996),.q(_w_5997));
  bfr _b_2428(.a(_w_3853),.q(_w_3854));
  bfr _b_6229(.a(_w_7654),.q(_w_7655));
  bfr _b_2257(.a(_w_3682),.q(_w_3683));
  bfr _b_3252(.a(_w_4677),.q(n461));
  bfr _b_3168(.a(_w_4593),.q(_w_4594));
  and_bi g355(.a(n354),.b(G137_1),.q(n355));
  bfr _b_2590(.a(_w_4015),.q(_w_4016));
  bfr _b_2450(.a(_w_3875),.q(_w_3876));
  and_bi g1055(.a(n1054),.b(n1052),.q(_w_5585));
  and_bi g1476(.a(G79_1),.b(n813_11),.q(n1476));
  bfr _b_6828(.a(_w_8253),.q(_w_8254));
  spl3L G150_s_1(.a(G150_3),.q0(_w_6172),.q1(G150_5),.q2(G150_6));
  bfr _b_3945(.a(_w_5370),.q(_w_5371));
  bfr _b_5661(.a(_w_7086),.q(_w_7087));
  and_bi g974(.a(G5251_6),.b(G176_5),.q(_w_5586));
  and_bi g1390(.a(G138_5),.b(n1389),.q(n1390));
  bfr _b_3877(.a(_w_5302),.q(_w_5303));
  bfr _b_3227(.a(_w_4652),.q(_w_4653));
  and_bi g982(.a(G177_15),.b(n981),.q(_w_5587));
  and_bb g361(.a(G105_5),.b(G167_13),.q(n361));
  bfr _b_2135(.a(_w_3560),.q(_w_3561));
  and_bi g749(.a(n747),.b(n748),.q(n749));
  and_bb g1256(.a(n1252_1),.b(n1254_1),.q(n1256));
  bfr _b_2829(.a(_w_4254),.q(n1474));
  bfr _b_5517(.a(_w_6942),.q(_w_6943));
  bfr _b_3426(.a(_w_4851),.q(_w_4852));
  bfr _b_5918(.a(G26),.q(_w_7344));
  bfr _b_4715(.a(_w_6140),.q(n356_1));
  or_bb g1395(.a(n1390),.b(n1394),.q(n1395));
  bfr _b_6910(.a(_w_8335),.q(_w_8336));
  bfr _b_2690(.a(_w_4115),.q(_w_4116));
  or_bb g598(.a(n479_1),.b(n597_0),.q(n598));
  and_bi g254(.a(G166_4),.b(G148_0),.q(n254));
  spl2 g789_s_0(.a(n789),.q0(n789_0),.q1(n789_1));
  or_bb g224(.a(n219),.b(n223),.q(n224));
  bfr _b_3179(.a(_w_4604),.q(_w_4605));
  spl4L g632_s_0(.a(n632),.q0(n632_0),.q1(n632_1),.q2(n632_2),.q3(n632_3));
  bfr _b_7059(.a(_w_8484),.q(_w_8485));
  bfr _b_6264(.a(_w_7689),.q(_w_7690));
  and_bb g1006(.a(G176_23),.b(n346_1),.q(n1006));
  and_bb g369(.a(n309),.b(n368),.q(_w_5595));
  and_bb g370(.a(G124_14),.b(G96_7),.q(_w_5614));
  bfr _b_7466(.a(_w_8891),.q(_w_8892));
  bfr _b_1988(.a(_w_3413),.q(_w_3414));
  and_bi g1073(.a(G18_1),.b(n632_8),.q(n1073));
  bfr _b_2606(.a(_w_4031),.q(_w_4032));
  bfr _b_4966(.a(G10),.q(_w_6392));
  bfr _b_5708(.a(_w_7133),.q(_w_7134));
  or_ii g194(.a(G5221_5),.b(n193),.q(_w_5629));
  bfr _b_3549(.a(_w_4974),.q(G5242_0));
  and_bb g840(.a(G26_0),.b(n586_5),.q(n840));
  bfr _b_5923(.a(_w_7348),.q(_w_7349));
  bfr _b_4583(.a(_w_6008),.q(_w_6009));
  bfr _b_2893(.a(_w_4318),.q(n1297));
  bfr _b_4847(.a(_w_6272),.q(_w_6273));
  or_bb g494(.a(n492),.b(n493),.q(n494));
  bfr _b_4080(.a(_w_5505),.q(_w_5506));
  spl2 G156_s_0(.a(_w_6704),.q0(G156_0),.q1(_w_5687));
  and_bi g381(.a(n380_0),.b(n379_0),.q(n381));
  bfr _b_7258(.a(_w_8683),.q(_w_8684));
  bfr _b_4183(.a(_w_5608),.q(_w_5609));
  spl2 G99_s_0(.a(_w_8956),.q0(G99_0),.q1(_w_5693));
  and_bb g812(.a(n809),.b(n811),.q(_w_5699));
  spl4L G172_s_2(.a(G172_2),.q0(G172_7),.q1(G172_8),.q2(G172_9),.q3(G172_10));
  and_bi g674(.a(n673),.b(n671),.q(n674));
  or_bb g1248(.a(n1226_0),.b(n1247_0),.q(n1248));
  bfr _b_6965(.a(_w_8390),.q(_w_8391));
  and_bb g585(.a(n582),.b(n584),.q(_w_5700));
  bfr _b_6247(.a(_w_7672),.q(_w_7673));
  and_bi g445(.a(n439_0),.b(n444_0),.q(n445));
  spl4L G158_s_4(.a(G158_3),.q0(_w_3666),.q1(_w_3668),.q2(_w_3670),.q3(G158_19));
  and_bi g1178(.a(n464_5),.b(n469_10),.q(n1178));
  bfr _b_2276(.a(_w_3701),.q(_w_3702));
  and_bi g255(.a(G148_1),.b(G169_4),.q(n255));
  bfr _b_3029(.a(_w_4454),.q(_w_4455));
  bfr _b_7099(.a(_w_8524),.q(_w_8525));
  and_bi g1308(.a(n1307),.b(n1306),.q(n1308));
  bfr _b_3828(.a(_w_5253),.q(G130_2));
  and_bi g1110(.a(G158_10),.b(G5286_4),.q(_w_5702));
  bfr _b_4770(.a(_w_6195),.q(G5311));
  or_bb g1058(.a(n1056),.b(n1057),.q(n1058));
  and_bi g1044(.a(G173_12),.b(G5286_1),.q(_w_5703));
  or_bb g1059(.a(n1055),.b(n1058),.q(_w_5704));
  bfr _b_4489(.a(_w_5914),.q(_w_5915));
  bfr _b_7095(.a(_w_8520),.q(_w_8521));
  and_bi g383(.a(_w_6400),.b(G124_21),.q(n383));
  bfr _b_6082(.a(_w_7507),.q(_w_7508));
  bfr _b_2985(.a(_w_4410),.q(_w_4411));
  or_bb g384(.a(n382),.b(n383),.q(n384));
  bfr _b_6612(.a(_w_8037),.q(_w_8038));
  and_bi g267(.a(n266),.b(G147_1),.q(n267));
  bfr _b_2988(.a(_w_4413),.q(_w_4414));
  and_bi g208(.a(G5221_9),.b(n207),.q(n208));
  and_bi g203(.a(G5221_8),.b(n202),.q(n203));
  spl4L g409_s_0(.a(n409),.q0(_w_5708),.q1(_w_5713),.q2(_w_5726),.q3(n409_3));
  or_bb g1035(.a(n1031),.b(n1034),.q(_w_6208));
  and_bb g386(.a(G139_4),.b(n384_1),.q(n386));
  spl2 G4_s_0(.a(_w_7562),.q0(G4_0),.q1(G4_1));
  and_bi g1192(.a(n1191),.b(n1189),.q(_w_5739));
  and_bi g387(.a(n385_0),.b(n386_0),.q(n387));
  bfr _b_2363(.a(_w_3788),.q(_w_3789));
  bfr _b_2435(.a(_w_3860),.q(_w_3861));
  and_bb g956(.a(G170_0),.b(G5251_2),.q(n956));
  bfr _b_3328(.a(_w_4753),.q(_w_4754));
  bfr _b_2035(.a(_w_3460),.q(n465_1));
  bfr _b_3685(.a(_w_5110),.q(_w_5111));
  and_bb g395(.a(G103_7),.b(G124_16),.q(n395));
  spl3L g643_s_0(.a(n643),.q0(n643_0),.q1(_w_5743),.q2(_w_5744));
  bfr _b_5883(.a(_w_7308),.q(_w_7309));
  or_bb g527(.a(n525),.b(n526),.q(_w_5745));
  bfr _b_2057(.a(_w_3482),.q(n459_1));
  bfr _b_2052(.a(_w_3477),.q(n462_3));
  bfr _b_5202(.a(_w_6627),.q(_w_6628));
  and_bb g229(.a(G102_5),.b(G119_2),.q(_w_6291));
  bfr _b_2281(.a(_w_3706),.q(_w_3707));
  and_bi g670(.a(n668),.b(n669),.q(n670));
  and_bi g237(.a(n235),.b(n236),.q(n237));
  bfr _b_2016(.a(_w_3441),.q(G142_2));
  bfr _b_2496(.a(_w_3921),.q(_w_3922));
  and_ii g650(.a(n636),.b(n649),.q(_w_4985));
  and_bi g1241(.a(G98_11),.b(G126_13),.q(n1241));
  and_bi g400(.a(n398_0),.b(n399_0),.q(n400));
  bfr _b_5579(.a(G173),.q(_w_7005));
  bfr _b_2114(.a(_w_3539),.q(_w_3540));
  or_bb g590(.a(n587),.b(n589),.q(n590));
  bfr _b_3532(.a(_w_4957),.q(_w_4958));
  or_bb g337(.a(n332),.b(n336),.q(_w_5748));
  bfr _b_2278(.a(_w_3703),.q(n425_2));
  or_bb g344(.a(n342),.b(n343),.q(n344));
  bfr _b_2587(.a(_w_4012),.q(_w_4013));
  bfr _b_4078(.a(_w_5503),.q(_w_5504));
  spl3L G132_s_0(.a(_w_6440),.q0(G132_0),.q1(G132_1),.q2(G132_2));
  or_bb g1461(.a(n1459),.b(n1460),.q(_w_5749));
  and_bb g402(.a(n388_0),.b(n401_0),.q(n402));
  bfr _b_1963(.a(_w_3388),.q(_w_3389));
  or_bb g763(.a(n761),.b(n762),.q(n763));
  bfr _b_1956(.a(_w_3381),.q(_w_3382));
  bfr _b_7296(.a(_w_8721),.q(_w_8722));
  bfr _b_3806(.a(_w_5231),.q(_w_5232));
  bfr _b_5028(.a(_w_6453),.q(_w_6454));
  bfr _b_2000(.a(_w_3425),.q(_w_3426));
  and_bi g698(.a(n696),.b(n697),.q(n698));
  spl4L g1447_s_0(.a(n1447),.q0(n1447_0),.q1(n1447_1),.q2(n1447_2),.q3(n1447_3));
  bfr _b_2465(.a(_w_3890),.q(_w_3891));
  bfr _b_2781(.a(_w_4206),.q(_w_4207));
  or_bb g980(.a(G176_7),.b(n786_1),.q(n980));
  and_bi g340(.a(n338),.b(n339),.q(n340));
  and_bi g814(.a(G81_1),.b(n813_0),.q(n814));
  bfr _b_5185(.a(_w_6610),.q(_w_6611));
  and_bi g662(.a(n661),.b(n659),.q(n662));
  bfr _b_4000(.a(_w_5425),.q(_w_5426));
  bfr _b_5687(.a(_w_7112),.q(_w_7113));
  and_bb g484(.a(G113_5),.b(G115_5),.q(n484));
  spl3L g233_s_0(.a(n233),.q0(n233_0),.q1(_w_5752),.q2(n233_2));
  spl2 g561_s_1(.a(G5248_3),.q0(G5248_4),.q1(G5248_5));
  bfr _b_4024(.a(_w_5449),.q(_w_5450));
  bfr _b_2049(.a(_w_3474),.q(_w_3475));
  bfr _b_2356(.a(_w_3781),.q(_w_3782));
  spl4L G119_s_0(.a(_w_6422),.q0(_w_4708),.q1(G119_1),.q2(G119_2),.q3(G119_3));
  and_bb g985(.a(_w_7778),.b(n552_12),.q(_w_5759));
  bfr _b_4275(.a(_w_5700),.q(n585));
  or_bb g414(.a(G143_4),.b(n412_1),.q(_w_5766));
  bfr _b_5849(.a(_w_7274),.q(_w_7275));
  or_bb g850(.a(n848),.b(n849),.q(n850));
  bfr _b_2886(.a(_w_4311),.q(_w_4312));
  and_bb g416(.a(G124_10),.b(G92_7),.q(n416));
  bfr _b_4929(.a(G1),.q(_w_6355));
  and_bi g525(.a(G105_8),.b(G107_8),.q(n525));
  bfr _b_7091(.a(_w_8516),.q(_w_8517));
  bfr _b_2698(.a(_w_4123),.q(_w_4124));
  and_bi g712(.a(n692_1),.b(n710_1),.q(n712));
  or_ii g190(.a(G5221_4),.b(n189),.q(_w_5770));
  bfr _b_6293(.a(_w_7718),.q(_w_7719));
  and_bb g431(.a(n403_0),.b(n430_0),.q(_w_5805));
  or_bb g418(.a(n416),.b(n417),.q(n418));
  or_bb g1251(.a(n224_2),.b(n233_2),.q(_w_5826));
  bfr _b_5681(.a(_w_7106),.q(_w_7107));
  or_bb g1462(.a(n1458),.b(n1461),.q(_w_5827));
  bfr _b_4003(.a(_w_5428),.q(_w_5429));
  bfr _b_6945(.a(_w_8370),.q(_w_8371));
  and_bi g423(.a(_w_8950),.b(G124_7),.q(n423));
  bfr _b_2926(.a(_w_4351),.q(_w_4352));
  bfr _b_7315(.a(_w_8740),.q(_w_8741));
  spl2 g658_s_0(.a(n658),.q0(n658_0),.q1(n658_1));
  spl2 g1254_s_0(.a(n1254),.q0(n1254_0),.q1(n1254_1));
  bfr _b_2929(.a(_w_4354),.q(n1149));
  and_bi g364(.a(n363),.b(G138_1),.q(n364));
  or_bb g920(.a(G160_24),.b(G5257_5),.q(n920));
  and_bi g471(.a(_w_6415),.b(G123_9),.q(_w_5828));
  bfr _b_5371(.a(_w_6796),.q(_w_6797));
  and_bi g1063(.a(n1062),.b(n1060),.q(_w_6228));
  bfr _b_3347(.a(_w_4772),.q(_w_4773));
  and_bb g428(.a(n421_0),.b(n427_0),.q(n428));
  spl2 g734_s_0(.a(n734),.q0(n734_0),.q1(n734_1));
  bfr _b_4698(.a(_w_6123),.q(G5290));
  or_bb g432(.a(G123_14),.b(G125_0),.q(n432));
  or_bb g851(.a(n847),.b(n850),.q(_w_5829));
  bfr _b_4094(.a(_w_5519),.q(_w_5520));
  bfr _b_6940(.a(_w_8365),.q(_w_8332));
  or_bb g720(.a(n716_0),.b(n719_0),.q(n720));
  and_bi g961(.a(n960),.b(n956),.q(n961));
  bfr _b_2433(.a(_w_3858),.q(_w_3859));
  bfr _b_2956(.a(_w_4381),.q(G5258_0));
  bfr _b_7511(.a(_w_8936),.q(_w_8937));
  bfr _b_6430(.a(_w_7855),.q(_w_7856));
  and_bi g641(.a(n640_0),.b(n375_2),.q(n641));
  bfr _b_6409(.a(_w_7834),.q(_w_7835));
  and_bb g726(.a(G111_2),.b(G124_6),.q(n726));
  bfr _b_2939(.a(_w_4364),.q(_w_4365));
  bfr _b_4644(.a(_w_6069),.q(G5286_0));
  and_bi g933(.a(G72_1),.b(n813_4),.q(n933));
  and_bi g730(.a(n728_1),.b(n424_3),.q(n730));
  bfr _b_7422(.a(_w_8847),.q(_w_8848));
  bfr _b_3213(.a(_w_4638),.q(_w_4639));
  or_bb g597(.a(n453_1),.b(n596),.q(n597));
  and_bb g754(.a(n658_1),.b(n753),.q(n754));
  and_ii g1015(.a(n1010),.b(n1014),.q(_w_5837));
  spl4L g675_s_0(.a(G5259_0),.q0(_w_5838),.q1(G5259_1),.q2(G5259_2),.q3(G5259_3));
  or_bb g699(.a(n695_0),.b(n698_0),.q(n699));
  bfr _b_3499(.a(_w_4924),.q(_w_4925));
  and_bi g733(.a(n372_3),.b(n406_3),.q(n733));
  or_bb g734(.a(n732),.b(n733),.q(n734));
  bfr _b_6688(.a(G60),.q(_w_8114));
  bfr _b_2138(.a(_w_3563),.q(_w_3564));
  spl4L g813_s_1(.a(n813_2),.q0(n813_4),.q1(n813_5),.q2(n813_6),.q3(n813_7));
  spl2 g663_s_1(.a(G5258_3),.q0(G5258_4),.q1(G5258_5));
  bfr _b_4165(.a(_w_5590),.q(_w_5591));
  and_bi g735(.a(n734_0),.b(n731_0),.q(n735));
  bfr _b_5491(.a(G17),.q(_w_6917));
  and_bi g1184(.a(n1183),.b(n1174),.q(_w_6317));
  bfr _b_2301(.a(_w_3726),.q(G173_17));
  bfr _b_3125(.a(_w_4550),.q(_w_4551));
  spl2 g1282_s_0(.a(n1282),.q0(n1282_0),.q1(n1282_1));
  bfr _b_5947(.a(_w_7372),.q(_w_7373));
  bfr _b_5316(.a(_w_6741),.q(_w_6742));
  or_bb g740(.a(n738),.b(n739),.q(n740));
  bfr _b_2637(.a(_w_4062),.q(G127_1));
  bfr _b_2873(.a(_w_4298),.q(_w_4299));
  bfr _b_3333(.a(_w_4758),.q(_w_4759));
  or_bb g1470(.a(n1466),.b(n1469),.q(n1470));
  bfr _b_2085(.a(_w_3510),.q(G140_2));
  or_bb g1183(.a(n1182),.b(n773_7),.q(n1183));
  bfr _b_4850(.a(_w_6275),.q(n947));
  and_ii g743(.a(n741),.b(n742),.q(_w_5845));
  spl2 G70_s_0(.a(_w_8332),.q0(G70_0),.q1(G70_1));
  spl4L G107_s_2(.a(G107_2),.q0(G107_6),.q1(_w_6104),.q2(G107_8),.q3(G107_9));
  bfr _b_3689(.a(_w_5114),.q(_w_5115));
  or_bb g818(.a(n812),.b(n817),.q(_w_5866));
  or_bb g747(.a(n409_1),.b(n746_0),.q(n747));
  bfr _b_6849(.a(_w_8274),.q(_w_8275));
  and_bb g1355(.a(G102_12),.b(G92_12),.q(n1355));
  bfr _b_3654(.a(_w_5079),.q(_w_5080));
  and_bb g855(.a(n852),.b(n854),.q(n855));
  and_bi g475(.a(G123_7),.b(G121_7),.q(_w_5868));
  and_bi g752(.a(n750),.b(n751),.q(n752));
  bfr _b_2482(.a(_w_3907),.q(_w_3908));
  spl4L g463_s_0(.a(n463),.q0(n463_0),.q1(_w_5869),.q2(_w_5876),.q3(_w_5878));
  bfr _b_5493(.a(_w_6918),.q(_w_6919));
  and_bi g977(.a(n976),.b(n974),.q(_w_5879));
  spl4L G163_s_3(.a(G163_3),.q0(G163_11),.q1(G163_12),.q2(G163_13),.q3(G163_14));
  bfr _b_6017(.a(_w_7442),.q(_w_7443));
  bfr _b_3261(.a(_w_4686),.q(_w_4687));
  bfr _b_3535(.a(_w_4960),.q(_w_4961));
  and_bb g1302(.a(n409_5),.b(n421_5),.q(n1302));
  bfr _b_2183(.a(_w_3608),.q(_w_3609));
  spl4L G167_s_3(.a(G167_3),.q0(G167_10),.q1(G167_11),.q2(G167_12),.q3(G167_13));
  and_bb g755(.a(n670_1),.b(n754),.q(n755));
  bfr _b_3673(.a(_w_5098),.q(_w_5099));
  and_bb g758(.a(n749_0),.b(n757),.q(_w_5882));
  spl2 g478_s_0(.a(n478),.q0(n478_0),.q1(_w_4914));
  bfr _b_2777(.a(_w_4202),.q(_w_4203));
  spl3L g386_s_1(.a(n386_3),.q0(_w_3369),.q1(n386_5),.q2(n386_6));
  bfr _b_4062(.a(_w_5487),.q(_w_5488));
  and_bb g759(.a(n428_1),.b(n744_4),.q(n759));
  bfr _b_3237(.a(_w_4662),.q(n979));
  spl4L g586_s_2(.a(n586_3),.q0(n586_8),.q1(n586_9),.q2(n586_10),.q3(n586_11));
  spl2 g752_s_0(.a(n752),.q0(n752_0),.q1(n752_1));
  bfr _b_2830(.a(_w_4255),.q(n1469));
  and_bb g460(.a(G119_5),.b(G123_4),.q(n460));
  bfr _b_5856(.a(_w_7281),.q(_w_7282));
  and_bi g1239(.a(G149_5),.b(n1238),.q(n1239));
  bfr _b_2329(.a(_w_3754),.q(_w_3755));
  bfr _b_5335(.a(_w_6760),.q(_w_6761));
  spl4L g996_s_0(.a(G5288_0),.q0(_w_4065),.q1(G5288_1),.q2(G5288_2),.q3(G5288_3));
  and_bi g766(.a(n765),.b(n764),.q(n766));
  and_bb g1103(.a(G159_11),.b(n1102),.q(n1103));
  bfr _b_5241(.a(_w_6666),.q(_w_6667));
  and_bi g320(.a(G96_4),.b(G168_10),.q(n320));
  or_bb g1236(.a(G100_4),.b(G126_10),.q(n1236));
  bfr _b_5596(.a(_w_7021),.q(_w_7022));
  or_bb g397(.a(n395),.b(n396),.q(_w_5883));
  or_bb g1023(.a(G176_28),.b(n752_1),.q(n1023));
  bfr _b_2195(.a(_w_3620),.q(_w_3621));
  inv inv_G153(.a(G153_1),.q(G5207));
  bfr _b_4879(.a(_w_6304),.q(_w_6305));
  and_bi g769(.a(n767),.b(n768),.q(n769));
  bfr _b_4845(.a(_w_6270),.q(n1270));
  bfr _b_5374(.a(_w_6799),.q(_w_6800));
  spl4L G124_s_0(.a(G124),.q0(G124_0),.q1(G124_1),.q2(G124_2),.q3(G124_3));
  or_bb g1407(.a(n1402),.b(n1406),.q(_w_5893));
  bfr _b_6023(.a(_w_7448),.q(_w_7447));
  bfr _b_5791(.a(_w_7216),.q(_w_7217));
  bfr _b_2729(.a(_w_4154),.q(_w_4155));
  bfr _b_1952(.a(_w_3377),.q(_w_3378));
  or_bb g775(.a(n463_1),.b(n773_1),.q(n775));
  bfr _b_2168(.a(_w_3593),.q(_w_3594));
  and_bi g326(.a(n325),.b(G141_1),.q(n326));
  bfr _b_2757(.a(_w_4182),.q(_w_4183));
  inv inv_G99(.a(G99_1),.q(G5206));
  or_bb g573(.a(G2_1),.b(n381_2),.q(_w_6065));
  and_bi g779(.a(n778),.b(n777),.q(n779));
  bfr _b_3589(.a(_w_5014),.q(_w_5015));
  and_bi g830(.a(G172_7),.b(n829),.q(n830));
  bfr _b_2783(.a(_w_4208),.q(_w_4209));
  bfr _b_4083(.a(_w_5508),.q(_w_5509));
  and_bb g782(.a(n466_1),.b(n773_2),.q(n782));
  bfr _b_7477(.a(_w_8902),.q(_w_8903));
  spl2 g419_s_0(.a(n419),.q0(n419_0),.q1(_w_3814));
  and_bi g252(.a(G130_1),.b(G101_7),.q(n252));
  or_bb g783(.a(n781),.b(n782),.q(n783));
  spl4L G128_s_0(.a(G128),.q0(G128_0),.q1(G128_1),.q2(G128_2),.q3(_w_5896));
  bfr _b_5227(.a(_w_6652),.q(_w_6653));
  and_bb g785(.a(n472_7),.b(n783_1),.q(n785));
  or_bb g965(.a(G170_3),.b(n246_1),.q(n965));
  bfr _b_2247(.a(_w_3672),.q(G158_0));
  spl4L g403_s_0(.a(n403),.q0(_w_4073),.q1(n403_1),.q2(_w_4074),.q3(_w_4076));
  and_bb g1206(.a(n1184_1),.b(n1204_1),.q(n1206));
  bfr _b_4401(.a(_w_5826),.q(n1251));
  bfr _b_4728(.a(_w_6153),.q(_w_6154));
  and_bi g786(.a(n784),.b(n785),.q(n786));
  and_bb g1322(.a(n1314_1),.b(n1320_1),.q(n1322));
  and_bi g845(.a(G173_4),.b(G5249_1),.q(n845));
  or_bb g788(.a(n465_2),.b(n773_5),.q(n788));
  or_bb g1245(.a(n1235_0),.b(n1244_0),.q(n1245));
  and_bb g1452(.a(G4_0),.b(n586_11),.q(n1452));
  bfr _b_5922(.a(_w_7347),.q(_w_7348));
  and_bi g1349(.a(n1348),.b(G143_6),.q(n1349));
  bfr _b_2475(.a(_w_3900),.q(_w_3901));
  spl4L G124_s_2(.a(G124_1),.q0(G124_8),.q1(G124_9),.q2(G124_10),.q3(G124_11));
  bfr _b_3440(.a(_w_4865),.q(_w_4866));
  bfr _b_5759(.a(G20),.q(_w_7185));
  bfr _b_4050(.a(_w_5475),.q(_w_5476));
  and_bi g981(.a(G176_8),.b(n249_1),.q(n981));
  and_bi g1182(.a(n1181),.b(n1180),.q(_w_5897));
  bfr _b_2710(.a(_w_4135),.q(_w_4136));
  spl2 G115_s_1(.a(G115_3),.q0(G115_4),.q1(G115_5));
  bfr _b_6096(.a(_w_7521),.q(_w_7522));
  and_bi g204(.a(n203),.b(n201),.q(_w_5297));
  and_bb g790(.a(G5251_1),.b(n556_1),.q(n790));
  bfr _b_6650(.a(_w_8075),.q(_w_8076));
  and_bi g1406(.a(n1405),.b(G141_6),.q(n1406));
  bfr _b_5061(.a(_w_6486),.q(_w_6484));
  spl2 G124_s_5(.a(G124_18),.q0(G124_20),.q1(G124_21));
  and_bb g792(.a(n620_1),.b(n791),.q(n792));
  bfr _b_5841(.a(_w_7266),.q(_w_7267));
  and_bi g324(.a(G166_11),.b(G96_6),.q(n324));
  and_bb g794(.a(n600_1),.b(n793),.q(_w_5899));
  bfr _b_5776(.a(_w_7201),.q(_w_7202));
  and_bb g910(.a(G64_21),.b(n909),.q(G5277));
  bfr _b_7182(.a(_w_8607),.q(_w_8608));
  bfr _b_6822(.a(_w_8247),.q(_w_8248));
  bfr _b_3479(.a(_w_4904),.q(_w_4905));
  bfr _b_6771(.a(_w_8196),.q(_w_8197));
  bfr _b_2084(.a(_w_3509),.q(G171_0));
  and_bi g796(.a(n795),.b(n786_0),.q(n796));
  bfr _b_7489(.a(_w_8914),.q(_w_8915));
  and_bi g968(.a(n967),.b(n963),.q(_w_6126));
  and_bi g1025(.a(G177_9),.b(n1024),.q(n1025));
  bfr _b_3852(.a(_w_5277),.q(_w_5278));
  spl4L G173_s_0(.a(_w_7004),.q0(_w_5903),.q1(_w_5905),.q2(_w_5907),.q3(G173_3));
  bfr _b_7479(.a(_w_8904),.q(_w_8905));
  bfr _b_6142(.a(_w_7567),.q(_w_7568));
  and_bb g259(.a(n243_0),.b(n258),.q(n259));
  or_bb g798(.a(G158_15),.b(G5250_4),.q(n798));
  spl4L G148_s_0(.a(_w_6562),.q0(G148_0),.q1(G148_1),.q2(_w_5663),.q3(G148_3));
  bfr _b_2096(.a(_w_3521),.q(G121_9));
  and_bi g799(.a(G158_27),.b(G5248_4),.q(n799));
  bfr _b_2104(.a(_w_3529),.q(_w_3530));
  and_bb g801(.a(n798),.b(n800),.q(_w_5921));
  or_bb g677(.a(n387_2),.b(n665_1),.q(_w_5707));
  or_bb g828(.a(G173_22),.b(G5258_1),.q(_w_5922));
  bfr _b_5245(.a(_w_6670),.q(_w_6671));
  bfr _b_2340(.a(_w_3765),.q(_w_3766));
  and_bi g803(.a(G81_0),.b(n802_0),.q(n803));
  bfr _b_5000(.a(G120),.q(_w_6426));
  and_bi g804(.a(G158_25),.b(G159_5),.q(n804));
  or_bb g483(.a(G113_4),.b(G115_4),.q(n483));
  spl4L G2_s_0(.a(_w_7175),.q0(G2_0),.q1(G2_1),.q2(_w_3888),.q3(_w_3894));
  bfr _b_3700(.a(_w_5125),.q(_w_5126));
  spl2 g637_s_0(.a(n637),.q0(_w_5945),.q1(n637_1));
  bfr _b_2717(.a(_w_4142),.q(n414_2));
  or_bb g807(.a(n801),.b(n806),.q(_w_5947));
  bfr _b_5555(.a(_w_6980),.q(_w_6981));
  and_bi g228(.a(G146_0),.b(n227),.q(n228));
  bfr _b_2650(.a(_w_4075),.q(n403_2));
  and_bi g199(.a(n198),.b(n196),.q(_w_5949));
  bfr _b_4813(.a(_w_6238),.q(_w_6239));
  spl2 G23_s_0(.a(_w_7244),.q0(G23_0),.q1(G23_1));
  and_bi g822(.a(G172_6),.b(n821),.q(n822));
  or_bb g1384(.a(n1382),.b(n1383),.q(n1384));
  bfr _b_4755(.a(_w_6180),.q(n227));
  and_bb g202(.a(_w_6391),.b(G163_10),.q(_w_5981));
  and_bi g832(.a(G6_0),.b(n588_4),.q(n832));
  bfr _b_4618(.a(_w_6043),.q(_w_6044));
  and_bb g787(.a(n465_1),.b(n773_4),.q(n787));
  bfr _b_2157(.a(_w_3582),.q(_w_3583));
  bfr _b_6209(.a(_w_7634),.q(_w_7635));
  bfr _b_5667(.a(_w_7092),.q(_w_7093));
  bfr _b_2532(.a(_w_3957),.q(G5213));
  spl4L G124_s_1(.a(G124_0),.q0(G124_4),.q1(G124_5),.q2(G124_6),.q3(G124_7));
  bfr _b_4978(.a(G110),.q(_w_6404));
  bfr _b_5735(.a(_w_7160),.q(_w_7161));
  or_bb g826(.a(n824),.b(n825),.q(n826));
  bfr _b_6185(.a(_w_7610),.q(_w_7611));
  bfr _b_2259(.a(_w_3684),.q(_w_3685));
  and_bb g833(.a(G27_0),.b(n586_4),.q(n833));
  bfr _b_5594(.a(_w_7019),.q(_w_7020));
  or_bb g836(.a(G173_20),.b(G5259_1),.q(n836));
  and_bb g1391(.a(G102_15),.b(G105_12),.q(n1391));
  bfr _b_3239(.a(_w_4664),.q(_w_4665));
  spl2 g719_s_0(.a(n719),.q0(n719_0),.q1(n719_1));
  bfr _b_6757(.a(_w_8182),.q(_w_8183));
  bfr _b_3380(.a(_w_4805),.q(_w_4806));
  and_bb g593(.a(n443_2),.b(n450_1),.q(n593));
  bfr _b_6208(.a(_w_7633),.q(_w_7634));
  and_bb g831(.a(n828),.b(n830),.q(_w_5982));
  bfr _b_2401(.a(_w_3826),.q(_w_3827));
  bfr _b_4414(.a(_w_5839),.q(_w_5840));
  bfr _b_5787(.a(G22),.q(_w_7213));
  bfr _b_4866(.a(_w_6291),.q(n229));
  bfr _b_5238(.a(_w_6663),.q(_w_6664));
  spl2 g725_s_0(.a(n725),.q0(n725_0),.q1(n725_1));
  and_bb g839(.a(n836),.b(n838),.q(_w_5983));
  and_bi g841(.a(G5_0),.b(n588_5),.q(n841));
  bfr _b_5367(.a(_w_6792),.q(_w_6793));
  bfr _b_5193(.a(_w_6618),.q(_w_6619));
  bfr _b_5150(.a(_w_6575),.q(_w_6576));
  or_bb g842(.a(n840),.b(n841),.q(n842));
  or_bb g843(.a(n839),.b(n842),.q(_w_5984));
  bfr _b_2240(.a(_w_3665),.q(G158_22));
  bfr _b_7309(.a(_w_8734),.q(_w_8735));
  or_bb g844(.a(G173_16),.b(G5260_1),.q(n844));
  and_bb g1266(.a(n381_4),.b(n386_4),.q(_w_5987));
  and_bb g847(.a(n844),.b(n846),.q(_w_5990));
  spl4L G94_s_3(.a(G94_3),.q0(G94_10),.q1(G94_11),.q2(G94_12),.q3(G94_13));
  or_bi g972(.a(n970),.b(n971),.q(_w_5991));
  and_bb g622(.a(G176_46),.b(n277_1),.q(n622));
  and_bi g1253(.a(n249_2),.b(n246_3),.q(_w_6011));
  spl2 G75_s_0(.a(_w_8502),.q0(G75_0),.q1(G75_1));
  and_bb g422(.a(G124_8),.b(G94_7),.q(n422));
  bfr _b_6403(.a(_w_7828),.q(_w_7829));
  and_bi g1419(.a(n1417),.b(n1418),.q(n1419));
  and_bi g849(.a(G25_0),.b(n588_6),.q(n849));
  bfr _b_4780(.a(_w_6205),.q(_w_6206));
  spl2 g666_s_0(.a(n666),.q0(n666_0),.q1(n666_1));
  and_bi g757(.a(n756),.b(n752_0),.q(_w_4821));
  bfr _b_4288(.a(_w_5713),.q(_w_5714));
  and_bi g1210(.a(G148_6),.b(G100_16),.q(n1210));
  or_bb g1201(.a(n1199),.b(n1200),.q(n1201));
  and_bb g857(.a(G16_1),.b(n630_1),.q(n857));
  bfr _b_2153(.a(_w_3578),.q(_w_3579));
  bfr _b_7553(.a(_w_8978),.q(_w_8979));
  and_bb g1188(.a(G162_0),.b(n442_7),.q(n1188));
  and_bi g1129(.a(G160_13),.b(G5288_5),.q(n1129));
  and_bi g441(.a(G131_0),.b(G123_20),.q(n441));
  bfr _b_6907(.a(G70),.q(_w_8333));
  bfr _b_6314(.a(_w_7739),.q(_w_7740));
  or_bb g860(.a(G174_22),.b(G5258_2),.q(_w_6020));
  bfr _b_6300(.a(_w_7725),.q(_w_7726));
  bfr _b_4237(.a(_w_5662),.q(G5229_0));
  bfr _b_5345(.a(_w_6770),.q(_w_6771));
  and_bb g1440(.a(n1341),.b(n1439),.q(n1440));
  and_bi g912(.a(G158_4),.b(G5254_4),.q(n912));
  spl2 g1407_s_0(.a(n1407),.q0(n1407_0),.q1(n1407_1));
  bfr _b_4378(.a(_w_5803),.q(_w_5804));
  bfr _b_2253(.a(_w_3678),.q(_w_3679));
  or_bb g1275(.a(n1273),.b(n1274),.q(n1275));
  and_bi g657(.a(n400_4),.b(n655_1),.q(n657));
  or_bb g866(.a(n864),.b(n865),.q(n866));
  bfr _b_2125(.a(_w_3550),.q(_w_3551));
  or_bb g408(.a(G142_3),.b(n406_1),.q(n408));
  or_bb g868(.a(G174_20),.b(G5259_2),.q(n868));
  bfr _b_5709(.a(_w_7134),.q(_w_7135));
  bfr _b_3729(.a(_w_5154),.q(n918));
  and_bi g869(.a(G174_17),.b(G5255_2),.q(n869));
  bfr _b_6439(.a(_w_7864),.q(_w_7865));
  and_bi g872(.a(G5_1),.b(n632_5),.q(n872));
  bfr _b_4763(.a(_w_6188),.q(G115_0));
  and_bi g600(.a(n598),.b(n599),.q(n600));
  bfr _b_2914(.a(_w_4339),.q(G159_3));
  and_bi g878(.a(G175_9),.b(n877),.q(n878));
  and_bb g879(.a(n876),.b(n878),.q(_w_6032));
  and_bi g1142(.a(G75_1),.b(n813_8),.q(n1142));
  spl2 G131_s_0(.a(_w_6438),.q0(G131_0),.q1(_w_3524));
  bfr _b_3667(.a(_w_5092),.q(_w_5093));
  and_bi g671(.a(n670_0),.b(G176_51),.q(n671));
  bfr _b_4574(.a(_w_5999),.q(_w_6000));
  bfr _b_2020(.a(_w_3445),.q(_w_3446));
  and_bb g955(.a(G64_4),.b(n954),.q(G5282));
  bfr _b_4169(.a(_w_5594),.q(n982));
  bfr _b_5609(.a(_w_7034),.q(_w_7035));
  and_bb g880(.a(G24_1),.b(n630_6),.q(n880));
  and_bi g1070(.a(G175_11),.b(n1069),.q(n1070));
  bfr _b_5044(.a(_w_6469),.q(_w_6470));
  or_bb g884(.a(G158_24),.b(G5257_4),.q(n884));
  and_bi g885(.a(G158_23),.b(G5253_4),.q(n885));
  bfr _b_2996(.a(_w_4421),.q(_w_4422));
  bfr _b_4057(.a(_w_5482),.q(_w_5483));
  spl2 g556_s_0(.a(n556),.q0(_w_6041),.q1(n556_1));
  bfr _b_2403(.a(_w_3828),.q(_w_3829));
  bfr _b_3387(.a(_w_4812),.q(_w_4813));
  and_bi g886(.a(G159_6),.b(n885),.q(n886));
  and_bi g648(.a(G177_23),.b(n647),.q(_w_6042));
  bfr _b_3865(.a(_w_5290),.q(_w_5291));
  bfr _b_4100(.a(_w_5525),.q(_w_5526));
  bfr _b_6716(.a(_w_8141),.q(_w_8142));
  and_bi g861(.a(G174_21),.b(G5254_2),.q(n861));
  and_bi g304(.a(G166_9),.b(G92_6),.q(n304));
  bfr _b_5444(.a(_w_6869),.q(_w_6870));
  or_bb g1170(.a(n1165),.b(n1169),.q(n1170));
  or_bb g891(.a(n887),.b(n890),.q(_w_6045));
  and_bi g895(.a(G159_7),.b(n894),.q(n895));
  bfr _b_5206(.a(_w_6631),.q(_w_6632));
  and_bi g1465(.a(G159_14),.b(n1464),.q(_w_6047));
  bfr _b_7478(.a(_w_8903),.q(_w_8904));
  bfr _b_5874(.a(_w_7299),.q(_w_7300));
  bfr _b_3054(.a(_w_4479),.q(_w_4480));
  and_bi g897(.a(G72_0),.b(n802_4),.q(n897));
  bfr _b_7257(.a(_w_8682),.q(_w_8683));
  and_bb g505(.a(n491_1),.b(n503_1),.q(n505));
  bfr _b_3849(.a(_w_5274),.q(_w_5275));
  and_bi g846(.a(G172_9),.b(n845),.q(n846));
  bfr _b_5764(.a(_w_7189),.q(_w_7190));
  and_bi g838(.a(G172_8),.b(n837),.q(n838));
  bfr _b_3074(.a(_w_4499),.q(_w_4500));
  or_bb g899(.a(n897),.b(n898),.q(n899));
  bfr _b_7440(.a(_w_8865),.q(_w_8866));
  bfr _b_5533(.a(_w_6958),.q(_w_6959));
  bfr _b_5133(.a(_w_6558),.q(_w_6550));
  bfr _b_2176(.a(_w_3601),.q(_w_3602));
  and_bb g721(.a(n716_1),.b(n719_1),.q(n721));
  or_bb g1137(.a(G160_12),.b(G5292_5),.q(_w_6050));
  bfr _b_3767(.a(_w_5192),.q(_w_5193));
  bfr _b_6109(.a(_w_7534),.q(_w_7535));
  spl4L G146_s_0(.a(_w_6550),.q0(G146_0),.q1(G146_1),.q2(_w_6024),.q3(_w_6026));
  and_bb g901(.a(G64_22),.b(n900),.q(G5276));
  bfr _b_6225(.a(_w_7650),.q(_w_7651));
  bfr _b_4573(.a(_w_5998),.q(_w_5999));
  bfr _b_4252(.a(_w_5677),.q(_w_5678));
  and_bi g904(.a(G159_8),.b(n903),.q(n904));
  and_bb g1154(.a(G64_8),.b(n1153),.q(_w_6051));
  and_bi g732(.a(n406_2),.b(n372_2),.q(n732));
  or_bb g908(.a(n906),.b(n907),.q(n908));
  and_bi g913(.a(G159_9),.b(n912),.q(n913));
  and_bb g466(.a(n459_0),.b(n465_0),.q(n466));
  and_bi g915(.a(G68_0),.b(n802_6),.q(n915));
  bfr _b_5633(.a(_w_7058),.q(_w_7059));
  spl4L G177_s_6(.a(G177_18),.q0(G177_22),.q1(G177_23),.q2(G177_24),.q3(G177_25));
  bfr _b_3091(.a(_w_4516),.q(_w_4517));
  bfr _b_4700(.a(_w_6125),.q(n456_6));
  and_bb g916(.a(G69_0),.b(n804_6),.q(n916));
  or_bb g665(.a(n379_2),.b(n572_1),.q(n665));
  spl3L g457_s_0(.a(n457),.q0(n457_0),.q1(_w_3490),.q2(n457_2));
  bfr _b_2626(.a(_w_4051),.q(_w_4052));
  bfr _b_7143(.a(_w_8568),.q(_w_8536));
  spl4L g391_s_0(.a(n391),.q0(n391_0),.q1(n391_1),.q2(n391_2),.q3(n391_3));
  and_bb g264(.a(G121_5),.b(G167_4),.q(n264));
  bfr _b_3285(.a(_w_4710),.q(_w_4711));
  bfr _b_4223(.a(_w_5648),.q(_w_5649));
  bfr _b_7498(.a(_w_8923),.q(_w_8924));
  and_bi g921(.a(G160_23),.b(G5253_5),.q(n921));
  and_bi g1262(.a(G177_8),.b(n1261),.q(_w_4694));
  bfr _b_4261(.a(_w_5686),.q(n541));
  and_bi g1078(.a(G175_12),.b(n1077),.q(n1078));
  bfr _b_7228(.a(_w_8653),.q(_w_8654));
  spl2 g1272_s_0(.a(n1272),.q0(n1272_0),.q1(n1272_1));
  and_bi g924(.a(G76_1),.b(n813_1),.q(n924));
  and_bb g934(.a(G82_1),.b(n815_4),.q(n934));
  and_bb g1171(.a(n1170_0),.b(n686_2),.q(n1171));
  spl4L G177_s_7(.a(G177_19),.q0(G177_26),.q1(G177_27),.q2(G177_28),.q3(G177_29));
  or_bb g1255(.a(n1252_0),.b(n1254_0),.q(n1255));
  or_bb g927(.a(n923),.b(n926),.q(_w_6066));
  bfr _b_3765(.a(_w_5190),.q(_w_5191));
  and_bb g234(.a(n224_0),.b(n233_0),.q(n234));
  bfr _b_4531(.a(_w_5956),.q(_w_5957));
  bfr _b_4795(.a(_w_6220),.q(_w_6221));
  and_bi g931(.a(G161_7),.b(n930),.q(n931));
  or_bb g917(.a(n915),.b(n916),.q(n917));
  bfr _b_7316(.a(_w_8741),.q(_w_8742));
  and_bi g1228(.a(G128_11),.b(G101_10),.q(n1228));
  and_bb g764(.a(n426_1),.b(n744_5),.q(n764));
  or_bb g935(.a(n933),.b(n934),.q(n935));
  bfr _b_4255(.a(_w_5680),.q(_w_5681));
  bfr _b_4723(.a(_w_6148),.q(n988));
  bfr _b_2091(.a(_w_3516),.q(_w_3517));
  bfr _b_3451(.a(_w_4876),.q(_w_4877));
  or_bb g1144(.a(n1140),.b(n1143),.q(n1144));
  bfr _b_2191(.a(_w_3616),.q(_w_3617));
  bfr _b_3482(.a(_w_4907),.q(_w_4908));
  and_bi g1344(.a(n1342),.b(n1343),.q(n1344));
  and_bb g937(.a(G64_16),.b(n936),.q(_w_6099));
  bfr _b_4331(.a(_w_5756),.q(_w_5757));
  spl2 g655_s_0(.a(n655),.q0(n655_0),.q1(n655_1));
  bfr _b_2354(.a(_w_3779),.q(_w_3780));
  bfr _b_5954(.a(_w_7379),.q(_w_7380));
  spl4L g448_s_0(.a(n448),.q0(n448_0),.q1(n448_1),.q2(n448_2),.q3(n448_3));
  bfr _b_2444(.a(_w_3869),.q(_w_3870));
  bfr _b_4858(.a(_w_6283),.q(n256));
  bfr _b_4303(.a(_w_5728),.q(_w_5729));
  and_bb g1466(.a(n1463),.b(n1465),.q(n1466));
  bfr _b_4920(.a(_w_6345),.q(_w_6346));
  bfr _b_2283(.a(_w_3708),.q(_w_3709));
  bfr _b_3043(.a(_w_4468),.q(_w_4469));
  or_bb g945(.a(n941),.b(n944),.q(n945));
  bfr _b_7112(.a(_w_8537),.q(_w_8538));
  and_bb g946(.a(G64_15),.b(n945),.q(_w_6113));
  and_bi g789(.a(n788),.b(n787),.q(n789));
  and_bi g949(.a(G161_9),.b(n948),.q(n949));
  bfr _b_7025(.a(_w_8450),.q(_w_8451));
  bfr _b_2033(.a(_w_3458),.q(_w_3459));
  bfr _b_5852(.a(G24),.q(_w_7278));
  or_bb g1227(.a(G100_14),.b(G128_10),.q(n1227));
  and_bb g285(.a(G167_6),.b(G94_5),.q(n285));
  and_bb g816(.a(G80_1),.b(n815_0),.q(n816));
  spl4L g813_s_0(.a(n813),.q0(n813_0),.q1(n813_1),.q2(n813_2),.q3(n813_3));
  bfr _b_2642(.a(_w_4067),.q(_w_4068));
  spl4L g1009_s_0(.a(G5290_0),.q0(_w_6116),.q1(G5290_1),.q2(G5290_2),.q3(G5290_3));
  bfr _b_3318(.a(_w_4743),.q(n196));
  bfr _b_6811(.a(_w_8236),.q(_w_8237));
  bfr _b_3874(.a(_w_5299),.q(_w_5300));
  or_bb g1235(.a(n1230),.b(n1234),.q(n1235));
  or_bb g953(.a(n951),.b(n952),.q(n953));
  bfr _b_7282(.a(_w_8707),.q(_w_8708));
  bfr _b_2515(.a(_w_3940),.q(_w_3941));
  bfr _b_7418(.a(_w_8843),.q(_w_8844));
  or_bb g817(.a(n814),.b(n816),.q(n817));
  spl2 g1440_s_0(.a(n1440),.q0(n1440_0),.q1(n1440_1));
  bfr _b_5156(.a(_w_6581),.q(_w_6582));
  and_bi g958(.a(G61_1),.b(n469_8),.q(n958));
  or_bb g959(.a(n957),.b(n958),.q(n959));
  bfr _b_1987(.a(_w_3412),.q(_w_3413));
  bfr _b_5654(.a(_w_7079),.q(_w_7080));
  bfr _b_2249(.a(_w_3674),.q(G158_1));
  bfr _b_6369(.a(_w_7794),.q(_w_7795));
  spl2 g401_s_0(.a(n401),.q0(n401_0),.q1(n401_1));
  spl3L g456_s_1(.a(n456_3),.q0(n456_4),.q1(n456_5),.q2(_w_6124));
  or_bb g1408(.a(G100_6),.b(G109_10),.q(n1408));
  and_bi g966(.a(n965),.b(n964),.q(n966));
  spl4L g424_s_0(.a(n424),.q0(n424_0),.q1(n424_1),.q2(n424_2),.q3(n424_3));
  bfr _b_4276(.a(_w_5701),.q(G5302));
  and_bi g555(.a(G21_1),.b(n442_2),.q(n555));
  or_bb g967(.a(G171_1),.b(n966),.q(n967));
  bfr _b_2643(.a(_w_4068),.q(_w_4069));
  bfr _b_6236(.a(G42),.q(_w_7662));
  bfr _b_3517(.a(_w_4942),.q(n356));
  spl4L G169_s_0(.a(G169),.q0(G169_0),.q1(G169_1),.q2(G169_2),.q3(G169_3));
  and_bi g975(.a(G176_6),.b(n246_2),.q(n975));
  bfr _b_5020(.a(_w_6445),.q(_w_6446));
  spl4L G88_s_1(.a(G88_3),.q0(_w_5881),.q1(G88_5),.q2(G88_6),.q3(G88_7));
  bfr _b_2562(.a(_w_3987),.q(_w_3988));
  bfr _b_4908(.a(_w_6333),.q(_w_6334));
  and_bb g987(.a(G176_10),.b(n224_1),.q(n987));
  or_bb g992(.a(G176_20),.b(n789_1),.q(n992));
  and_bi g518(.a(n516),.b(n517),.q(n518));
  bfr _b_2094(.a(_w_3519),.q(_w_3520));
  and_bb g999(.a(G5199_1),.b(n998),.q(n999));
  and_bi g1000(.a(n999),.b(G5242_1),.q(n1000));
  spl4L g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1),.q2(_w_6134),.q3(_w_6138));
  or_bb g1128(.a(G160_14),.b(G5293_5),.q(_w_6139));
  and_bi g1002(.a(n1001),.b(G5261_1),.q(n1002));
  bfr _b_4313(.a(_w_5738),.q(n409_2));
  spl2 g356_s_0(.a(n356),.q0(n356_0),.q1(_w_6140));
  and_bi g1005(.a(n749_1),.b(G176_22),.q(n1005));
  and_bi g988(.a(G177_14),.b(n987),.q(_w_6141));
  or_bb g556(.a(n554),.b(n555),.q(_w_6151));
  bfr _b_3626(.a(_w_5051),.q(n575));
  and_bb g1010(.a(_w_7736),.b(n552_9),.q(_w_6157));
  bfr _b_5725(.a(_w_7150),.q(_w_7151));
  spl2 g1170_s_0(.a(n1170),.q0(n1170_0),.q1(n1170_1));
  bfr _b_3113(.a(_w_4538),.q(_w_4539));
  and_bi g624(.a(n623),.b(n621),.q(_w_6164));
  bfr _b_2378(.a(_w_3803),.q(n375_4));
  bfr _b_3441(.a(_w_4866),.q(_w_4867));
  and_bb g991(.a(_w_7694),.b(n552_11),.q(_w_6129));
  and_bi g1011(.a(n763_1),.b(G176_4),.q(n1011));
  and_bi g691(.a(n686_1),.b(n689_1),.q(n691));
  bfr _b_4156(.a(_w_5581),.q(_w_5582));
  bfr _b_6281(.a(_w_7706),.q(_w_7707));
  bfr _b_4864(.a(_w_6289),.q(n1113));
  and_bi g490(.a(n485_1),.b(n488_1),.q(n490));
  bfr _b_2790(.a(_w_4215),.q(_w_4216));
  and_bb g1012(.a(G176_25),.b(n298_1),.q(_w_6168));
  bfr _b_6424(.a(_w_7849),.q(_w_7850));
  spl4L G130_s_0(.a(G130),.q0(_w_5248),.q1(_w_5250),.q2(_w_5252),.q3(G130_3));
  bfr _b_4424(.a(_w_5849),.q(_w_5850));
  and_bi g1013(.a(G177_11),.b(n1012),.q(_w_6173));
  bfr _b_5083(.a(_w_6508),.q(_w_6509));
  and_bi g1237(.a(G126_11),.b(G101_11),.q(n1237));
  and_bb g1124(.a(G83_0),.b(n804_10),.q(n1124));
  bfr _b_4671(.a(_w_6096),.q(_w_6097));
  and_bi g701(.a(n699),.b(n700),.q(n701));
  and_bb g923(.a(n920),.b(n922),.q(n923));
  bfr _b_2827(.a(_w_4252),.q(n547_1));
  and_bi g227(.a(n225),.b(n226),.q(_w_6177));
  bfr _b_5412(.a(_w_6837),.q(_w_6838));
  or_bb g1028(.a(G174_14),.b(G5290_1),.q(_w_6189));
  spl2 g565_s_0(.a(n565),.q0(n565_0),.q1(n565_1));
  bfr _b_2941(.a(_w_4366),.q(G5299));
  and_ii g1021(.a(n1016),.b(n1020),.q(_w_6190));
  bfr _b_3889(.a(_w_5314),.q(_w_5315));
  and_ii g1442(.a(n1440_0),.b(n1441),.q(_w_6191));
  bfr _b_4015(.a(_w_5440),.q(_w_5441));
  or_bb g875(.a(n871),.b(n874),.q(_w_6196));
  bfr _b_6984(.a(_w_8409),.q(_w_8410));
  spl4L g615_s_0(.a(G5254_0),.q0(_w_4010),.q1(G5254_1),.q2(G5254_2),.q3(G5254_3));
  and_bb g314(.a(G109_5),.b(G167_9),.q(n314));
  bfr _b_4067(.a(_w_5492),.q(n1007));
  bfr _b_4380(.a(_w_5805),.q(_w_5806));
  and_bb g1024(.a(G176_29),.b(n289_1),.q(n1024));
  and_bb g1026(.a(n1023),.b(n1025),.q(n1026));
  bfr _b_1985(.a(_w_3410),.q(_w_3411));
  bfr _b_5950(.a(_w_7375),.q(_w_7343));
  or_bb g464(.a(G146_3),.b(n462_1),.q(n464));
  spl2 G61_s_0(.a(_w_8134),.q0(G61_0),.q1(G61_1));
  bfr _b_3369(.a(_w_4794),.q(_w_4795));
  and_bb g546(.a(n414_1),.b(n545_0),.q(n546));
  and_bi g1030(.a(G175_10),.b(n1029),.q(n1030));
  bfr _b_4756(.a(_w_6181),.q(_w_6182));
  bfr _b_2549(.a(_w_3974),.q(_w_3975));
  and_bb g1031(.a(n1028),.b(n1030),.q(_w_6207));
  and_bb g1033(.a(G42_0),.b(n630_7),.q(n1033));
  bfr _b_3335(.a(_w_4760),.q(n307));
  spl2 g760_s_0(.a(n760),.q0(n760_0),.q1(n760_1));
  and_bb g1280(.a(n380_1),.b(n385_2),.q(_w_6353));
  or_bb g1036(.a(G173_14),.b(G5290_2),.q(_w_6211));
  bfr _b_4686(.a(_w_6111),.q(_w_6112));
  and_bi g1037(.a(G173_13),.b(G5285_2),.q(n1037));
  or_bb g1414(.a(n1412),.b(n1413),.q(n1414));
  or_bb g1045(.a(G173_11),.b(G5291_1),.q(n1045));
  bfr _b_4396(.a(_w_5821),.q(_w_5822));
  spl3L g597_s_0(.a(n597),.q0(n597_0),.q1(n597_1),.q2(n597_2));
  bfr _b_4810(.a(_w_6235),.q(n1293));
  and_bb g1048(.a(G17_0),.b(n586_8),.q(n1048));
  bfr _b_2116(.a(_w_3541),.q(_w_3542));
  bfr _b_4600(.a(_w_6025),.q(G146_2));
  or_bb g1190(.a(G162_1),.b(n439_3),.q(n1190));
  bfr _b_3843(.a(_w_5268),.q(_w_5269));
  bfr _b_5382(.a(_w_6807),.q(_w_6808));
  or_bb g1050(.a(n1048),.b(n1049),.q(n1050));
  spl4L g400_s_0(.a(n400),.q0(n400_0),.q1(_w_6212),.q2(_w_6215),.q3(n400_3));
  and_bb g1062(.a(G172_13),.b(n1061),.q(n1062));
  spl4L G98_s_2(.a(G98_1),.q0(G98_8),.q1(G98_9),.q2(G98_10),.q3(G98_11));
  bfr _b_2075(.a(_w_3500),.q(_w_3501));
  and_bi g951(.a(G68_1),.b(n813_6),.q(n951));
  or_bb g1313(.a(n413_3),.b(n545_3),.q(_w_6222));
  and_bb g652(.a(n388_1),.b(n394_1),.q(n652));
  bfr _b_2628(.a(_w_4053),.q(_w_4054));
  bfr _b_3484(.a(_w_4909),.q(_w_4910));
  bfr _b_4881(.a(_w_6306),.q(n1158));
  bfr _b_3878(.a(_w_5303),.q(_w_5304));
  bfr _b_5920(.a(_w_7345),.q(_w_7346));
  bfr _b_4754(.a(_w_6179),.q(_w_6180));
  or_bb g784(.a(n472_6),.b(n783_0),.q(n784));
  and_bi g1052(.a(G173_10),.b(G5287_1),.q(_w_6226));
  and_bb g1468(.a(G78_0),.b(n804_11),.q(n1468));
  or_bb g1053(.a(G173_9),.b(G5292_1),.q(n1053));
  spl2 g605_s_1(.a(G5253_3),.q0(G5253_4),.q1(G5253_5));
  or_bb g1294(.a(n1285_1),.b(n1292_1),.q(n1294));
  bfr _b_2720(.a(_w_4145),.q(_w_4146));
  bfr _b_4407(.a(_w_5832),.q(_w_5833));
  or_bb g1061(.a(G173_7),.b(G5293_1),.q(n1061));
  bfr _b_2844(.a(_w_4269),.q(n429_1));
  bfr _b_4256(.a(_w_5681),.q(n413_3));
  bfr _b_6682(.a(_w_8107),.q(_w_8108));
  bfr _b_4949(.a(_w_6374),.q(_w_6375));
  and_bi g1165(.a(n463_4),.b(n1164_0),.q(_w_6229));
  bfr _b_3050(.a(_w_4475),.q(_w_4476));
  bfr _b_5455(.a(_w_6880),.q(_w_6881));
  bfr _b_2376(.a(_w_3801),.q(G5293));
  and_bb g1064(.a(G36_0),.b(n586_10),.q(n1064));
  bfr _b_5336(.a(_w_6761),.q(_w_6762));
  bfr _b_1959(.a(_w_3384),.q(_w_3385));
  spl4L g744_s_0(.a(n744),.q0(n744_0),.q1(n744_1),.q2(n744_2),.q3(n744_3));
  bfr _b_5082(.a(_w_6507),.q(_w_6508));
  and_bi g1065(.a(G15_0),.b(n588_10),.q(n1065));
  or_bb g1066(.a(n1064),.b(n1065),.q(n1066));
  bfr _b_4185(.a(_w_5610),.q(_w_5611));
  spl4L G174_s_6(.a(G174_19),.q0(_w_3733),.q1(G174_25),.q2(G174_26),.q3(G174_27));
  and_bb g1293(.a(n1285_0),.b(n1292_0),.q(_w_6235));
  bfr _b_6939(.a(_w_8364),.q(_w_8365));
  bfr _b_2330(.a(_w_3755),.q(_w_3756));
  or_ii g184(.a(G136),.b(G154),.q(_w_6236));
  bfr _b_5424(.a(_w_6849),.q(_w_6850));
  spl4L g813_s_2(.a(n813_3),.q0(n813_8),.q1(n813_9),.q2(n813_10),.q3(n813_11));
  bfr _b_4369(.a(_w_5794),.q(_w_5795));
  spl4L G101_s_3(.a(G101_2),.q0(G101_12),.q1(G101_13),.q2(G101_14),.q3(G101_15));
  bfr _b_3527(.a(_w_4952),.q(G5253_0));
  bfr _b_6221(.a(_w_7646),.q(_w_7647));
  and_bi g1270(.a(n1269),.b(n534_1),.q(_w_6268));
  bfr _b_5956(.a(_w_7381),.q(_w_7382));
  bfr _b_5844(.a(_w_7269),.q(_w_7270));
  bfr _b_5138(.a(G149),.q(_w_6564));
  bfr _b_2177(.a(_w_3602),.q(_w_3603));
  and_bb g407(.a(G142_2),.b(n406_0),.q(n407));
  bfr _b_4159(.a(_w_5584),.q(n491));
  and_bi g1429(.a(n1407_0),.b(n1428_0),.q(n1429));
  or_bb g1082(.a(n1080),.b(n1081),.q(n1082));
  and_bi g1168(.a(n456_6),.b(n465_3),.q(n1168));
  and_bi g709(.a(n707_1),.b(n701_1),.q(n709));
  or_bb g1083(.a(n1079),.b(n1082),.q(_w_6272));
  bfr _b_3893(.a(_w_5318),.q(_w_5319));
  and_bi g198(.a(G5221_7),.b(n197),.q(n198));
  or_bb g883(.a(n879),.b(n882),.q(_w_6277));
  and_bb g1088(.a(G36_1),.b(n630_10),.q(n1088));
  or_bb g216(.a(G100_13),.b(G117_0),.q(n216));
  and_bb g587(.a(G3_0),.b(n586_0),.q(n587));
  bfr _b_4140(.a(_w_5565),.q(_w_5566));
  bfr _b_7084(.a(_w_8509),.q(_w_8510));
  and_bb g998(.a(G5213_1),.b(n997),.q(n998));
  bfr _b_4725(.a(_w_6150),.q(G5290_0));
  or_bb g1479(.a(n1475),.b(n1478),.q(n1479));
  or_bb g1090(.a(n1088),.b(n1089),.q(n1090));
  bfr _b_2124(.a(_w_3549),.q(_w_3550));
  and_bb g452(.a(n445_0),.b(n451_0),.q(n452));
  bfr _b_1971(.a(_w_3396),.q(_w_3397));
  and_bb g220(.a(G102_4),.b(G117_2),.q(_w_6285));
  bfr _b_2487(.a(_w_3912),.q(_w_3913));
  bfr _b_3142(.a(_w_4567),.q(_w_4568));
  bfr _b_2172(.a(_w_3597),.q(_w_3598));
  and_bb g401(.a(n394_0),.b(n400_0),.q(n401));
  and_bi g1049(.a(G18_0),.b(n588_8),.q(n1049));
  bfr _b_3108(.a(_w_4533),.q(_w_4534));
  bfr _b_4049(.a(_w_5474),.q(n442));
  or_bb g1102(.a(G158_11),.b(G5292_4),.q(n1102));
  bfr _b_6320(.a(_w_7745),.q(_w_7746));
  bfr _b_4325(.a(_w_5750),.q(n1461));
  bfr _b_2131(.a(_w_3556),.q(_w_3557));
  bfr _b_4483(.a(_w_5908),.q(G173_2));
  bfr _b_4748(.a(_w_6173),.q(_w_6174));
  and_bb g1106(.a(G85_0),.b(n804_8),.q(n1106));
  bfr _b_7362(.a(_w_8787),.q(_w_8788));
  or_bb g1068(.a(G174_12),.b(G5291_2),.q(_w_6287));
  bfr _b_4236(.a(_w_5661),.q(_w_5662));
  spl4L g586_s_1(.a(n586_2),.q0(n586_4),.q1(n586_5),.q2(n586_6),.q3(n586_7));
  or_bb g260(.a(G121_0),.b(G169_5),.q(n260));
  bfr _b_5289(.a(_w_6714),.q(_w_6715));
  or_bb g1108(.a(n1104),.b(n1107),.q(n1108));
  and_bb g697(.a(n438_3),.b(n448_3),.q(n697));
  and_bi g725(.a(n724),.b(n723),.q(_w_5832));
  and_bb g1109(.a(G64_13),.b(n1108),.q(_w_6288));
  bfr _b_4662(.a(_w_6087),.q(_w_6088));
  bfr _b_6349(.a(_w_7774),.q(_w_7775));
  or_bb g1098(.a(n1096),.b(n1097),.q(n1098));
  bfr _b_6654(.a(_w_8079),.q(_w_8058));
  bfr _b_6212(.a(_w_7637),.q(_w_7638));
  bfr _b_3748(.a(_w_5173),.q(_w_5174));
  or_bb g1111(.a(G158_9),.b(G5291_4),.q(n1111));
  bfr _b_5949(.a(_w_7374),.q(_w_7375));
  bfr _b_5770(.a(_w_7195),.q(_w_7196));
  and_bi g969(.a(n968),.b(n962),.q(_w_5229));
  bfr _b_2216(.a(_w_3641),.q(n402_2));
  and_bi g1113(.a(n1112),.b(n1110),.q(_w_6289));
  bfr _b_6296(.a(_w_7721),.q(_w_7722));
  and_bb g1114(.a(G84_0),.b(n804_9),.q(n1114));
  bfr _b_2162(.a(_w_3587),.q(_w_3588));
  spl2 g749_s_0(.a(n749),.q0(n749_0),.q1(n749_1));
  and_bb g309(.a(n289_0),.b(n308),.q(n309));
  bfr _b_3407(.a(_w_4832),.q(_w_4833));
  bfr _b_4381(.a(_w_5806),.q(_w_5807));
  spl3L g1268_s_0(.a(n1268),.q0(n1268_0),.q1(n1268_1),.q2(n1268_2));
  and_bb g1118(.a(G64_12),.b(n1117),.q(_w_6290));
  bfr _b_3866(.a(_w_5291),.q(_w_5292));
  bfr _b_2170(.a(_w_3595),.q(_w_3596));
  bfr _b_6243(.a(_w_7668),.q(_w_7669));
  bfr _b_2672(.a(_w_4097),.q(_w_4098));
  bfr _b_4035(.a(_w_5460),.q(_w_5461));
  bfr _b_3132(.a(_w_4557),.q(G174_2));
  bfr _b_2409(.a(_w_3834),.q(_w_3835));
  and_bi g613(.a(G177_25),.b(n612),.q(n613));
  or_bb g607(.a(n452_1),.b(n594_1),.q(n607));
  and_bi g1121(.a(G159_13),.b(n1120),.q(n1121));
  or_bb g244(.a(G113_0),.b(G98_6),.q(n244));
  and_bb g1039(.a(n1036),.b(n1038),.q(_w_6292));
  bfr _b_4796(.a(_w_6221),.q(n400_2));
  bfr _b_2973(.a(_w_4398),.q(G5239_0));
  bfr _b_2165(.a(_w_3590),.q(_w_3591));
  spl4L g185_s_2(.a(G5221_3),.q0(G5221_7),.q1(G5221_8),.q2(G5221_9),.q3(G5221_10));
  spl3L g640_s_0(.a(n640),.q0(n640_0),.q1(n640_1),.q2(n640_2));
  spl2 g572_s_0(.a(n572),.q0(n572_0),.q1(n572_1));
  and_bb g1131(.a(n1128),.b(n1130),.q(_w_6294));
  and_bb g599(.a(n479_2),.b(n597_1),.q(n599));
  and_bi g1185(.a(n433_2),.b(n607_2),.q(n1185));
  bfr _b_3897(.a(_w_5322),.q(_w_5323));
  bfr _b_3442(.a(_w_4867),.q(_w_4868));
  bfr _b_2007(.a(_w_3432),.q(_w_3433));
  bfr _b_6881(.a(_w_8306),.q(_w_8307));
  bfr _b_2622(.a(_w_4047),.q(_w_4048));
  bfr _b_6363(.a(_w_7788),.q(_w_7789));
  and_bi g1132(.a(G77_1),.b(n813_7),.q(n1132));
  bfr _b_3725(.a(_w_5150),.q(_w_5151));
  and_bi g661(.a(G177_22),.b(n660),.q(_w_6295));
  and_bb g1133(.a(G87_1),.b(n815_7),.q(n1133));
  bfr _b_2809(.a(_w_4234),.q(_w_4235));
  and_bb g983(.a(n980),.b(n982),.q(n983));
  bfr _b_3903(.a(_w_5328),.q(_w_5329));
  and_bi g248(.a(G115_1),.b(G101_6),.q(_w_6296));
  bfr _b_5627(.a(_w_7052),.q(_w_7053));
  bfr _b_2912(.a(_w_4337),.q(G159_2));
  and_bi g1260(.a(G176_31),.b(n1259),.q(n1260));
  and_bi g1173(.a(n1172),.b(n1171),.q(n1173));
  bfr _b_4622(.a(_w_6047),.q(_w_6048));
  bfr _b_5768(.a(_w_7193),.q(_w_7194));
  spl4L G123_s_3(.a(G123_2),.q0(G123_12),.q1(G123_13),.q2(_w_6297),.q3(G123_15));
  and_bi g1139(.a(G161_11),.b(n1138),.q(n1139));
  and_bi g1150(.a(G74_1),.b(n813_9),.q(n1150));
  bfr _b_4852(.a(_w_6277),.q(_w_6278));
  bfr _b_5536(.a(G171),.q(_w_6962));
  spl3L G166_s_1(.a(G166_1),.q0(G166_4),.q1(G166_5),.q2(G166_6));
  or_bb g1152(.a(n1150),.b(n1151),.q(n1152));
  bfr _b_6632(.a(_w_8057),.q(_w_8036));
  bfr _b_2616(.a(_w_4041),.q(_w_4042));
  bfr _b_3814(.a(_w_5239),.q(_w_5240));
  or_bb g1153(.a(n1149),.b(n1152),.q(n1153));
  bfr _b_2481(.a(_w_3906),.q(_w_3907));
  bfr _b_7556(.a(_w_8981),.q(_w_8982));
  bfr _b_5516(.a(_w_6941),.q(_w_6942));
  spl2 g1434_s_0(.a(n1434),.q0(n1434_0),.q1(n1434_1));
  and_bi g250(.a(n246_0),.b(n249_0),.q(n250));
  bfr _b_2796(.a(_w_4221),.q(_w_4222));
  bfr _b_4856(.a(_w_6281),.q(_w_6282));
  or_bb g1285(.a(n1283),.b(n1284),.q(_w_6303));
  and_bb g1046(.a(G172_11),.b(n1045),.q(n1046));
  and_bi g1157(.a(G161_13),.b(n1156),.q(n1157));
  or_bb g1207(.a(G176_30),.b(n1206),.q(n1207));
  spl4L g630_s_0(.a(n630),.q0(n630_0),.q1(n630_1),.q2(n630_2),.q3(n630_3));
  bfr _b_2795(.a(_w_4220),.q(_w_4221));
  bfr _b_4324(.a(_w_5749),.q(_w_5750));
  bfr _b_5699(.a(_w_7124),.q(_w_7125));
  bfr _b_2044(.a(_w_3469),.q(_w_3470));
  bfr _b_3584(.a(_w_5009),.q(_w_5010));
  bfr _b_2055(.a(_w_3480),.q(_w_3481));
  or_bb g835(.a(n831),.b(n834),.q(_w_4405));
  bfr _b_4577(.a(_w_6002),.q(_w_6003));
  and_bi g1164(.a(n456_5),.b(G145_5),.q(n1164));
  bfr _b_2488(.a(_w_3913),.q(_w_3914));
  bfr _b_5873(.a(_w_7298),.q(_w_7299));
  bfr _b_4071(.a(_w_5496),.q(_w_5497));
  bfr _b_7120(.a(_w_8545),.q(_w_8546));
  bfr _b_5251(.a(_w_6676),.q(_w_6677));
  bfr _b_2469(.a(_w_3894),.q(_w_3895));
  bfr _b_2179(.a(_w_3604),.q(_w_3605));
  bfr _b_4957(.a(_w_6382),.q(_w_6383));
  or_bb g1167(.a(n1164_1),.b(n1166),.q(n1167));
  and_bi g1169(.a(n1167),.b(n1168),.q(n1169));
  or_bb g1405(.a(n1403),.b(n1404),.q(n1405));
  bfr _b_3645(.a(_w_5070),.q(_w_5071));
  or_bb g644(.a(n638),.b(n643_0),.q(n644));
  bfr _b_5343(.a(_w_6768),.q(_w_6769));
  bfr _b_4269(.a(_w_5694),.q(_w_5695));
  spl4L g462_s_0(.a(n462),.q0(n462_0),.q1(n462_1),.q2(_w_3474),.q3(_w_3476));
  and_bi g1174(.a(n773_6),.b(n1173),.q(n1174));
  or_bb g1179(.a(n1177),.b(n1178),.q(_w_6309));
  bfr _b_6906(.a(_w_8331),.q(_w_8330));
  bfr _b_4665(.a(_w_6090),.q(_w_6091));
  and_ii g625(.a(n616),.b(n624),.q(_w_6310));
  bfr _b_2627(.a(_w_4052),.q(_w_4053));
  bfr _b_2639(.a(_w_4064),.q(G149_2));
  bfr _b_2924(.a(_w_4349),.q(_w_4350));
  bfr _b_3647(.a(_w_5072),.q(_w_5073));
  or_bb g1093(.a(G158_13),.b(G5293_4),.q(n1093));
  or_bb g1181(.a(n1176_1),.b(n1179_1),.q(n1181));
  bfr _b_3968(.a(_w_5393),.q(_w_5394));
  bfr _b_4045(.a(_w_5470),.q(_w_5471));
  bfr _b_2706(.a(_w_4131),.q(_w_4132));
  spl4L G163_s_2(.a(G163_2),.q0(G163_7),.q1(G163_8),.q2(G163_9),.q3(G163_10));
  bfr _b_2963(.a(_w_4388),.q(_w_4389));
  and_bb g388(.a(n381_0),.b(n387_0),.q(n388));
  bfr _b_3338(.a(_w_4763),.q(_w_4764));
  bfr _b_2184(.a(_w_3609),.q(_w_3610));
  bfr _b_2675(.a(_w_4100),.q(G5292));
  and_bi g1186(.a(n607_3),.b(n434_2),.q(n1186));
  bfr _b_6631(.a(_w_8056),.q(_w_8057));
  bfr _b_5875(.a(_w_7300),.q(_w_7301));
  bfr _b_4767(.a(_w_6192),.q(_w_6193));
  bfr _b_2149(.a(_w_3574),.q(_w_3575));
  and_bb g1189(.a(n1188),.b(n439_2),.q(n1189));
  and_bb g1191(.a(n1190),.b(n444_1),.q(n1191));
  bfr _b_6517(.a(_w_7942),.q(_w_7943));
  bfr _b_4064(.a(_w_5489),.q(_w_5490));
  bfr _b_6534(.a(_w_7959),.q(_w_7960));
  bfr _b_2089(.a(_w_3514),.q(_w_3515));
  and_bi g1193(.a(n479_4),.b(n435_4),.q(n1193));
  spl4L G123_s_4(.a(G123_3),.q0(_w_6322),.q1(G123_17),.q2(G123_18),.q3(G123_19));
  bfr _b_5651(.a(_w_7076),.q(_w_7077));
  bfr _b_2108(.a(_w_3533),.q(_w_3534));
  or_bb g1197(.a(n1192_1),.b(n1195_1),.q(n1197));
  bfr _b_3110(.a(_w_4535),.q(_w_4536));
  bfr _b_5470(.a(_w_6895),.q(_w_6896));
  bfr _b_3713(.a(_w_5138),.q(_w_5139));
  and_bi g1473(.a(G160_5),.b(n1447_3),.q(n1473));
  bfr _b_7339(.a(_w_8764),.q(_w_8765));
  bfr _b_2027(.a(_w_3452),.q(_w_3453));
  and_bi g1200(.a(n451_5),.b(n1198_1),.q(n1200));
  spl3L g432_s_0(.a(n432),.q0(n432_0),.q1(n432_1),.q2(n432_2));
  bfr _b_2728(.a(_w_4153),.q(_w_4154));
  bfr _b_3382(.a(_w_4807),.q(_w_4808));
  and_bi g1366(.a(G140_5),.b(n1365),.q(n1366));
  bfr _b_6323(.a(_w_7748),.q(_w_7749));
  and_bb g907(.a(G71_0),.b(n804_5),.q(n907));
  and_bb g780(.a(n458_1),.b(n463_2),.q(n780));
  bfr _b_6557(.a(_w_7982),.q(_w_7983));
  bfr _b_3891(.a(_w_5316),.q(_w_5317));
  and_bi g686(.a(n685),.b(n684),.q(_w_6324));
  bfr _b_4789(.a(_w_6214),.q(n400_1));
  bfr _b_7407(.a(_w_8832),.q(_w_8833));
  or_bb g372(.a(n370),.b(n371),.q(n372));
  and_bi g1217(.a(n1215),.b(n1216),.q(n1217));
  bfr _b_5803(.a(_w_7228),.q(_w_7229));
  bfr _b_4508(.a(_w_5933),.q(n451_3));
  bfr _b_2181(.a(_w_3606),.q(n253_1));
  bfr _b_2958(.a(_w_4383),.q(_w_4384));
  bfr _b_3242(.a(_w_4667),.q(G135_4));
  and_bi g964(.a(G170_2),.b(G54_0),.q(n964));
  and_bb g443(.a(G150_4),.b(n438_1),.q(n443));
  and_bi g1220(.a(G98_9),.b(G121_13),.q(n1220));
  bfr _b_3659(.a(_w_5084),.q(_w_5085));
  or_bb g1223(.a(n1218),.b(n1222),.q(_w_6327));
  and_bi g810(.a(G160_27),.b(G5248_5),.q(n810));
  or_bb g1224(.a(n1214_0),.b(n1223_0),.q(n1224));
  or_bb g765(.a(n425_2),.b(n744_6),.q(n765));
  and_bb g1225(.a(n1214_1),.b(n1223_1),.q(n1225));
  bfr _b_2223(.a(_w_3648),.q(G143_2));
  spl2 G103_s_1(.a(G103_1),.q0(G103_4),.q1(G103_5));
  bfr _b_4820(.a(_w_6245),.q(_w_6246));
  bfr _b_3345(.a(_w_4770),.q(G160_24));
  bfr _b_2535(.a(_w_3960),.q(_w_3961));
  and_bi g1226(.a(n1224),.b(n1225),.q(n1226));
  bfr _b_4239(.a(_w_5664),.q(_w_5665));
  and_bb g436(.a(G123_23),.b(G128_7),.q(n436));
  or_bb g1119(.a(G158_8),.b(G5290_4),.q(_w_6328));
  and_bi g825(.a(G14_0),.b(n588_1),.q(n825));
  and_bi g962(.a(G171_0),.b(n961),.q(n962));
  or_bb g458(.a(G145_4),.b(n456_1),.q(n458));
  bfr _b_3060(.a(_w_4485),.q(_w_4486));
  bfr _b_3580(.a(_w_5005),.q(_w_5006));
  or_bb g1258(.a(n1250_0),.b(n1257_0),.q(_w_6329));
  bfr _b_2041(.a(_w_3466),.q(n465_2));
  spl4L G105_s_2(.a(G105_2),.q0(G105_6),.q1(_w_6330),.q2(G105_8),.q3(G105_9));
  and_bi g1439(.a(G177_7),.b(n1438),.q(_w_4270));
  or_bb g1233(.a(n1231),.b(n1232),.q(n1233));
  bfr _b_5045(.a(_w_6470),.q(_w_6471));
  bfr _b_2674(.a(_w_4099),.q(_w_4100));
  bfr _b_5847(.a(_w_7272),.q(_w_7273));
  spl4L G177_s_1(.a(G177_0),.q0(G177_4),.q1(G177_5),.q2(G177_6),.q3(_w_6331));
  bfr _b_3906(.a(_w_5331),.q(n226));
  bfr _b_5071(.a(_w_6496),.q(_w_6497));
  or_bb g874(.a(n872),.b(n873),.q(n874));
  and_bb g1240(.a(G102_10),.b(G126_12),.q(n1240));
  and_bb g989(.a(n986),.b(n988),.q(n989));
  bfr _b_6177(.a(_w_7602),.q(_w_7603));
  and_bi g1250(.a(n1248),.b(n1249),.q(_w_6335));
  or_bb g1242(.a(n1240),.b(n1241),.q(n1242));
  spl4L g386_s_0(.a(n386),.q0(n386_0),.q1(n386_1),.q2(_w_6340),.q3(n386_3));
  bfr _b_7546(.a(_w_8971),.q(_w_8972));
  bfr _b_2725(.a(_w_4150),.q(_w_4151));
  bfr _b_7074(.a(_w_8499),.q(_w_8500));
  spl4L G158_s_5(.a(G158_18),.q0(_w_3664),.q1(G158_21),.q2(_w_3665),.q3(G158_23));
  spl2 g318_s_0(.a(n318),.q0(n318_0),.q1(n318_1));
  and_bb g440(.a(G123_21),.b(G130_2),.q(n440));
  or_bb g542(.a(n539),.b(n541),.q(n542));
  bfr _b_4068(.a(_w_5493),.q(G176_43));
  and_bi g1247(.a(n1245),.b(n1246),.q(_w_6348));
  bfr _b_3317(.a(_w_4742),.q(_w_4743));
  bfr _b_4654(.a(_w_6079),.q(_w_6080));
  and_bi g1331(.a(n1330),.b(n1328),.q(n1331));
  bfr _b_2742(.a(_w_4167),.q(_w_4168));
  bfr _b_3065(.a(_w_4490),.q(_w_4491));
  and_bb g1249(.a(n1226_1),.b(n1247_1),.q(n1249));
  bfr _b_4293(.a(_w_5718),.q(_w_5719));
  and_bi g1252(.a(n1251),.b(n234_1),.q(n1252));
  bfr _b_7116(.a(_w_8541),.q(_w_8542));
  spl2 g530_s_0(.a(n530),.q0(n530_0),.q1(n530_1));
  bfr _b_3872(.a(_w_5297),.q(_w_5298));
  bfr _b_6565(.a(_w_7990),.q(_w_7991));
  or_bb g1254(.a(n1253),.b(n250_1),.q(n1254));
  spl4L g588_s_2(.a(n588_3),.q0(n588_8),.q1(n588_9),.q2(n588_10),.q3(n588_11));
  spl2 g1324_s_0(.a(n1324),.q0(_w_6349),.q1(n1324_1));
  bfr _b_6246(.a(_w_7671),.q(_w_7672));
  and_bi g1257(.a(n1255),.b(n1256),.q(n1257));
  or_bb g193(.a(n191),.b(n192),.q(n193));
  bfr _b_6504(.a(_w_7929),.q(_w_7930));
  and_bi g1130(.a(G161_10),.b(n1129),.q(n1130));
  and_bi g1343(.a(G90_11),.b(G101_12),.q(n1343));
  bfr _b_4321(.a(_w_5746),.q(_w_5747));
  and_bb g1403(.a(G102_16),.b(G96_12),.q(n1403));
  and_bb g1261(.a(n1258),.b(n1260),.q(n1261));
  bfr _b_2132(.a(_w_3557),.q(_w_3558));
  bfr _b_3483(.a(_w_4908),.q(_w_4909));
  bfr _b_3977(.a(_w_5402),.q(G5248_0));
  bfr _b_4128(.a(_w_5553),.q(_w_5554));
  bfr _b_2709(.a(_w_4134),.q(_w_4135));
  bfr _b_1942(.a(_w_3367),.q(_w_3368));
  bfr _b_2357(.a(_w_3782),.q(_w_3783));
  bfr _b_2835(.a(_w_4260),.q(G161_0));
  bfr _b_4905(.a(_w_6330),.q(G105_7));
  bfr _b_2359(.a(_w_3784),.q(_w_3785));
  bfr _b_2411(.a(_w_3836),.q(_w_3837));
  bfr _b_7213(.a(_w_8638),.q(_w_8639));
  bfr _b_6305(.a(_w_7730),.q(_w_7731));
  bfr _b_2360(.a(_w_3785),.q(_w_3786));
  bfr _b_2364(.a(_w_3789),.q(_w_3790));
  spl4L g384_s_0(.a(n384),.q0(n384_0),.q1(n384_1),.q2(n384_2),.q3(n384_3));
  bfr _b_2365(.a(_w_3790),.q(_w_3791));
  bfr _b_7276(.a(_w_8701),.q(_w_8702));
  bfr _b_3260(.a(_w_4685),.q(_w_4686));
  bfr _b_2367(.a(_w_3792),.q(_w_3793));
  bfr _b_2369(.a(_w_3794),.q(_w_3795));
  bfr _b_2370(.a(_w_3795),.q(_w_3796));
  bfr _b_4696(.a(_w_6121),.q(_w_6122));
  bfr _b_2371(.a(_w_3796),.q(_w_3797));
  bfr _b_2372(.a(_w_3797),.q(_w_3798));
  bfr _b_2373(.a(_w_3798),.q(_w_3799));
  bfr _b_5109(.a(_w_6534),.q(_w_6531));
  bfr _b_2374(.a(_w_3799),.q(_w_3800));
  and_bb g303(.a(G167_8),.b(G92_5),.q(n303));
  bfr _b_3632(.a(_w_5057),.q(_w_5058));
  bfr _b_4464(.a(_w_5889),.q(_w_5890));
  bfr _b_2379(.a(_w_3804),.q(n375_0));
  bfr _b_6795(.a(_w_8220),.q(_w_8221));
  bfr _b_2380(.a(_w_3805),.q(_w_3806));
  bfr _b_2381(.a(_w_3806),.q(_w_3807));
  bfr _b_2382(.a(_w_3807),.q(n375_2));
  bfr _b_5509(.a(_w_6934),.q(_w_6935));
  bfr _b_5169(.a(_w_6594),.q(_w_6595));
  bfr _b_2383(.a(_w_3808),.q(_w_3809));
  bfr _b_2385(.a(_w_3810),.q(_w_3811));
  and_bb g819(.a(G64_24),.b(n818),.q(G5266));
  bfr _b_2386(.a(_w_3811),.q(_w_3812));
  spl2 G17_s_0(.a(_w_6916),.q0(G17_0),.q1(G17_1));
  bfr _b_2387(.a(_w_3812),.q(_w_3813));
  bfr _b_7201(.a(_w_8626),.q(_w_8627));
  bfr _b_2571(.a(_w_3996),.q(_w_3997));
  bfr _b_2388(.a(_w_3813),.q(n453_0));
  bfr _b_3086(.a(_w_4511),.q(_w_4512));
  bfr _b_6389(.a(_w_7814),.q(_w_7815));
  bfr _b_2389(.a(_w_3814),.q(_w_3815));
  bfr _b_5310(.a(_w_6735),.q(_w_6704));
  and_bb g430(.a(n409_0),.b(n429_0),.q(n430));
  bfr _b_2390(.a(_w_3815),.q(n419_1));
  bfr _b_6098(.a(_w_7523),.q(_w_7524));
  bfr _b_2454(.a(_w_3879),.q(_w_3880));
  bfr _b_6872(.a(_w_8297),.q(_w_8298));
  bfr _b_3251(.a(_w_4676),.q(n277_1));
  bfr _b_2391(.a(_w_3816),.q(_w_3817));
  bfr _b_4568(.a(_w_5993),.q(_w_5994));
  or_bb g1298(.a(n428_2),.b(n545_2),.q(n1298));
  bfr _b_2392(.a(_w_3817),.q(_w_3818));
  bfr _b_2393(.a(_w_3818),.q(_w_3819));
  spl4L g632_s_1(.a(n632_2),.q0(n632_4),.q1(n632_5),.q2(n632_6),.q3(n632_7));
  bfr _b_2394(.a(_w_3819),.q(_w_3820));
  bfr _b_2875(.a(_w_4300),.q(_w_4301));
  bfr _b_3990(.a(_w_5415),.q(_w_5416));
  bfr _b_2396(.a(_w_3821),.q(_w_3822));
  bfr _b_2993(.a(_w_4418),.q(_w_4419));
  bfr _b_2791(.a(_w_4216),.q(_w_4217));
  bfr _b_2397(.a(_w_3822),.q(_w_3823));
  bfr _b_2398(.a(_w_3823),.q(_w_3824));
  bfr _b_2399(.a(_w_3824),.q(_w_3825));
  and_bi g476(.a(n474_0),.b(n475),.q(n476));
  bfr _b_2540(.a(_w_3965),.q(_w_3966));
  bfr _b_2533(.a(_w_3958),.q(_w_3959));
  bfr _b_6173(.a(_w_7598),.q(_w_7599));
  bfr _b_5409(.a(_w_6834),.q(_w_6835));
  bfr _b_3160(.a(_w_4585),.q(_w_4586));
  bfr _b_2220(.a(_w_3645),.q(G141_4));
  bfr _b_2404(.a(_w_3829),.q(_w_3830));
  bfr _b_3784(.a(_w_5209),.q(_w_5210));
  bfr _b_6553(.a(_w_7978),.q(_w_7979));
  bfr _b_2405(.a(_w_3830),.q(_w_3831));
  bfr _b_2407(.a(_w_3832),.q(_w_3833));
  bfr _b_2045(.a(_w_3470),.q(_w_3471));
  bfr _b_2408(.a(_w_3833),.q(_w_3834));
  bfr _b_6009(.a(_w_7434),.q(_w_7435));
  bfr _b_2410(.a(_w_3835),.q(_w_3836));
  bfr _b_4834(.a(_w_6259),.q(_w_6260));
  bfr _b_4871(.a(_w_6296),.q(n248));
  bfr _b_2413(.a(_w_3838),.q(_w_3839));
  and_bi g1409(.a(G109_11),.b(G101_18),.q(n1409));
  bfr _b_2078(.a(_w_3503),.q(n443_3));
  bfr _b_2415(.a(_w_3840),.q(_w_3841));
  bfr _b_2416(.a(_w_3841),.q(_w_3842));
  bfr _b_2418(.a(_w_3843),.q(_w_3844));
  bfr _b_2425(.a(_w_3850),.q(_w_3851));
  bfr _b_4868(.a(_w_6293),.q(G5305));
  and_bb g419(.a(G144_2),.b(n418_0),.q(n419));
  bfr _b_3796(.a(_w_5221),.q(_w_5222));
  bfr _b_2419(.a(_w_3844),.q(_w_3845));
  bfr _b_6615(.a(_w_8040),.q(_w_8041));
  bfr _b_6156(.a(_w_7581),.q(_w_7582));
  bfr _b_2421(.a(_w_3846),.q(_w_3847));
  bfr _b_5648(.a(_w_7073),.q(_w_7074));
  bfr _b_2422(.a(_w_3847),.q(_w_3848));
  bfr _b_2423(.a(_w_3848),.q(_w_3849));
  bfr _b_2424(.a(_w_3849),.q(_w_3850));
  bfr _b_2430(.a(_w_3855),.q(_w_3856));
  bfr _b_2432(.a(_w_3857),.q(_w_3858));
  bfr _b_2434(.a(_w_3859),.q(_w_3860));
  or_bb g692(.a(n690),.b(n691),.q(n692));
  bfr _b_4726(.a(_w_6151),.q(_w_6152));
  bfr _b_2436(.a(_w_3861),.q(_w_3862));
  bfr _b_2437(.a(_w_3862),.q(_w_3863));
  bfr _b_4533(.a(_w_5958),.q(_w_5959));
  and_bi g722(.a(n720),.b(n721),.q(_w_5156));
  bfr _b_3027(.a(_w_4452),.q(_w_4453));
  bfr _b_2440(.a(_w_3865),.q(_w_3866));
  bfr _b_5486(.a(_w_6911),.q(_w_6912));
  bfr _b_2442(.a(_w_3867),.q(_w_3868));
  bfr _b_2443(.a(_w_3868),.q(_w_3869));
  bfr _b_2446(.a(_w_3871),.q(_w_3872));
  or_bb g582(.a(G173_15),.b(G5250_1),.q(n582));
  bfr _b_2576(.a(_w_4001),.q(n472_7));
  or_bb g1333(.a(n394_5),.b(n400_5),.q(n1333));
  bfr _b_3739(.a(_w_5164),.q(_w_5165));
  and_bi g311(.a(G109_4),.b(G168_9),.q(n311));
  bfr _b_2447(.a(_w_3872),.q(_w_3873));
  and_bb g482(.a(n453_0),.b(n481),.q(_w_4383));
  bfr _b_2448(.a(_w_3873),.q(_w_3874));
  bfr _b_5148(.a(_w_6573),.q(_w_6574));
  bfr _b_2449(.a(_w_3874),.q(_w_3875));
  bfr _b_3629(.a(_w_5054),.q(_w_5055));
  bfr _b_3998(.a(_w_5423),.q(_w_5424));
  bfr _b_2451(.a(_w_3876),.q(_w_3877));
  bfr _b_3350(.a(_w_4775),.q(_w_4776));
  bfr _b_2452(.a(_w_3877),.q(_w_3878));
  bfr _b_6982(.a(_w_8407),.q(_w_8408));
  bfr _b_3984(.a(_w_5409),.q(_w_5410));
  bfr _b_2456(.a(_w_3881),.q(_w_3882));
  bfr _b_3754(.a(_w_5179),.q(_w_5180));
  bfr _b_3837(.a(_w_5262),.q(_w_5263));
  bfr _b_2457(.a(_w_3882),.q(_w_3883));
  bfr _b_7042(.a(_w_8467),.q(_w_8434));
  bfr _b_4196(.a(_w_5621),.q(_w_5622));
  bfr _b_2459(.a(_w_3884),.q(_w_3885));
  bfr _b_5157(.a(_w_6582),.q(_w_6583));
  bfr _b_3822(.a(_w_5247),.q(G5283));
  bfr _b_2460(.a(_w_3885),.q(_w_3886));
  bfr _b_2462(.a(_w_3887),.q(G114_1));
  bfr _b_4091(.a(_w_5516),.q(_w_5517));
  bfr _b_2464(.a(_w_3889),.q(_w_3890));
  bfr _b_7413(.a(_w_8838),.q(_w_8839));
  bfr _b_6354(.a(_w_7779),.q(_w_7780));
  bfr _b_2949(.a(_w_4374),.q(_w_4375));
  bfr _b_3450(.a(_w_4875),.q(_w_4876));
  bfr _b_2467(.a(_w_3892),.q(_w_3893));
  bfr _b_2468(.a(_w_3893),.q(G2_2));
  bfr _b_6524(.a(_w_7949),.q(_w_7950));
  bfr _b_2471(.a(_w_3896),.q(G2_3));
  bfr _b_2473(.a(_w_3898),.q(_w_3899));
  bfr _b_2476(.a(_w_3901),.q(_w_3902));
  bfr _b_2477(.a(_w_3902),.q(_w_3903));
  bfr _b_4844(.a(_w_6269),.q(_w_6270));
  and_bi g1209(.a(G98_8),.b(G148_5),.q(n1209));
  bfr _b_2480(.a(_w_3905),.q(G128_7));
  and_bi g498(.a(G126_8),.b(G128_8),.q(n498));
  bfr _b_2483(.a(_w_3908),.q(_w_3909));
  bfr _b_2484(.a(_w_3909),.q(_w_3910));
  bfr _b_5643(.a(_w_7068),.q(_w_7069));
  bfr _b_2485(.a(_w_3910),.q(_w_3911));
  bfr _b_3763(.a(_w_5188),.q(_w_5189));
  bfr _b_6026(.a(_w_7451),.q(_w_7452));
  or_bb g516(.a(G103_8),.b(G96_8),.q(n516));
  bfr _b_4150(.a(_w_5575),.q(_w_5576));
  and_bb g606(.a(_w_8058),.b(n552_22),.q(n606));
  and_bb g1136(.a(G64_10),.b(n1135),.q(_w_5758));
  bfr _b_2486(.a(_w_3911),.q(_w_3912));
  bfr _b_2032(.a(_w_3457),.q(_w_3458));
  bfr _b_2819(.a(_w_4244),.q(_w_4245));
  bfr _b_4460(.a(_w_5885),.q(_w_5886));
  bfr _b_2489(.a(_w_3914),.q(_w_3915));
  bfr _b_2490(.a(_w_3915),.q(n346_1));
  bfr _b_2492(.a(_w_3917),.q(_w_3918));
  spl2 g1179_s_0(.a(n1179),.q0(n1179_0),.q1(n1179_1));
  inv inv_G131(.a(G131_1),.q(G5198));
  bfr _b_2493(.a(_w_3918),.q(_w_3919));
  bfr _b_2649(.a(_w_4074),.q(_w_4075));
  bfr _b_5877(.a(_w_7302),.q(_w_7303));
  and_bi g718(.a(n378_3),.b(n384_3),.q(n718));
  bfr _b_4466(.a(_w_5891),.q(_w_5892));
  bfr _b_2494(.a(_w_3919),.q(_w_3920));
  and_bb g772(.a(n478_1),.b(n597_2),.q(n772));
  bfr _b_3608(.a(_w_5033),.q(_w_5034));
  bfr _b_2498(.a(_w_3923),.q(_w_3924));
  bfr _b_6886(.a(_w_8311),.q(_w_8312));
  bfr _b_5225(.a(_w_6650),.q(_w_6651));
  spl2 g650_s_1(.a(G5257_3),.q0(G5257_4),.q1(G5257_5));
  bfr _b_2499(.a(_w_3924),.q(_w_3925));
  bfr _b_2500(.a(_w_3925),.q(n234_0));
  bfr _b_2501(.a(_w_3926),.q(_w_3927));
  bfr _b_3424(.a(_w_4849),.q(_w_4850));
  bfr _b_4298(.a(_w_5723),.q(_w_5724));
  bfr _b_2503(.a(_w_3928),.q(_w_3929));
  bfr _b_4594(.a(_w_6019),.q(G5250_0));
  bfr _b_3665(.a(_w_5090),.q(_w_5091));
  bfr _b_4226(.a(_w_5651),.q(_w_5652));
  bfr _b_4889(.a(_w_6314),.q(_w_6315));
  bfr _b_2504(.a(_w_3929),.q(_w_3930));
  bfr _b_3156(.a(_w_4581),.q(_w_4582));
  bfr _b_5340(.a(_w_6765),.q(_w_6766));
  bfr _b_2243(.a(_w_3668),.q(_w_3669));
  bfr _b_3257(.a(_w_4682),.q(_w_4683));
  bfr _b_2507(.a(_w_3932),.q(G123_11));
  bfr _b_2508(.a(_w_3933),.q(_w_3934));
  bfr _b_4742(.a(_w_6167),.q(n1276));
  bfr _b_2509(.a(_w_3934),.q(G123_4));
  bfr _b_5987(.a(_w_7412),.q(_w_7411));
  bfr _b_2510(.a(_w_3935),.q(G123_2));
  bfr _b_2511(.a(_w_3936),.q(n456_1));
  bfr _b_3831(.a(_w_5256),.q(n406));
  bfr _b_5435(.a(_w_6860),.q(_w_6861));
  bfr _b_2518(.a(_w_3943),.q(G88_2));
  bfr _b_2975(.a(_w_4400),.q(_w_4401));
  bfr _b_6533(.a(_w_7958),.q(_w_7959));
  bfr _b_4776(.a(_w_6201),.q(n1022));
  bfr _b_2520(.a(_w_3945),.q(G92_3));
  and_bi g1432(.a(n1431_0),.b(n1398_0),.q(n1432));
  bfr _b_2521(.a(_w_3946),.q(_w_3947));
  bfr _b_6336(.a(_w_7761),.q(_w_7762));
  bfr _b_2522(.a(_w_3947),.q(_w_3948));
  bfr _b_2525(.a(_w_3950),.q(_w_3951));
  bfr _b_2531(.a(_w_3956),.q(_w_3957));
  bfr _b_3772(.a(_w_5197),.q(_w_5198));
  bfr _b_3809(.a(_w_5234),.q(_w_5235));
  bfr _b_2536(.a(_w_3961),.q(_w_3962));
  bfr _b_2539(.a(_w_3964),.q(_w_3965));
  bfr _b_2541(.a(_w_3966),.q(_w_3967));
  bfr _b_7554(.a(_w_8979),.q(_w_8980));
  bfr _b_2543(.a(_w_3968),.q(_w_3969));
  bfr _b_5686(.a(_w_7111),.q(_w_7112));
  bfr _b_2806(.a(_w_4231),.q(n435_2));
  spl3L G137_s_1(.a(G137_3),.q0(_w_3981),.q1(G137_5),.q2(G137_6));
  bfr _b_4308(.a(_w_5733),.q(_w_5734));
  bfr _b_2550(.a(_w_3975),.q(_w_3976));
  bfr _b_2552(.a(_w_3977),.q(_w_3978));
  bfr _b_4994(.a(G118),.q(_w_6420));
  bfr _b_2553(.a(_w_3978),.q(_w_3979));
  bfr _b_3526(.a(_w_4951),.q(_w_4952));
  bfr _b_2555(.a(_w_3980),.q(n394_4));
  bfr _b_7364(.a(_w_8789),.q(_w_8790));
  bfr _b_6540(.a(_w_7965),.q(_w_7966));
  or_bb g318(.a(n313),.b(n317),.q(_w_4863));
  bfr _b_2556(.a(_w_3981),.q(G137_4));
  bfr _b_6763(.a(_w_8188),.q(_w_8189));
  or_bb g247(.a(G100_20),.b(G115_0),.q(n247));
  bfr _b_3186(.a(_w_4611),.q(_w_4612));
  bfr _b_2557(.a(_w_3982),.q(_w_3983));
  bfr _b_2558(.a(_w_3983),.q(_w_3984));
  bfr _b_2560(.a(_w_3985),.q(_w_3986));
  bfr _b_2561(.a(_w_3986),.q(_w_3987));
  and_ii g579(.a(n571),.b(n578),.q(_w_6013));
  bfr _b_3962(.a(_w_5387),.q(G5249));
  bfr _b_2324(.a(_w_3749),.q(_w_3750));
  bfr _b_2563(.a(_w_3988),.q(_w_3989));
  bfr _b_2083(.a(_w_3508),.q(_w_3509));
  bfr _b_2568(.a(_w_3993),.q(_w_3994));
  spl2 g779_s_0(.a(n779),.q0(_w_3443),.q1(n779_1));
  bfr _b_2653(.a(_w_4078),.q(_w_4079));
  bfr _b_2570(.a(_w_3995),.q(_w_3996));
  bfr _b_2572(.a(_w_3997),.q(_w_3998));
  bfr _b_2577(.a(_w_4002),.q(n442_4));
  bfr _b_3353(.a(_w_4778),.q(_w_4779));
  bfr _b_4060(.a(_w_5485),.q(n911));
  bfr _b_2583(.a(_w_4008),.q(_w_4009));
  bfr _b_4053(.a(_w_5478),.q(_w_5479));
  bfr _b_4993(.a(_w_6418),.q(_w_6417));
  bfr _b_2584(.a(_w_4009),.q(G5243));
  bfr _b_7433(.a(_w_8858),.q(_w_8859));
  bfr _b_2586(.a(_w_4011),.q(_w_4012));
  or_bb g1162(.a(n1158),.b(n1161),.q(_w_6308));
  bfr _b_2588(.a(_w_4013),.q(_w_4014));
  bfr _b_5569(.a(_w_6994),.q(_w_6995));
  and_bi g1194(.a(n435_5),.b(n479_5),.q(n1194));
  bfr _b_3931(.a(_w_5356),.q(_w_5357));
  bfr _b_2591(.a(_w_4016),.q(_w_4017));
  spl2 g464_s_1(.a(n464_3),.q0(n464_4),.q1(n464_5));
  bfr _b_2592(.a(_w_4017),.q(G5254));
  spl2 g610_s_0(.a(n610),.q0(n610_0),.q1(_w_3444));
  bfr _b_2593(.a(_w_4018),.q(_w_4019));
  bfr _b_7096(.a(_w_8521),.q(_w_8522));
  bfr _b_2595(.a(_w_4020),.q(_w_4021));
  spl4L G66_s_0(.a(_w_8187),.q0(_w_5468),.q1(G66_0),.q2(G66_1),.q3(G66_2));
  bfr _b_2395(.a(_w_3820),.q(_w_3821));
  bfr _b_2596(.a(_w_4021),.q(_w_4022));
  bfr _b_2597(.a(_w_4022),.q(_w_4023));
  bfr _b_4585(.a(_w_6010),.q(G5284));
  bfr _b_6532(.a(_w_7957),.q(_w_7958));
  bfr _b_3838(.a(_w_5263),.q(_w_5264));
  bfr _b_2479(.a(_w_3904),.q(G54_1));
  bfr _b_2599(.a(_w_4024),.q(_w_4025));
  bfr _b_2600(.a(_w_4025),.q(G5258));
  bfr _b_2602(.a(_w_4027),.q(_w_4028));
  bfr _b_2605(.a(_w_4030),.q(_w_4031));
  bfr _b_2607(.a(_w_4032),.q(_w_4033));
  bfr _b_7097(.a(_w_8522),.q(_w_8523));
  bfr _b_4409(.a(_w_5834),.q(_w_5835));
  bfr _b_2611(.a(_w_4036),.q(_w_4037));
  bfr _b_5388(.a(_w_6813),.q(_w_6814));
  bfr _b_2614(.a(_w_4039),.q(_w_4040));
  spl4L G159_s_2(.a(G159_2),.q0(G159_7),.q1(G159_8),.q2(G159_9),.q3(G159_10));
  bfr _b_3858(.a(_w_5283),.q(_w_5284));
  bfr _b_4637(.a(_w_6062),.q(_w_6063));
  bfr _b_2617(.a(_w_4042),.q(_w_4043));
  bfr _b_3076(.a(_w_4501),.q(_w_4502));
  bfr _b_2235(.a(_w_3660),.q(_w_3661));
  bfr _b_2618(.a(_w_4043),.q(_w_4044));
  bfr _b_3336(.a(_w_4761),.q(_w_4762));
  bfr _b_2619(.a(_w_4044),.q(_w_4045));
  spl3L G148_s_1(.a(G148_3),.q0(_w_3742),.q1(G148_5),.q2(G148_6));
  and_bi g455(.a(_w_6419),.b(G123_15),.q(_w_4674));
  bfr _b_2620(.a(_w_4045),.q(_w_4046));
  bfr _b_2431(.a(_w_3856),.q(_w_3857));
  bfr _b_2623(.a(_w_4048),.q(_w_4049));
  bfr _b_4406(.a(_w_5831),.q(G5270));
  bfr _b_2624(.a(_w_4049),.q(_w_4050));
  bfr _b_2625(.a(_w_4050),.q(_w_4051));
  bfr _b_2678(.a(_w_4103),.q(_w_4104));
  bfr _b_5002(.a(_w_6427),.q(_w_6425));
  bfr _b_2630(.a(_w_4055),.q(_w_4056));
  bfr _b_5564(.a(_w_6989),.q(_w_6990));
  bfr _b_2631(.a(_w_4056),.q(_w_4057));
  bfr _b_3841(.a(_w_5266),.q(_w_5267));
  bfr _b_2633(.a(_w_4058),.q(_w_4059));
  bfr _b_2634(.a(_w_4059),.q(_w_4060));
  bfr _b_4891(.a(_w_6316),.q(G5255_0));
  bfr _b_2635(.a(_w_4060),.q(_w_4061));
  bfr _b_4982(.a(G112),.q(_w_6408));
  bfr _b_2579(.a(_w_4004),.q(_w_4005));
  bfr _b_3611(.a(_w_5036),.q(_w_5037));
  bfr _b_3819(.a(_w_5244),.q(_w_5245));
  bfr _b_2640(.a(_w_4065),.q(_w_4066));
  bfr _b_2645(.a(_w_4070),.q(_w_4071));
  bfr _b_2752(.a(_w_4177),.q(_w_4178));
  bfr _b_6709(.a(G61),.q(_w_8135));
  bfr _b_2646(.a(_w_4071),.q(_w_4072));
  bfr _b_2930(.a(_w_4355),.q(_w_4356));
  bfr _b_5273(.a(_w_6698),.q(_w_6699));
  bfr _b_4524(.a(_w_5949),.q(_w_5950));
  bfr _b_2659(.a(_w_4084),.q(_w_4085));
  bfr _b_4323(.a(_w_5748),.q(n337));
  bfr _b_2662(.a(_w_4087),.q(_w_4088));
  bfr _b_3246(.a(_w_4671),.q(_w_4672));
  bfr _b_2755(.a(_w_4180),.q(n434_2));
  and_bi g1436(.a(n1377_1),.b(n1434_1),.q(_w_5767));
  bfr _b_2815(.a(_w_4240),.q(_w_4241));
  bfr _b_7391(.a(_w_8816),.q(_w_8817));
  bfr _b_3476(.a(_w_4901),.q(_w_4902));
  bfr _b_2665(.a(_w_4090),.q(_w_4091));
  bfr _b_6930(.a(_w_8355),.q(_w_8356));
  bfr _b_4305(.a(_w_5730),.q(_w_5731));
  bfr _b_3789(.a(_w_5214),.q(_w_5215));
  bfr _b_2676(.a(_w_4101),.q(_w_4102));
  bfr _b_5805(.a(_w_7230),.q(_w_7231));
  bfr _b_2677(.a(_w_4102),.q(_w_4103));
  and_bb g660(.a(G176_50),.b(n356_1),.q(n660));
  bfr _b_2679(.a(_w_4104),.q(_w_4105));
  bfr _b_3224(.a(_w_4649),.q(_w_4650));
  bfr _b_5278(.a(_w_6703),.q(_w_6672));
  bfr _b_3829(.a(_w_5254),.q(_w_5255));
  bfr _b_2680(.a(_w_4105),.q(n246_2));
  bfr _b_3753(.a(_w_5178),.q(_w_5179));
  bfr _b_5975(.a(_w_7400),.q(_w_7401));
  bfr _b_2681(.a(_w_4106),.q(_w_4107));
  bfr _b_2682(.a(_w_4107),.q(n479_0));
  bfr _b_2670(.a(_w_4095),.q(_w_4096));
  bfr _b_4589(.a(_w_6014),.q(_w_6015));
  bfr _b_2684(.a(_w_4109),.q(_w_4110));
  bfr _b_5060(.a(_w_6485),.q(_w_6486));
  bfr _b_2537(.a(_w_3962),.q(G5199));
  bfr _b_3296(.a(_w_4721),.q(_w_4722));
  bfr _b_2685(.a(_w_4110),.q(_w_4111));
  bfr _b_3529(.a(_w_4954),.q(_w_4955));
  spl2 G121_s_1(.a(G121_1),.q0(G121_4),.q1(G121_5));
  bfr _b_4704(.a(_w_6129),.q(_w_6130));
  bfr _b_2686(.a(_w_4111),.q(_w_4112));
  bfr _b_3249(.a(_w_4674),.q(n455));
  bfr _b_4174(.a(_w_5599),.q(_w_5600));
  bfr _b_2691(.a(_w_4116),.q(_w_4117));
  bfr _b_2693(.a(_w_4118),.q(_w_4119));
  or_bb g412(.a(n410),.b(n411),.q(n412));
  bfr _b_4085(.a(_w_5510),.q(_w_5511));
  bfr _b_5175(.a(_w_6600),.q(_w_6601));
  bfr _b_2694(.a(_w_4119),.q(_w_4120));
  bfr _b_2696(.a(_w_4121),.q(_w_4122));
  bfr _b_2697(.a(_w_4122),.q(_w_4123));
  bfr _b_2699(.a(_w_4124),.q(_w_4125));
  bfr _b_2702(.a(_w_4127),.q(_w_4128));
  and_bb g887(.a(n884),.b(n886),.q(n887));
  bfr _b_2703(.a(_w_4128),.q(_w_4129));
  bfr _b_2547(.a(_w_3972),.q(n537_0));
  bfr _b_4109(.a(_w_5534),.q(_w_5535));
  bfr _b_2704(.a(_w_4129),.q(_w_4130));
  and_bb g745(.a(n429_1),.b(n744_0),.q(n745));
  bfr _b_2708(.a(_w_4133),.q(n365_1));
  bfr _b_2711(.a(_w_4136),.q(n414_1));
  bfr _b_2713(.a(_w_4138),.q(_w_4139));
  spl4L G90_s_2(.a(G90_2),.q0(G90_6),.q1(G90_7),.q2(G90_8),.q3(G90_9));
  bfr _b_2714(.a(_w_4139),.q(_w_4140));
  bfr _b_2715(.a(_w_4140),.q(_w_4141));
  bfr _b_3974(.a(_w_5399),.q(_w_5400));
  bfr _b_2718(.a(_w_4143),.q(G160_20));
  bfr _b_3385(.a(_w_4810),.q(_w_4811));
  bfr _b_2719(.a(_w_4144),.q(G160_22));
  bfr _b_2913(.a(_w_4338),.q(_w_4339));
  bfr _b_4956(.a(_w_6381),.q(_w_6382));
  bfr _b_5416(.a(_w_6841),.q(_w_6842));
  bfr _b_2722(.a(_w_4147),.q(G160_6));
  bfr _b_5438(.a(_w_6863),.q(_w_6864));
  bfr _b_1980(.a(_w_3405),.q(_w_3406));
  bfr _b_2724(.a(_w_4149),.q(_w_4150));
  bfr _b_3105(.a(_w_4530),.q(_w_4531));
  bfr _b_2726(.a(_w_4151),.q(_w_4152));
  bfr _b_4730(.a(_w_6155),.q(_w_6156));
  bfr _b_2566(.a(_w_3991),.q(n472_6));
  bfr _b_3386(.a(_w_4811),.q(_w_4812));
  bfr _b_5728(.a(G19),.q(_w_7154));
  bfr _b_2737(.a(_w_4162),.q(_w_4163));
  bfr _b_4088(.a(_w_5513),.q(_w_5514));
  bfr _b_5551(.a(_w_6976),.q(_w_6977));
  bfr _b_2739(.a(_w_4164),.q(_w_4165));
  bfr _b_7353(.a(_w_8778),.q(_w_8779));
  bfr _b_2741(.a(_w_4166),.q(_w_4167));
  bfr _b_3453(.a(_w_4878),.q(_w_4879));
  bfr _b_2744(.a(_w_4169),.q(_w_4170));
  bfr _b_2745(.a(_w_4170),.q(G5251));
  bfr _b_4898(.a(_w_6323),.q(G123_16));
  bfr _b_2748(.a(_w_4173),.q(_w_4174));
  bfr _b_7383(.a(_w_8808),.q(_w_8809));
  bfr _b_4278(.a(_w_5703),.q(n1044));
  bfr _b_2749(.a(_w_4174),.q(n307_1));
  bfr _b_4922(.a(_w_6347),.q(n386_2));
  bfr _b_2750(.a(_w_4175),.q(n434_1));
  bfr _b_2753(.a(_w_4178),.q(_w_4179));
  bfr _b_4452(.a(_w_5877),.q(n463_2));
  bfr _b_3749(.a(_w_5174),.q(_w_5175));
  bfr _b_2754(.a(_w_4179),.q(_w_4180));
  and_bi g1032(.a(G41_0),.b(n632_7),.q(n1032));
  bfr _b_2782(.a(_w_4207),.q(_w_4208));
  bfr _b_3015(.a(_w_4440),.q(_w_4441));
  bfr _b_2756(.a(_w_4181),.q(n380_2));
  bfr _b_6447(.a(_w_7872),.q(_w_7873));
  bfr _b_2758(.a(_w_4183),.q(_w_4184));
  bfr _b_7535(.a(_w_8960),.q(_w_8961));
  bfr _b_4750(.a(_w_6175),.q(_w_6176));
  bfr _b_4335(.a(_w_5760),.q(_w_5761));
  bfr _b_3777(.a(_w_5202),.q(_w_5203));
  and_bi g211(.a(_w_7411),.b(G163_13),.q(_w_5475));
  bfr _b_2766(.a(_w_4191),.q(n415_0));
  bfr _b_2767(.a(_w_4192),.q(_w_4193));
  spl4L G143_s_0(.a(_w_6535),.q0(G143_0),.q1(G143_1),.q2(_w_3648),.q3(G143_3));
  bfr _b_2960(.a(_w_4385),.q(_w_4386));
  bfr _b_5696(.a(_w_7121),.q(_w_7122));
  bfr _b_2768(.a(_w_4193),.q(_w_4194));
  and_bb g352(.a(G103_5),.b(G167_12),.q(n352));
  bfr _b_4943(.a(_w_6368),.q(_w_6369));
  bfr _b_2771(.a(_w_4196),.q(_w_4197));
  bfr _b_2773(.a(_w_4198),.q(_w_4199));
  bfr _b_4061(.a(_w_5486),.q(_w_5487));
  spl4L g479_s_0(.a(n479),.q0(_w_4106),.q1(_w_4108),.q2(_w_4113),.q3(n479_3));
  bfr _b_2774(.a(_w_4199),.q(_w_4200));
  bfr _b_2776(.a(_w_4201),.q(_w_4202));
  and_bi g1216(.a(G121_11),.b(G101_9),.q(n1216));
  bfr _b_2683(.a(_w_4108),.q(_w_4109));
  bfr _b_2784(.a(_w_4209),.q(_w_4210));
  bfr _b_2573(.a(_w_3998),.q(_w_3999));
  bfr _b_2787(.a(_w_4212),.q(_w_4213));
  bfr _b_2788(.a(_w_4213),.q(_w_4214));
  and_bb g1140(.a(n1137),.b(n1139),.q(_w_6300));
  bfr _b_2918(.a(_w_4343),.q(n695));
  bfr _b_5158(.a(_w_6583),.q(_w_6584));
  bfr _b_1955(.a(_w_3380),.q(G176_49));
  bfr _b_3956(.a(_w_5381),.q(_w_5382));
  bfr _b_5706(.a(_w_7131),.q(_w_7132));
  bfr _b_2789(.a(_w_4214),.q(_w_4215));
  bfr _b_3702(.a(_w_5127),.q(_w_5128));
  and_bb g399(.a(G137_4),.b(n397_1),.q(n399));
  bfr _b_4121(.a(_w_5546),.q(_w_5547));
  bfr _b_4827(.a(_w_6252),.q(_w_6253));
  bfr _b_2798(.a(_w_4223),.q(_w_4224));
  bfr _b_4295(.a(_w_5720),.q(_w_5721));
  bfr _b_2799(.a(_w_4224),.q(n433_2));
  bfr _b_7194(.a(_w_8619),.q(_w_8620));
  bfr _b_2800(.a(_w_4225),.q(n435_0));
  bfr _b_6418(.a(_w_7843),.q(_w_7844));
  bfr _b_2801(.a(_w_4226),.q(_w_4227));
  bfr _b_2804(.a(_w_4229),.q(_w_4230));
  bfr _b_7447(.a(_w_8872),.q(_w_8873));
  and_bi g1305(.a(n1304),.b(n544_1),.q(n1305));
  and_bb g534(.a(n379_1),.b(n385_1),.q(n534));
  bfr _b_2805(.a(_w_4230),.q(_w_4231));
  bfr _b_3744(.a(_w_5169),.q(_w_5170));
  bfr _b_2810(.a(_w_4235),.q(_w_4236));
  and_bi g1274(.a(n1272_1),.b(n537_6),.q(n1274));
  bfr _b_2813(.a(_w_4238),.q(_w_4239));
  bfr _b_2816(.a(_w_4241),.q(G172_0));
  bfr _b_5461(.a(_w_6886),.q(_w_6887));
  bfr _b_2818(.a(_w_4243),.q(G172_2));
  bfr _b_4371(.a(_w_5796),.q(_w_5797));
  bfr _b_3230(.a(_w_4655),.q(G175_14));
  bfr _b_2821(.a(_w_4246),.q(G138_4));
  bfr _b_2647(.a(_w_4072),.q(G5288));
  bfr _b_4991(.a(_w_6416),.q(_w_6415));
  bfr _b_2669(.a(_w_4094),.q(_w_4095));
  bfr _b_2824(.a(_w_4249),.q(_w_4250));
  bfr _b_2826(.a(_w_4251),.q(_w_4252));
  bfr _b_2831(.a(_w_4256),.q(G5312));
  bfr _b_2832(.a(_w_4257),.q(G105_0));
  bfr _b_3275(.a(_w_4700),.q(n206));
  bfr _b_2940(.a(_w_4365),.q(_w_4366));
  bfr _b_6690(.a(_w_8115),.q(_w_8116));
  bfr _b_2833(.a(_w_4258),.q(G105_3));
  or_bb g298(.a(n293),.b(n297),.q(_w_4903));
  bfr _b_2834(.a(_w_4259),.q(_w_4260));
  bfr _b_2836(.a(_w_4261),.q(_w_4262));
  bfr _b_2837(.a(_w_4262),.q(G161_2));
  bfr _b_2838(.a(_w_4263),.q(_w_4264));
  bfr _b_2840(.a(_w_4265),.q(_w_4266));
  and_bb g1122(.a(n1119),.b(n1121),.q(_w_4874));
  bfr _b_2950(.a(_w_4375),.q(_w_4376));
  bfr _b_4395(.a(_w_5820),.q(_w_5821));
  bfr _b_7299(.a(_w_8724),.q(_w_8725));
  bfr _b_6606(.a(_w_8031),.q(_w_8032));
  bfr _b_2841(.a(_w_4266),.q(_w_4267));
  bfr _b_2205(.a(_w_3630),.q(_w_3631));
  bfr _b_2997(.a(_w_4422),.q(_w_4423));
  spl2 g1247_s_0(.a(n1247),.q0(n1247_0),.q1(n1247_1));
  spl4L G100_s_0(.a(_w_6393),.q0(G100_0),.q1(G100_1),.q2(G100_2),.q3(G100_3));
  bfr _b_4449(.a(_w_5874),.q(_w_5875));
  bfr _b_7066(.a(_w_8491),.q(_w_8492));
  bfr _b_2842(.a(_w_4267),.q(_w_4268));
  bfr _b_6021(.a(_w_7446),.q(_w_7445));
  and_bi g940(.a(G161_8),.b(n939),.q(n940));
  bfr _b_4790(.a(_w_6215),.q(_w_6216));
  bfr _b_3845(.a(_w_5270),.q(_w_5271));
  bfr _b_5234(.a(_w_6659),.q(_w_6660));
  bfr _b_4287(.a(_w_5712),.q(n409_0));
  bfr _b_2846(.a(_w_4271),.q(_w_4272));
  bfr _b_2848(.a(_w_4273),.q(_w_4274));
  bfr _b_5149(.a(_w_6574),.q(_w_6575));
  bfr _b_2101(.a(_w_3526),.q(_w_3527));
  bfr _b_2849(.a(_w_4274),.q(_w_4275));
  bfr _b_4974(.a(_w_6399),.q(_w_6398));
  bfr _b_2851(.a(_w_4276),.q(_w_4277));
  bfr _b_5452(.a(G161),.q(_w_6878));
  bfr _b_4669(.a(_w_6094),.q(_w_6095));
  bfr _b_2852(.a(_w_4277),.q(n1439));
  bfr _b_4652(.a(_w_6077),.q(_w_6078));
  bfr _b_2853(.a(_w_4278),.q(_w_4279));
  and_bb g1372(.a(n1371_0),.b(n346_2),.q(n1372));
  and_bi g1060(.a(G173_8),.b(G5288_1),.q(_w_6012));
  bfr _b_3850(.a(_w_5275),.q(_w_5276));
  bfr _b_4753(.a(_w_6178),.q(_w_6179));
  bfr _b_2855(.a(_w_4280),.q(_w_4281));
  bfr _b_6425(.a(_w_7850),.q(_w_7851));
  bfr _b_2384(.a(_w_3809),.q(_w_3810));
  bfr _b_2856(.a(_w_4281),.q(n1435));
  bfr _b_7417(.a(_w_8842),.q(_w_8843));
  bfr _b_2858(.a(_w_4283),.q(_w_4284));
  bfr _b_6602(.a(_w_8027),.q(_w_8028));
  bfr _b_6232(.a(_w_7657),.q(_w_7658));
  bfr _b_2859(.a(_w_4284),.q(_w_4285));
  bfr _b_3078(.a(_w_4503),.q(_w_4504));
  bfr _b_2860(.a(_w_4285),.q(_w_4286));
  bfr _b_2863(.a(_w_4288),.q(_w_4289));
  bfr _b_6920(.a(_w_8345),.q(_w_8346));
  bfr _b_4995(.a(_w_6420),.q(_w_6421));
  bfr _b_3379(.a(_w_4804),.q(_w_4805));
  bfr _b_2864(.a(_w_4289),.q(G161_6));
  bfr _b_5118(.a(_w_6543),.q(_w_6544));
  bfr _b_2870(.a(_w_4295),.q(_w_4296));
  bfr _b_2872(.a(_w_4297),.q(_w_4298));
  bfr _b_2874(.a(_w_4299),.q(_w_4300));
  bfr _b_7342(.a(_w_8767),.q(_w_8768));
  bfr _b_2877(.a(_w_4302),.q(_w_4303));
  bfr _b_4822(.a(_w_6247),.q(_w_6248));
  and_bb g774(.a(n464_1),.b(n773_0),.q(n774));
  bfr _b_2878(.a(_w_4303),.q(_w_4304));
  bfr _b_2879(.a(_w_4304),.q(n394_2));
  bfr _b_2880(.a(_w_4305),.q(n1338));
  bfr _b_3579(.a(_w_5004),.q(n564));
  bfr _b_2881(.a(_w_4306),.q(G173_20));
  bfr _b_3541(.a(_w_4966),.q(_w_4967));
  bfr _b_2882(.a(_w_4307),.q(_w_4308));
  bfr _b_2738(.a(_w_4163),.q(_w_4164));
  bfr _b_3259(.a(_w_4684),.q(_w_4685));
  bfr _b_5076(.a(_w_6501),.q(_w_6502));
  bfr _b_2883(.a(_w_4308),.q(_w_4309));
  bfr _b_2885(.a(_w_4310),.q(n1321));
  bfr _b_3144(.a(_w_4569),.q(_w_4570));
  bfr _b_3389(.a(_w_4814),.q(_w_4815));
  bfr _b_6234(.a(_w_7659),.q(_w_7660));
  bfr _b_2889(.a(_w_4314),.q(_w_4315));
  bfr _b_3832(.a(_w_5257),.q(n373));
  bfr _b_4431(.a(_w_5856),.q(_w_5857));
  and_bb g680(.a(G176_24),.b(n337_1),.q(n680));
  bfr _b_2890(.a(_w_4315),.q(n1300));
  and_bi g1420(.a(G137_5),.b(n1419),.q(n1420));
  bfr _b_2891(.a(_w_4316),.q(_w_4317));
  bfr _b_4838(.a(_w_6263),.q(_w_6264));
  bfr _b_7509(.a(_w_8934),.q(_w_8935));
  and_bi g1381(.a(G139_5),.b(n1380),.q(n1381));
  bfr _b_2892(.a(_w_4317),.q(_w_4318));
  bfr _b_2895(.a(_w_4320),.q(n1457));
  bfr _b_4617(.a(_w_6042),.q(_w_6043));
  bfr _b_3162(.a(_w_4587),.q(_w_4588));
  bfr _b_6683(.a(_w_8108),.q(_w_8109));
  bfr _b_2896(.a(_w_4321),.q(n472_2));
  bfr _b_2899(.a(_w_4324),.q(_w_4325));
  bfr _b_6398(.a(_w_7823),.q(_w_7824));
  bfr _b_2902(.a(_w_4327),.q(_w_4328));
  bfr _b_1947(.a(_w_3372),.q(n959_2));
  bfr _b_2903(.a(_w_4328),.q(_w_4329));
  bfr _b_5682(.a(_w_7107),.q(_w_7108));
  bfr _b_3530(.a(_w_4955),.q(_w_4956));
  or_bb g1117(.a(n1113),.b(n1116),.q(n1117));
  bfr _b_2905(.a(_w_4330),.q(_w_4331));
  bfr _b_2906(.a(_w_4331),.q(_w_4332));
  bfr _b_2910(.a(_w_4335),.q(G159_0));
  bfr _b_2888(.a(_w_4313),.q(_w_4314));
  bfr _b_2915(.a(_w_4340),.q(_w_4341));
  bfr _b_2143(.a(_w_3568),.q(_w_3569));
  bfr _b_2666(.a(_w_4091),.q(_w_4092));
  bfr _b_2916(.a(_w_4341),.q(_w_4342));
  bfr _b_2947(.a(_w_4372),.q(_w_4373));
  bfr _b_2920(.a(_w_4345),.q(_w_4346));
  bfr _b_2121(.a(_w_3546),.q(_w_3547));
  bfr _b_2921(.a(_w_4346),.q(_w_4347));
  bfr _b_2923(.a(_w_4348),.q(_w_4349));
  bfr _b_3927(.a(_w_5352),.q(_w_5353));
  spl4L G173_s_1(.a(G173_0),.q0(G173_4),.q1(_w_3728),.q2(_w_3729),.q3(G173_7));
  bfr _b_4317(.a(_w_5742),.q(n1192));
  bfr _b_2925(.a(_w_4350),.q(_w_4351));
  bfr _b_2928(.a(_w_4353),.q(n863));
  bfr _b_6034(.a(_w_7459),.q(_w_7460));
  inv inv_G152(.a(G152_0),.q(G5200));
  bfr _b_4339(.a(_w_5764),.q(_w_5765));
  bfr _b_3053(.a(_w_4478),.q(_w_4479));
  bfr _b_4863(.a(_w_6288),.q(G5303));
  bfr _b_6748(.a(_w_8173),.q(_w_8174));
  bfr _b_6216(.a(_w_7641),.q(_w_7642));
  bfr _b_2931(.a(_w_4356),.q(_w_4357));
  bfr _b_2932(.a(_w_4357),.q(_w_4358));
  bfr _b_2074(.a(_w_3499),.q(n443_1));
  bfr _b_2933(.a(_w_4358),.q(_w_4359));
  bfr _b_2937(.a(_w_4362),.q(_w_4363));
  bfr _b_3870(.a(_w_5295),.q(G5212));
  bfr _b_5675(.a(_w_7100),.q(_w_7101));
  bfr _b_2942(.a(_w_4367),.q(n1166));
  bfr _b_2548(.a(_w_3973),.q(G5262));
  bfr _b_2943(.a(_w_4368),.q(_w_4369));
  bfr _b_3083(.a(_w_4508),.q(_w_4509));
  bfr _b_6094(.a(_w_7519),.q(_w_7520));
  bfr _b_3925(.a(_w_5350),.q(_w_5351));
  bfr _b_2944(.a(_w_4369),.q(_w_4370));
  bfr _b_3143(.a(_w_4568),.q(_w_4569));
  bfr _b_3033(.a(_w_4458),.q(_w_4459));
  bfr _b_3153(.a(_w_4578),.q(_w_4579));
  bfr _b_6275(.a(_w_7700),.q(_w_7701));
  bfr _b_2945(.a(_w_4370),.q(_w_4371));
  bfr _b_3210(.a(_w_4635),.q(_w_4636));
  and_bb g1087(.a(n1084),.b(n1086),.q(_w_6115));
  bfr _b_4714(.a(_w_6139),.q(n1128));
  bfr _b_7089(.a(_w_8514),.q(_w_8515));
  bfr _b_2948(.a(_w_4373),.q(n703));
  bfr _b_2951(.a(_w_4376),.q(_w_4377));
  bfr _b_4357(.a(_w_5782),.q(_w_5783));
  bfr _b_4279(.a(_w_5704),.q(_w_5705));
  bfr _b_2952(.a(_w_4377),.q(_w_4378));
  bfr _b_6573(.a(_w_7998),.q(_w_7999));
  bfr _b_2953(.a(_w_4378),.q(_w_4379));
  bfr _b_2957(.a(_w_4382),.q(n448));
  bfr _b_2959(.a(_w_4384),.q(_w_4385));
  bfr _b_3461(.a(_w_4886),.q(_w_4887));
  or_bb g500(.a(n498),.b(n499),.q(_w_4618));
  bfr _b_2961(.a(_w_4386),.q(_w_4387));
  bfr _b_2962(.a(_w_4387),.q(_w_4388));
  bfr _b_7524(.a(_w_8949),.q(_w_8948));
  bfr _b_6056(.a(_w_7481),.q(_w_7482));
  bfr _b_2966(.a(_w_4391),.q(_w_4392));
  bfr _b_5809(.a(_w_7234),.q(_w_7235));
  and_bi g604(.a(n603),.b(n601),.q(n604));
  bfr _b_4712(.a(_w_6137),.q(n379_2));
  spl4L g579_s_0(.a(G5250_0),.q0(_w_6105),.q1(G5250_1),.q2(G5250_2),.q3(G5250_3));
  bfr _b_2967(.a(_w_4392),.q(_w_4393));
  bfr _b_5085(.a(_w_6510),.q(_w_6511));
  bfr _b_2968(.a(_w_4393),.q(_w_4394));
  bfr _b_3558(.a(_w_4983),.q(_w_4984));
  bfr _b_2971(.a(_w_4396),.q(_w_4397));
  and_bb g941(.a(n938),.b(n940),.q(_w_6103));
  and_bb g963(.a(G178),.b(G62),.q(_w_6084));
  bfr _b_2976(.a(_w_4401),.q(_w_4402));
  bfr _b_6704(.a(_w_8129),.q(_w_8130));
  bfr _b_2977(.a(_w_4402),.q(_w_4403));
  bfr _b_2978(.a(_w_4403),.q(_w_4404));
  bfr _b_2980(.a(_w_4405),.q(_w_4406));
  bfr _b_2981(.a(_w_4406),.q(_w_4407));
  bfr _b_7088(.a(_w_8513),.q(_w_8514));
  bfr _b_4041(.a(_w_5466),.q(_w_5467));
  bfr _b_2982(.a(_w_4407),.q(G5268));
  or_bb g1310(.a(n1300_1),.b(n1308_1),.q(n1310));
  bfr _b_2983(.a(_w_4408),.q(_w_4409));
  bfr _b_3587(.a(_w_5012),.q(_w_5013));
  bfr _b_2984(.a(_w_4409),.q(n620));
  bfr _b_5926(.a(_w_7351),.q(_w_7352));
  bfr _b_3429(.a(_w_4854),.q(_w_4855));
  bfr _b_6343(.a(_w_7768),.q(_w_7769));
  bfr _b_4377(.a(_w_5802),.q(_w_5803));
  bfr _b_2986(.a(_w_4411),.q(_w_4412));
  bfr _b_2987(.a(_w_4412),.q(_w_4413));
  bfr _b_4595(.a(_w_6020),.q(n860));
  and_bi g529(.a(n527_1),.b(n524_1),.q(n529));
  bfr _b_2990(.a(_w_4415),.q(_w_4416));
  and_bi g1300(.a(n414_2),.b(n1299),.q(_w_4313));
  bfr _b_2991(.a(_w_4416),.q(G5254_0));
  bfr _b_2992(.a(_w_4417),.q(_w_4418));
  and_bb g805(.a(G80_0),.b(n804_0),.q(n805));
  bfr _b_2994(.a(_w_4419),.q(_w_4420));
  bfr _b_7560(.a(_w_8985),.q(_w_8986));
  bfr _b_2999(.a(_w_4424),.q(_w_4425));
  bfr _b_4506(.a(_w_5931),.q(_w_5932));
  bfr _b_3001(.a(_w_4426),.q(n428_1));
  bfr _b_3003(.a(_w_4428),.q(n578));
  bfr _b_3004(.a(_w_4429),.q(_w_4430));
  bfr _b_3007(.a(_w_4432),.q(_w_4433));
  bfr _b_6271(.a(_w_7696),.q(_w_7697));
  bfr _b_3008(.a(_w_4433),.q(_w_4434));
  bfr _b_6643(.a(_w_8068),.q(_w_8069));
  bfr _b_2765(.a(_w_4190),.q(n387_3));
  bfr _b_3009(.a(_w_4434),.q(_w_4435));
  bfr _b_3010(.a(_w_4435),.q(G5249_0));
  bfr _b_3011(.a(_w_4436),.q(_w_4437));
  bfr _b_3012(.a(_w_4437),.q(n569));
  bfr _b_5309(.a(_w_6734),.q(_w_6735));
  bfr _b_3013(.a(_w_4438),.q(_w_4439));
  bfr _b_3017(.a(_w_4442),.q(_w_4443));
  and_bb g544(.a(n420_1),.b(n425_1),.q(n544));
  bfr _b_3018(.a(_w_4443),.q(n1004));
  and_bb g602(.a(G176_42),.b(n268_1),.q(n602));
  bfr _b_4412(.a(_w_5837),.q(G5291_0));
  bfr _b_3019(.a(_w_4444),.q(_w_4445));
  bfr _b_5833(.a(_w_7258),.q(_w_7259));
  bfr _b_4761(.a(_w_6186),.q(_w_6187));
  bfr _b_3020(.a(_w_4445),.q(_w_4446));
  bfr _b_3021(.a(_w_4446),.q(_w_4447));
  bfr _b_4355(.a(_w_5780),.q(_w_5781));
  bfr _b_4432(.a(_w_5857),.q(_w_5858));
  bfr _b_3022(.a(_w_4447),.q(_w_4448));
  bfr _b_3023(.a(_w_4448),.q(_w_4449));
  bfr _b_3024(.a(_w_4449),.q(_w_4450));
  bfr _b_3025(.a(_w_4450),.q(_w_4451));
  bfr _b_3026(.a(_w_4451),.q(_w_4452));
  bfr _b_4497(.a(_w_5922),.q(n828));
  and_bi g334(.a(G166_12),.b(G107_6),.q(n334));
  bfr _b_4774(.a(_w_6199),.q(_w_6200));
  bfr _b_3028(.a(_w_4453),.q(_w_4454));
  bfr _b_3030(.a(_w_4455),.q(_w_4456));
  bfr _b_3036(.a(_w_4461),.q(n426_2));
  bfr _b_3037(.a(_w_4462),.q(_w_4463));
  bfr _b_2786(.a(_w_4211),.q(_w_4212));
  bfr _b_3038(.a(_w_4463),.q(_w_4464));
  bfr _b_5360(.a(_w_6785),.q(_w_6757));
  spl3L G64_s_5(.a(G64_17),.q0(G64_19),.q1(G64_20),.q2(G64_21));
  bfr _b_3155(.a(_w_4580),.q(_w_4581));
  bfr _b_5254(.a(_w_6679),.q(_w_6680));
  bfr _b_3039(.a(_w_4464),.q(_w_4465));
  and_bb g1158(.a(n1155),.b(n1157),.q(_w_6306));
  bfr _b_3040(.a(_w_4465),.q(n426_3));
  bfr _b_3041(.a(_w_4466),.q(n560));
  bfr _b_3217(.a(_w_4642),.q(G5210));
  bfr _b_2495(.a(_w_3920),.q(_w_3921));
  bfr _b_3070(.a(_w_4495),.q(_w_4496));
  or_bb g1051(.a(n1047),.b(n1050),.q(_w_6223));
  bfr _b_3044(.a(_w_4469),.q(_w_4470));
  bfr _b_3940(.a(_w_5365),.q(_w_5366));
  bfr _b_3045(.a(_w_4470),.q(_w_4471));
  bfr _b_7374(.a(_w_8799),.q(_w_8800));
  bfr _b_3633(.a(_w_5058),.q(_w_5059));
  bfr _b_7482(.a(_w_8907),.q(_w_8875));
  bfr _b_3046(.a(_w_4471),.q(_w_4472));
  and_bb g943(.a(G71_1),.b(n815_5),.q(n943));
  bfr _b_3048(.a(_w_4473),.q(_w_4474));
  bfr _b_5775(.a(_w_7200),.q(_w_7201));
  bfr _b_3681(.a(_w_5106),.q(_w_5107));
  bfr _b_3049(.a(_w_4474),.q(_w_4475));
  bfr _b_3052(.a(_w_4477),.q(_w_4478));
  bfr _b_7344(.a(_w_8769),.q(_w_8770));
  bfr _b_3055(.a(_w_4480),.q(_w_4481));
  bfr _b_3056(.a(_w_4481),.q(_w_4482));
  bfr _b_6544(.a(_w_7969),.q(_w_7970));
  or_bb g820(.a(G173_24),.b(G5257_1),.q(n820));
  bfr _b_3057(.a(_w_4482),.q(_w_4483));
  bfr _b_3058(.a(_w_4483),.q(_w_4484));
  bfr _b_7435(.a(_w_8860),.q(_w_8861));
  bfr _b_4065(.a(_w_5490),.q(_w_5491));
  bfr _b_3063(.a(_w_4488),.q(_w_4489));
  bfr _b_6614(.a(_w_8039),.q(_w_8040));
  bfr _b_3064(.a(_w_4489),.q(_w_4490));
  bfr _b_6780(.a(_w_8205),.q(_w_8206));
  bfr _b_4581(.a(_w_6006),.q(_w_6007));
  bfr _b_4762(.a(_w_6187),.q(n1016));
  bfr _b_3067(.a(_w_4492),.q(_w_4493));
  spl2 g1021_s_1(.a(G5292_3),.q0(G5292_4),.q1(G5292_5));
  bfr _b_3068(.a(_w_4493),.q(_w_4494));
  bfr _b_5232(.a(_w_6657),.q(_w_6658));
  bfr _b_3304(.a(_w_4729),.q(_w_4730));
  bfr _b_7158(.a(_w_8583),.q(_w_8584));
  and_bi g1365(.a(n1363),.b(n1364),.q(n1365));
  bfr _b_3069(.a(_w_4494),.q(_w_4495));
  bfr _b_2491(.a(_w_3916),.q(G144_2));
  bfr _b_3071(.a(_w_4496),.q(_w_4497));
  bfr _b_3072(.a(_w_4497),.q(_w_4498));
  bfr _b_3075(.a(_w_4500),.q(_w_4501));
  bfr _b_7054(.a(_w_8479),.q(_w_8480));
  bfr _b_5075(.a(_w_6500),.q(_w_6501));
  bfr _b_3077(.a(_w_4502),.q(_w_4503));
  bfr _b_3699(.a(_w_5124),.q(_w_5125));
  bfr _b_3081(.a(_w_4506),.q(_w_4507));
  spl2 g716_s_0(.a(n716),.q0(n716_0),.q1(n716_1));
  bfr _b_4606(.a(_w_6031),.q(n871));
  bfr _b_3082(.a(_w_4507),.q(_w_4508));
  bfr _b_3381(.a(_w_4806),.q(_w_4807));
  bfr _b_3394(.a(_w_4819),.q(_w_4820));
  bfr _b_6707(.a(_w_8132),.q(_w_8133));
  bfr _b_5381(.a(_w_6806),.q(_w_6807));
  bfr _b_3846(.a(_w_5271),.q(_w_5272));
  bfr _b_3087(.a(_w_4512),.q(_w_4513));
  spl2 g552_s_5(.a(n552_18),.q0(n552_20),.q1(n552_21));
  bfr _b_3088(.a(_w_4513),.q(_w_4514));
  bfr _b_3983(.a(_w_5408),.q(_w_5409));
  bfr _b_3073(.a(_w_4498),.q(_w_4499));
  bfr _b_3089(.a(_w_4514),.q(i_G151));
  bfr _b_6261(.a(_w_7686),.q(_w_7687));
  bfr _b_3090(.a(_w_4515),.q(_w_4516));
  spl4L G109_s_0(.a(G109),.q0(_w_3511),.q1(G109_1),.q2(G109_2),.q3(_w_3512));
  bfr _b_3093(.a(_w_4518),.q(_w_4519));
  bfr _b_3912(.a(_w_5337),.q(n413));
  and_bi g274(.a(G166_6),.b(G126_6),.q(n274));
  bfr _b_4525(.a(_w_5950),.q(_w_5951));
  bfr _b_3095(.a(_w_4520),.q(_w_4521));
  bfr _b_5287(.a(_w_6712),.q(_w_6713));
  bfr _b_4953(.a(_w_6378),.q(_w_6379));
  bfr _b_3096(.a(_w_4521),.q(_w_4522));
  bfr _b_3097(.a(_w_4522),.q(G176_22));
  bfr _b_6858(.a(_w_8283),.q(_w_8284));
  bfr _b_3098(.a(_w_4523),.q(_w_4524));
  spl2 g1416_s_0(.a(n1416),.q0(n1416_0),.q1(n1416_1));
  bfr _b_3209(.a(_w_4634),.q(_w_4635));
  bfr _b_3099(.a(_w_4524),.q(_w_4525));
  bfr _b_3100(.a(_w_4525),.q(_w_4526));
  bfr _b_3101(.a(_w_4526),.q(_w_4527));
  bfr _b_3244(.a(_w_4669),.q(_w_4670));
  bfr _b_3536(.a(_w_4961),.q(_w_4962));
  bfr _b_3102(.a(_w_4527),.q(_w_4528));
  bfr _b_4778(.a(_w_6203),.q(_w_6204));
  bfr _b_3103(.a(_w_4528),.q(_w_4529));
  bfr _b_3106(.a(_w_4531),.q(_w_4532));
  bfr _b_3107(.a(_w_4532),.q(_w_4533));
  bfr _b_6016(.a(_w_7441),.q(_w_7442));
  bfr _b_4876(.a(_w_6301),.q(n1146));
  bfr _b_3109(.a(_w_4534),.q(_w_4535));
  bfr _b_4653(.a(_w_6078),.q(_w_6079));
  bfr _b_3112(.a(_w_4537),.q(_w_4538));
  bfr _b_6288(.a(_w_7713),.q(_w_7714));
  bfr _b_3967(.a(_w_5392),.q(_w_5393));
  bfr _b_3114(.a(_w_4539),.q(_w_4540));
  bfr _b_3116(.a(_w_4541),.q(_w_4542));
  bfr _b_4234(.a(_w_5659),.q(_w_5660));
  bfr _b_4710(.a(_w_6135),.q(_w_6136));
  bfr _b_4440(.a(_w_5865),.q(G5262_0));
  bfr _b_6342(.a(_w_7767),.q(_w_7768));
  bfr _b_3118(.a(_w_4543),.q(n549));
  bfr _b_4368(.a(_w_5793),.q(_w_5794));
  bfr _b_2272(.a(_w_3697),.q(_w_3698));
  bfr _b_3120(.a(_w_4545),.q(_w_4546));
  spl4L g413_s_0(.a(n413),.q0(n413_0),.q1(_w_5669),.q2(_w_5674),.q3(_w_5679));
  bfr _b_4623(.a(_w_6048),.q(n1465));
  bfr _b_3121(.a(_w_4546),.q(_w_4547));
  bfr _b_3122(.a(_w_4547),.q(G170_0));
  bfr _b_3126(.a(_w_4551),.q(G170_1));
  bfr _b_4133(.a(_w_5558),.q(_w_5559));
  bfr _b_4862(.a(_w_6287),.q(n1068));
  bfr _b_3127(.a(_w_4552),.q(_w_4553));
  and_bi g359(.a(n357),.b(n358),.q(n359));
  bfr _b_3128(.a(_w_4553),.q(G174_0));
  bfr _b_5128(.a(_w_6553),.q(_w_6554));
  bfr _b_3129(.a(_w_4554),.q(_w_4555));
  bfr _b_4567(.a(_w_5992),.q(_w_5993));
  bfr _b_3131(.a(_w_4556),.q(_w_4557));
  bfr _b_3134(.a(_w_4559),.q(_w_4560));
  bfr _b_2763(.a(_w_4188),.q(_w_4189));
  bfr _b_3148(.a(_w_4573),.q(_w_4574));
  bfr _b_3138(.a(_w_4563),.q(_w_4564));
  bfr _b_7180(.a(_w_8605),.q(_w_8606));
  bfr _b_4886(.a(_w_6311),.q(_w_6312));
  bfr _b_5916(.a(_w_7341),.q(_w_7342));
  bfr _b_3135(.a(_w_4560),.q(_w_4561));
  bfr _b_6245(.a(_w_7670),.q(_w_7671));
  bfr _b_3622(.a(_w_5047),.q(_w_5048));
  bfr _b_6136(.a(_w_7561),.q(_w_7529));
  bfr _b_4601(.a(_w_6026),.q(_w_6027));
  and_bi g1411(.a(G135_5),.b(n1410),.q(n1411));
  bfr _b_3137(.a(_w_4562),.q(_w_4563));
  bfr _b_6355(.a(_w_7780),.q(_w_7781));
  bfr _b_3139(.a(_w_4564),.q(_w_4565));
  bfr _b_3140(.a(_w_4565),.q(_w_4566));
  bfr _b_3145(.a(_w_4570),.q(_w_4571));
  bfr _b_6769(.a(_w_8194),.q(_w_8195));
  bfr _b_3149(.a(_w_4574),.q(_w_4575));
  bfr _b_4250(.a(_w_5675),.q(_w_5676));
  bfr _b_4936(.a(_w_6361),.q(_w_6362));
  bfr _b_5933(.a(_w_7358),.q(_w_7359));
  bfr _b_3047(.a(_w_4472),.q(_w_4473));
  bfr _b_3150(.a(_w_4575),.q(_w_4576));
  bfr _b_3151(.a(_w_4576),.q(_w_4577));
  bfr _b_3152(.a(_w_4577),.q(_w_4578));
  bfr _b_2406(.a(_w_3831),.q(_w_3832));
  bfr _b_3154(.a(_w_4579),.q(_w_4580));
  bfr _b_3158(.a(_w_4583),.q(_w_4584));
  bfr _b_4831(.a(_w_6256),.q(_w_6257));
  bfr _b_3159(.a(_w_4584),.q(G5243_0));
  bfr _b_2663(.a(_w_4088),.q(_w_4089));
  bfr _b_3163(.a(_w_4588),.q(_w_4589));
  bfr _b_3264(.a(_w_4689),.q(_w_4690));
  bfr _b_7253(.a(_w_8678),.q(_w_8679));
  and_bi g689(.a(n688),.b(n687),.q(_w_6350));
  bfr _b_3165(.a(_w_4590),.q(_w_4591));
  bfr _b_3619(.a(_w_5044),.q(_w_5045));
  bfr _b_3169(.a(_w_4594),.q(_w_4595));
  bfr _b_3170(.a(_w_4595),.q(_w_4596));
  bfr _b_3472(.a(_w_4897),.q(n347));
  bfr _b_3171(.a(_w_4596),.q(G5261_0));
  bfr _b_4397(.a(_w_5822),.q(_w_5823));
  bfr _b_3172(.a(_w_4597),.q(_w_4598));
  bfr _b_3175(.a(_w_4600),.q(_w_4601));
  bfr _b_5442(.a(_w_6867),.q(_w_6868));
  bfr _b_3176(.a(_w_4601),.q(_w_4602));
  bfr _b_3177(.a(_w_4602),.q(_w_4603));
  bfr _b_3178(.a(_w_4603),.q(_w_4604));
  bfr _b_3180(.a(_w_4605),.q(n243));
  bfr _b_3181(.a(_w_4606),.q(_w_4607));
  bfr _b_3182(.a(_w_4607),.q(n429));
  bfr _b_5186(.a(_w_6611),.q(_w_6612));
  bfr _b_3851(.a(_w_5276),.q(_w_5277));
  bfr _b_7033(.a(_w_8458),.q(_w_8459));
  bfr _b_3183(.a(_w_4608),.q(_w_4609));
  bfr _b_3184(.a(_w_4609),.q(_w_4610));
  bfr _b_5447(.a(_w_6872),.q(_w_6873));
  bfr _b_3185(.a(_w_4610),.q(n515));
  bfr _b_3566(.a(_w_4991),.q(G5257_0));
  bfr _b_3187(.a(_w_4612),.q(_w_4613));
  bfr _b_4987(.a(_w_6412),.q(_w_6411));
  spl2 G83_s_0(.a(_w_8773),.q0(G83_0),.q1(G83_1));
  spl2 g1337_s_0(.a(n1337),.q0(n1337_0),.q1(n1337_1));
  bfr _b_4492(.a(_w_5917),.q(_w_5918));
  bfr _b_3190(.a(_w_4615),.q(_w_4616));
  bfr _b_3795(.a(_w_5220),.q(_w_5221));
  bfr _b_4114(.a(_w_5539),.q(G5195));
  bfr _b_6590(.a(G57),.q(_w_8016));
  bfr _b_3193(.a(_w_4618),.q(_w_4619));
  bfr _b_3194(.a(_w_4619),.q(_w_4620));
  bfr _b_6624(.a(_w_8049),.q(_w_8050));
  bfr _b_3195(.a(_w_4620),.q(n500));
  bfr _b_5586(.a(_w_7011),.q(_w_7012));
  spl2 g449_s_0(.a(n449),.q0(n449_0),.q1(_w_3498));
  and_bi g514(.a(n509_1),.b(n512_1),.q(n514));
  bfr _b_4510(.a(_w_5935),.q(_w_5936));
  bfr _b_5727(.a(_w_7152),.q(_w_7120));
  bfr _b_3200(.a(_w_4625),.q(n542_1));
  bfr _b_3201(.a(_w_4626),.q(_w_4627));
  bfr _b_3204(.a(_w_4629),.q(_w_4630));
  bfr _b_5078(.a(_w_6503),.q(_w_6504));
  bfr _b_3205(.a(_w_4630),.q(n542_2));
  bfr _b_7343(.a(_w_8768),.q(_w_8769));
  spl4L G175_s_3(.a(G175_3),.q0(G175_11),.q1(G175_12),.q2(G175_13),.q3(_w_4655));
  bfr _b_3206(.a(_w_4631),.q(_w_4632));
  bfr _b_3208(.a(_w_4633),.q(n537_5));
  bfr _b_3581(.a(_w_5006),.q(_w_5007));
  bfr _b_3211(.a(_w_4636),.q(n537_6));
  bfr _b_6011(.a(_w_7436),.q(_w_7437));
  bfr _b_5871(.a(_w_7296),.q(_w_7297));
  bfr _b_3212(.a(_w_4637),.q(_w_4638));
  or_bb g1161(.a(n1159),.b(n1160),.q(n1161));
  bfr _b_3218(.a(_w_4643),.q(_w_4644));
  bfr _b_6663(.a(_w_8088),.q(_w_8089));
  bfr _b_5474(.a(_w_6899),.q(_w_6900));
  bfr _b_4421(.a(_w_5846),.q(_w_5847));
  bfr _b_3221(.a(_w_4646),.q(_w_4647));
  bfr _b_6362(.a(_w_7787),.q(_w_7788));
  bfr _b_6269(.a(G43),.q(_w_7695));
  bfr _b_4494(.a(_w_5919),.q(G5264));
  bfr _b_6738(.a(_w_8163),.q(_w_8164));
  bfr _b_3222(.a(_w_4647),.q(n477));
  bfr _b_3223(.a(_w_4648),.q(_w_4649));
  bfr _b_6932(.a(_w_8357),.q(_w_8358));
  bfr _b_3226(.a(_w_4651),.q(_w_4652));
  bfr _b_4562(.a(_w_5987),.q(_w_5988));
  bfr _b_5443(.a(_w_6868),.q(_w_6869));
  bfr _b_3228(.a(_w_4653),.q(_w_4654));
  bfr _b_4063(.a(_w_5488),.q(_w_5489));
  bfr _b_3232(.a(_w_4657),.q(_w_4658));
  bfr _b_5159(.a(_w_6584),.q(_w_6585));
  bfr _b_4184(.a(_w_5609),.q(_w_5610));
  bfr _b_4263(.a(_w_5688),.q(_w_5689));
  bfr _b_3233(.a(_w_4658),.q(_w_4659));
  bfr _b_3234(.a(_w_4659),.q(_w_4660));
  and_bi g511(.a(G94_9),.b(G92_9),.q(n511));
  bfr _b_3236(.a(_w_4661),.q(_w_4662));
  bfr _b_7244(.a(_w_8669),.q(_w_8670));
  bfr _b_3238(.a(_w_4663),.q(_w_4664));
  bfr _b_3240(.a(_w_4665),.q(_w_4666));
  bfr _b_2344(.a(_w_3769),.q(_w_3770));
  bfr _b_4108(.a(_w_5533),.q(_w_5534));
  bfr _b_2188(.a(_w_3613),.q(_w_3614));
  bfr _b_3993(.a(_w_5418),.q(_w_5419));
  bfr _b_3243(.a(_w_4668),.q(_w_4669));
  bfr _b_3248(.a(_w_4673),.q(n456));
  bfr _b_3250(.a(_w_4675),.q(_w_4676));
  bfr _b_3253(.a(_w_4678),.q(G5205));
  bfr _b_3255(.a(_w_4680),.q(n451));
  bfr _b_7142(.a(_w_8567),.q(_w_8568));
  bfr _b_3256(.a(_w_4681),.q(n439));
  bfr _b_3262(.a(_w_4687),.q(_w_4688));
  bfr _b_3263(.a(_w_4688),.q(_w_4689));
  spl2 G26_s_0(.a(_w_7343),.q0(G26_0),.q1(G26_1));
  bfr _b_5019(.a(_w_6444),.q(_w_6445));
  bfr _b_4218(.a(_w_5643),.q(_w_5644));
  bfr _b_3265(.a(_w_4690),.q(_w_4691));
  bfr _b_3266(.a(_w_4691),.q(_w_4692));
  bfr _b_3267(.a(_w_4692),.q(_w_4693));
  bfr _b_6089(.a(_w_7514),.q(_w_7515));
  and_bi g753(.a(n678_1),.b(n574_1),.q(_w_5880));
  bfr _b_4013(.a(_w_5438),.q(_w_5439));
  bfr _b_3268(.a(_w_4693),.q(n289));
  bfr _b_7126(.a(_w_8551),.q(_w_8552));
  bfr _b_3272(.a(_w_4697),.q(_w_4698));
  bfr _b_3274(.a(_w_4699),.q(_w_4700));
  bfr _b_6782(.a(_w_8207),.q(_w_8208));
  spl4L g472_s_1(.a(n472_3),.q0(n472_4),.q1(n472_5),.q2(_w_3982),.q3(_w_3992));
  bfr _b_3370(.a(_w_4795),.q(_w_4796));
  bfr _b_3276(.a(_w_4701),.q(G107_0));
  bfr _b_3277(.a(_w_4702),.q(G107_3));
  bfr _b_3278(.a(_w_4703),.q(n207));
  bfr _b_3280(.a(_w_4705),.q(n557));
  bfr _b_6499(.a(_w_7924),.q(_w_7925));
  bfr _b_3598(.a(_w_5023),.q(_w_5024));
  bfr _b_3281(.a(_w_4706),.q(n636));
  or_bb g420(.a(G144_4),.b(n418_1),.q(n420));
  bfr _b_4969(.a(G101),.q(_w_6394));
  bfr _b_4989(.a(_w_6414),.q(_w_6413));
  bfr _b_3282(.a(_w_4707),.q(n1101));
  bfr _b_3283(.a(_w_4708),.q(G119_0));
  bfr _b_6879(.a(_w_8304),.q(_w_8305));
  bfr _b_3284(.a(_w_4709),.q(_w_4710));
  bfr _b_3288(.a(_w_4713),.q(_w_4714));
  bfr _b_3966(.a(_w_5391),.q(_w_5392));
  bfr _b_3289(.a(_w_4714),.q(_w_4715));
  bfr _b_3766(.a(_w_5191),.q(_w_5192));
  bfr _b_6294(.a(_w_7719),.q(_w_7720));
  spl2 g713_s_0(.a(G5261_0),.q0(_w_3365),.q1(G5261_1));
  spl2 G69_s_0(.a(_w_8296),.q0(G69_0),.q1(G69_1));
  bfr _b_3189(.a(_w_4614),.q(_w_4615));
  bfr _b_3293(.a(_w_4718),.q(_w_4719));
  bfr _b_3294(.a(_w_4719),.q(_w_4720));
  bfr _b_3297(.a(_w_4722),.q(_w_4723));
  or_bb g545(.a(n419_1),.b(n544_0),.q(n545));
  bfr _b_3298(.a(_w_4723),.q(_w_4724));
  bfr _b_3299(.a(_w_4724),.q(G5287));
  bfr _b_7262(.a(_w_8687),.q(_w_8688));
  bfr _b_3300(.a(_w_4725),.q(_w_4726));
  bfr _b_3302(.a(_w_4727),.q(_w_4728));
  spl4L G90_s_3(.a(G90_3),.q0(G90_10),.q1(G90_11),.q2(G90_12),.q3(G90_13));
  spl4L G159_s_0(.a(_w_6786),.q0(_w_4334),.q1(G159_1),.q2(_w_4336),.q3(_w_4338));
  bfr _b_2429(.a(_w_3854),.q(_w_3855));
  bfr _b_3305(.a(_w_4730),.q(_w_4731));
  bfr _b_7183(.a(_w_8608),.q(_w_8609));
  bfr _b_3306(.a(_w_4731),.q(_w_4732));
  bfr _b_3310(.a(_w_4735),.q(_w_4736));
  bfr _b_3311(.a(_w_4736),.q(_w_4737));
  bfr _b_3313(.a(_w_4738),.q(_w_4739));
  or_bb g231(.a(n229),.b(n230),.q(_w_5403));
  bfr _b_3314(.a(_w_4739),.q(_w_4740));
  bfr _b_3315(.a(_w_4740),.q(_w_4741));
  bfr _b_3316(.a(_w_4741),.q(n638));
  bfr _b_6630(.a(_w_8055),.q(_w_8056));
  spl2 g452_s_0(.a(n452),.q0(n452_0),.q1(n452_1));
  bfr _b_3319(.a(_w_4744),.q(n950));
  bfr _b_5806(.a(_w_7231),.q(_w_7232));
  bfr _b_5497(.a(_w_6922),.q(_w_6923));
  bfr _b_3320(.a(_w_4745),.q(_w_4746));
  bfr _b_7164(.a(_w_8589),.q(_w_8590));
  bfr _b_3322(.a(_w_4747),.q(_w_4748));
  bfr _b_3323(.a(_w_4748),.q(_w_4749));
  bfr _b_3324(.a(_w_4749),.q(n462));
  spl2 g497_s_0(.a(n497),.q0(n497_0),.q1(n497_1));
  bfr _b_3325(.a(_w_4750),.q(_w_4751));
  bfr _b_2445(.a(_w_3870),.q(_w_3871));
  bfr _b_3326(.a(_w_4751),.q(_w_4752));
  bfr _b_5822(.a(_w_7247),.q(_w_7248));
  bfr _b_3360(.a(_w_4785),.q(n954));
  bfr _b_3402(.a(_w_4827),.q(_w_4828));
  bfr _b_3330(.a(_w_4755),.q(_w_4756));
  bfr _b_4565(.a(_w_5990),.q(n847));
  bfr _b_3331(.a(_w_4756),.q(_w_4757));
  bfr _b_5850(.a(_w_7275),.q(_w_7276));
  bfr _b_3334(.a(_w_4759),.q(_w_4760));
  and_bi g1318(.a(n1303_2),.b(n1317_0),.q(n1318));
  bfr _b_3337(.a(_w_4762),.q(_w_4763));
  bfr _b_3340(.a(_w_4765),.q(_w_4766));
  bfr _b_3342(.a(_w_4767),.q(_w_4768));
  bfr _b_3343(.a(_w_4768),.q(G5310));
  bfr _b_6674(.a(_w_8099),.q(_w_8100));
  spl2 g1425_s_0(.a(n1425),.q0(n1425_0),.q1(n1425_1));
  bfr _b_3346(.a(_w_4771),.q(_w_4772));
  bfr _b_4253(.a(_w_5678),.q(n413_2));
  bfr _b_5266(.a(_w_6691),.q(_w_6692));
  bfr _b_3349(.a(_w_4774),.q(_w_4775));
  bfr _b_3199(.a(_w_4624),.q(n781));
  bfr _b_4925(.a(_w_6350),.q(_w_6351));
  bfr _b_3287(.a(_w_4712),.q(_w_4713));
  bfr _b_3351(.a(_w_4776),.q(_w_4777));
  bfr _b_3352(.a(_w_4777),.q(_w_4778));
  bfr _b_3953(.a(_w_5378),.q(_w_5379));
  bfr _b_5542(.a(_w_6967),.q(_w_6968));
  bfr _b_2197(.a(_w_3622),.q(_w_3623));
  bfr _b_4399(.a(_w_5824),.q(_w_5825));
  bfr _b_3354(.a(_w_4779),.q(_w_4780));
  bfr _b_6584(.a(_w_8009),.q(_w_8010));
  bfr _b_4200(.a(_w_5625),.q(_w_5626));
  and_bi g742(.a(n722_1),.b(n740_1),.q(n742));
  bfr _b_3356(.a(_w_4781),.q(n327));
  bfr _b_3985(.a(_w_5410),.q(_w_5411));
  bfr _b_3358(.a(_w_4783),.q(n439_2));
  bfr _b_3359(.a(_w_4784),.q(n566));
  bfr _b_3650(.a(_w_5075),.q(_w_5076));
  bfr _b_3363(.a(_w_4788),.q(_w_4789));
  bfr _b_5781(.a(_w_7206),.q(_w_7207));
  bfr _b_3365(.a(_w_4790),.q(_w_4791));
  bfr _b_7165(.a(_w_8590),.q(_w_8591));
  bfr _b_3366(.a(_w_4791),.q(_w_4792));
  bfr _b_4458(.a(_w_5883),.q(n397));
  bfr _b_2857(.a(_w_4282),.q(_w_4283));
  bfr _b_3367(.a(_w_4792),.q(_w_4793));
  bfr _b_3371(.a(_w_4796),.q(_w_4797));
  bfr _b_3935(.a(_w_5360),.q(_w_5361));
  bfr _b_3372(.a(_w_4797),.q(_w_4798));
  or_bb g744(.a(n542_1),.b(n637_1),.q(n744));
  bfr _b_4208(.a(_w_5633),.q(_w_5634));
  bfr _b_3373(.a(_w_4798),.q(_w_4799));
  bfr _b_6893(.a(_w_8318),.q(_w_8319));
  bfr _b_6884(.a(_w_8309),.q(_w_8310));
  bfr _b_3374(.a(_w_4799),.q(_w_4800));
  bfr _b_3621(.a(_w_5046),.q(_w_5047));
  bfr _b_3376(.a(_w_4801),.q(_w_4802));
  bfr _b_3377(.a(_w_4802),.q(_w_4803));
  bfr _b_3378(.a(_w_4803),.q(_w_4804));
  bfr _b_3383(.a(_w_4808),.q(_w_4809));
  spl2 g515_s_0(.a(n515),.q0(n515_0),.q1(n515_1));
  and_bi g1105(.a(G75_0),.b(n802_8),.q(n1105));
  bfr _b_2156(.a(_w_3581),.q(_w_3582));
  bfr _b_3384(.a(_w_4809),.q(_w_4810));
  and_bi g322(.a(G141_0),.b(n321),.q(n322));
  bfr _b_3388(.a(_w_4813),.q(_w_4814));
  bfr _b_3393(.a(_w_4818),.q(_w_4819));
  bfr _b_2998(.a(_w_4423),.q(_w_4424));
  bfr _b_3395(.a(_w_4820),.q(G5231));
  bfr _b_7390(.a(_w_8815),.q(_w_8816));
  bfr _b_4485(.a(_w_5910),.q(_w_5911));
  bfr _b_3396(.a(_w_4821),.q(_w_4822));
  and_bi g283(.a(n281),.b(n282),.q(n283));
  bfr _b_4821(.a(_w_6246),.q(_w_6247));
  bfr _b_4888(.a(_w_6313),.q(_w_6314));
  bfr _b_7191(.a(_w_8616),.q(_w_8617));
  bfr _b_3401(.a(_w_4826),.q(_w_4827));
  or_bb g1244(.a(n1239),.b(n1243),.q(n1244));
  bfr _b_3404(.a(_w_4829),.q(n469));
  bfr _b_5622(.a(_w_7047),.q(_w_7048));
  bfr _b_3505(.a(_w_4930),.q(_w_4931));
  bfr _b_4743(.a(_w_6168),.q(_w_6169));
  bfr _b_3406(.a(_w_4831),.q(_w_4832));
  bfr _b_4389(.a(_w_5814),.q(_w_5815));
  bfr _b_3408(.a(_w_4833),.q(_w_4834));
  bfr _b_3410(.a(_w_4835),.q(_w_4836));
  bfr _b_5797(.a(_w_7222),.q(_w_7223));
  bfr _b_5052(.a(_w_6477),.q(_w_6478));
  bfr _b_3412(.a(_w_4837),.q(_w_4838));
  bfr _b_5879(.a(_w_7304),.q(_w_7305));
  bfr _b_3413(.a(_w_4838),.q(_w_4839));
  bfr _b_3417(.a(_w_4842),.q(_w_4843));
  bfr _b_5331(.a(_w_6756),.q(_w_6736));
  bfr _b_3419(.a(_w_4844),.q(_w_4845));
  bfr _b_4792(.a(_w_6217),.q(_w_6218));
  bfr _b_3420(.a(_w_4845),.q(_w_4846));
  or_bb g491(.a(n489),.b(n490),.q(_w_5584));
  spl2 g1214_s_0(.a(n1214),.q0(n1214_0),.q1(n1214_1));
  bfr _b_4937(.a(_w_6362),.q(_w_6363));
  bfr _b_3423(.a(_w_4848),.q(_w_4849));
  bfr _b_4027(.a(_w_5452),.q(_w_5453));
  bfr _b_3425(.a(_w_4850),.q(_w_4851));
  bfr _b_3431(.a(_w_4856),.q(G145_2));
  bfr _b_2063(.a(_w_3488),.q(G94_0));
  bfr _b_3432(.a(_w_4857),.q(_w_4858));
  spl2 G171_s_0(.a(_w_6961),.q0(_w_3506),.q1(G171_1));
  bfr _b_3433(.a(_w_4858),.q(_w_4859));
  bfr _b_2907(.a(_w_4332),.q(_w_4333));
  bfr _b_3437(.a(_w_4862),.q(G5288_0));
  or_bb g1317(.a(n1315),.b(n1316),.q(n1317));
  bfr _b_3438(.a(_w_4863),.q(_w_4864));
  bfr _b_5637(.a(_w_7062),.q(_w_7063));
  spl2 g710_s_0(.a(n710),.q0(n710_0),.q1(n710_1));
  bfr _b_3439(.a(_w_4864),.q(_w_4865));
  bfr _b_5581(.a(_w_7006),.q(_w_7007));
  bfr _b_3443(.a(_w_4868),.q(_w_4869));
  bfr _b_3444(.a(_w_4869),.q(_w_4870));
  spl3L G113_s_1(.a(G113_3),.q0(G113_4),.q1(G113_5),.q2(_w_3753));
  bfr _b_4877(.a(_w_6302),.q(n1155));
  spl2 g1250_s_0(.a(n1250),.q0(n1250_0),.q1(n1250_1));
  bfr _b_3445(.a(_w_4870),.q(_w_4871));
  bfr _b_5276(.a(_w_6701),.q(_w_6702));
  bfr _b_3471(.a(_w_4896),.q(_w_4897));
  and_bb g1426(.a(n1416_0),.b(n1425_0),.q(n1426));
  bfr _b_4137(.a(_w_5562),.q(_w_5563));
  or_ii g1471(.a(G64_6),.b(n1470),.q(G5314));
  bfr _b_3446(.a(_w_4871),.q(_w_4872));
  bfr _b_5275(.a(_w_6700),.q(_w_6701));
  bfr _b_3447(.a(_w_4872),.q(_w_4873));
  bfr _b_4561(.a(_w_5986),.q(G5269));
  bfr _b_2732(.a(_w_4157),.q(_w_4158));
  bfr _b_3454(.a(_w_4879),.q(_w_4880));
  bfr _b_3462(.a(_w_4887),.q(_w_4888));
  bfr _b_3463(.a(_w_4888),.q(n246));
  bfr _b_4259(.a(_w_5684),.q(_w_5685));
  bfr _b_3465(.a(_w_4890),.q(_w_4891));
  bfr _b_3466(.a(_w_4891),.q(_w_4892));
  and_bb g1396(.a(n1386_0),.b(n1395_0),.q(n1396));
  bfr _b_3546(.a(_w_4971),.q(_w_4972));
  bfr _b_3502(.a(_w_4927),.q(_w_4928));
  bfr _b_4612(.a(_w_6037),.q(_w_6038));
  bfr _b_3468(.a(_w_4893),.q(_w_4894));
  spl4L g570_s_0(.a(G5249_0),.q0(_w_5380),.q1(G5249_1),.q2(G5249_2),.q3(G5249_3));
  bfr _b_3469(.a(_w_4894),.q(_w_4895));
  bfr _b_3470(.a(_w_4895),.q(_w_4896));
  bfr _b_3174(.a(_w_4599),.q(_w_4600));
  bfr _b_3473(.a(_w_4898),.q(_w_4899));
  bfr _b_5355(.a(_w_6780),.q(_w_6781));
  bfr _b_4470(.a(_w_5895),.q(n1407));
  bfr _b_3474(.a(_w_4899),.q(_w_4900));
  bfr _b_6883(.a(_w_8308),.q(_w_8309));
  bfr _b_3599(.a(_w_5024),.q(_w_5025));
  bfr _b_3481(.a(_w_4906),.q(_w_4907));
  bfr _b_4105(.a(_w_5530),.q(_w_5531));
  bfr _b_4430(.a(_w_5855),.q(_w_5856));
  bfr _b_3488(.a(_w_4913),.q(n298));
  bfr _b_3491(.a(_w_4916),.q(_w_4917));
  bfr _b_3492(.a(_w_4917),.q(_w_4918));
  bfr _b_5021(.a(_w_6446),.q(_w_6447));
  and_bb g950(.a(n947),.b(n949),.q(_w_4744));
  or_bb g1204(.a(n1202),.b(n1203),.q(n1204));
  bfr _b_3215(.a(_w_4640),.q(_w_4641));
  bfr _b_4625(.a(_w_6050),.q(n1137));
  bfr _b_3495(.a(_w_4920),.q(n478_1));
  bfr _b_2542(.a(_w_3967),.q(_w_3968));
  bfr _b_3496(.a(_w_4921),.q(_w_4922));
  bfr _b_3497(.a(_w_4922),.q(_w_4923));
  bfr _b_3498(.a(_w_4923),.q(_w_4924));
  bfr _b_4608(.a(_w_6033),.q(_w_6034));
  bfr _b_3500(.a(_w_4925),.q(_w_4926));
  bfr _b_3501(.a(_w_4926),.q(_w_4927));
  bfr _b_2225(.a(_w_3650),.q(G150_2));
  bfr _b_2792(.a(_w_4217),.q(_w_4218));
  bfr _b_3503(.a(_w_4928),.q(_w_4929));
  bfr _b_3510(.a(_w_4935),.q(_w_4936));
  bfr _b_3504(.a(_w_4929),.q(_w_4930));
  and_bi g797(.a(n796),.b(n779_0),.q(_w_5909));
  bfr _b_3506(.a(_w_4931),.q(_w_4932));
  bfr _b_3507(.a(_w_4932),.q(n1334));
  bfr _b_6591(.a(_w_8016),.q(_w_8017));
  bfr _b_3508(.a(_w_4933),.q(_w_4934));
  bfr _b_6815(.a(_w_8240),.q(_w_8241));
  bfr _b_3905(.a(_w_5330),.q(n1277));
  bfr _b_3511(.a(_w_4936),.q(_w_4937));
  spl4L G174_s_4(.a(G174_3),.q0(_w_3736),.q1(_w_3739),.q2(_w_3741),.q3(G174_19));
  bfr _b_4529(.a(_w_5954),.q(_w_5955));
  bfr _b_3512(.a(_w_4937),.q(_w_4938));
  bfr _b_3513(.a(_w_4938),.q(_w_4939));
  bfr _b_7458(.a(_w_8883),.q(_w_8884));
  spl2 G81_s_0(.a(_w_8706),.q0(G81_0),.q1(G81_1));
  bfr _b_3515(.a(_w_4940),.q(_w_4941));
  and_bi g1385(.a(n1384),.b(G139_6),.q(n1385));
  bfr _b_3516(.a(_w_4941),.q(_w_4942));
  bfr _b_3519(.a(_w_4944),.q(G172_6));
  bfr _b_3834(.a(_w_5259),.q(_w_5260));
  bfr _b_3520(.a(_w_4945),.q(n1478));
  bfr _b_5228(.a(_w_6653),.q(_w_6654));
  and_bi g1069(.a(G174_11),.b(G5286_2),.q(n1069));
  bfr _b_3521(.a(_w_4946),.q(_w_4947));
  bfr _b_3522(.a(_w_4947),.q(_w_4948));
  bfr _b_3523(.a(_w_4948),.q(_w_4949));
  bfr _b_3524(.a(_w_4949),.q(_w_4950));
  bfr _b_5457(.a(_w_6882),.q(_w_6883));
  bfr _b_3525(.a(_w_4950),.q(_w_4951));
  and_bi g1077(.a(G174_9),.b(G5287_2),.q(n1077));
  bfr _b_3528(.a(_w_4953),.q(_w_4954));
  bfr _b_5535(.a(_w_6960),.q(_w_6949));
  bfr _b_3531(.a(_w_4956),.q(_w_4957));
  bfr _b_4727(.a(_w_6152),.q(_w_6153));
  bfr _b_3533(.a(_w_4958),.q(_w_4959));
  bfr _b_3534(.a(_w_4959),.q(_w_4960));
  bfr _b_7431(.a(_w_8856),.q(_w_8857));
  bfr _b_2946(.a(_w_4371),.q(n222));
  bfr _b_3538(.a(_w_4963),.q(_w_4964));
  bfr _b_3544(.a(_w_4969),.q(_w_4970));
  bfr _b_5729(.a(_w_7154),.q(_w_7155));
  bfr _b_3545(.a(_w_4970),.q(_w_4971));
  bfr _b_3547(.a(_w_4972),.q(_w_4973));
  bfr _b_6321(.a(_w_7746),.q(_w_7747));
  and_bi g1389(.a(n1387),.b(n1388),.q(n1389));
  bfr _b_3551(.a(_w_4976),.q(n1095));
  bfr _b_3553(.a(_w_4978),.q(G98_5));
  bfr _b_6958(.a(_w_8383),.q(_w_8384));
  bfr _b_2100(.a(_w_3525),.q(_w_3526));
  bfr _b_3556(.a(_w_4981),.q(n201));
  bfr _b_6129(.a(_w_7554),.q(_w_7555));
  bfr _b_2567(.a(_w_3992),.q(_w_3993));
  bfr _b_3166(.a(_w_4591),.q(_w_4592));
  bfr _b_5067(.a(_w_6492),.q(_w_6490));
  bfr _b_3557(.a(_w_4982),.q(_w_4983));
  bfr _b_7199(.a(_w_8624),.q(_w_8625));
  bfr _b_2569(.a(_w_3994),.q(_w_3995));
  bfr _b_3560(.a(_w_4985),.q(_w_4986));
  bfr _b_6916(.a(_w_8341),.q(_w_8342));
  bfr _b_3561(.a(_w_4986),.q(_w_4987));
  bfr _b_5427(.a(_w_6852),.q(_w_6853));
  bfr _b_3220(.a(_w_4645),.q(_w_4646));
  bfr _b_4079(.a(_w_5504),.q(_w_5505));
  bfr _b_3397(.a(_w_4822),.q(n757));
  bfr _b_3562(.a(_w_4987),.q(_w_4988));
  bfr _b_3853(.a(_w_5278),.q(_w_5279));
  bfr _b_3564(.a(_w_4989),.q(_w_4990));
  bfr _b_7167(.a(_w_8592),.q(_w_8593));
  bfr _b_3565(.a(_w_4990),.q(_w_4991));
  bfr _b_3568(.a(_w_4993),.q(_w_4994));
  bfr _b_3743(.a(_w_5168),.q(_w_5169));
  bfr _b_3459(.a(_w_4884),.q(_w_4885));
  bfr _b_3571(.a(_w_4996),.q(_w_4997));
  bfr _b_4896(.a(_w_6321),.q(n1187));
  bfr _b_3572(.a(_w_4997),.q(_w_4998));
  bfr _b_2402(.a(_w_3827),.q(_w_3828));
  bfr _b_3921(.a(_w_5346),.q(_w_5347));
  bfr _b_3573(.a(_w_4998),.q(_w_4999));
  bfr _b_3574(.a(_w_4999),.q(_w_5000));
  and_bb g453(.a(n435_0),.b(n452_0),.q(n453));
  bfr _b_3575(.a(_w_5000),.q(n277));
  bfr _b_1979(.a(_w_3404),.q(G176_28));
  bfr _b_3577(.a(_w_5002),.q(n1449));
  bfr _b_4684(.a(_w_6109),.q(_w_6110));
  bfr _b_3578(.a(_w_5003),.q(G5307));
  bfr _b_3583(.a(_w_5008),.q(_w_5009));
  bfr _b_3585(.a(_w_5010),.q(_w_5011));
  bfr _b_3588(.a(_w_5013),.q(_w_5014));
  and_bb g580(.a(n469_4),.b(n472_2),.q(n580));
  bfr _b_3937(.a(_w_5362),.q(_w_5363));
  bfr _b_3590(.a(_w_5015),.q(_w_5016));
  and_bi g292(.a(n290),.b(n291),.q(n292));
  bfr _b_3591(.a(_w_5016),.q(_w_5017));
  bfr _b_3592(.a(_w_5017),.q(_w_5018));
  bfr _b_5458(.a(_w_6883),.q(_w_6884));
  bfr _b_3593(.a(_w_5018),.q(_w_5019));
  bfr _b_7103(.a(_w_8528),.q(_w_8529));
  spl4L G173_s_4(.a(G173_3),.q0(_w_3722),.q1(_w_3725),.q2(_w_3727),.q3(G173_19));
  bfr _b_3594(.a(_w_5019),.q(_w_5020));
  bfr _b_4426(.a(_w_5851),.q(_w_5852));
  bfr _b_4894(.a(_w_6319),.q(_w_6320));
  bfr _b_7082(.a(_w_8507),.q(_w_8508));
  bfr _b_3597(.a(_w_5022),.q(_w_5023));
  bfr _b_3600(.a(_w_5025),.q(_w_5026));
  bfr _b_3601(.a(_w_5026),.q(_w_5027));
  bfr _b_3604(.a(_w_5029),.q(_w_5030));
  bfr _b_3606(.a(_w_5031),.q(_w_5032));
  bfr _b_3607(.a(_w_5032),.q(_w_5033));
  bfr _b_3609(.a(_w_5034),.q(_w_5035));
  bfr _b_3610(.a(_w_5035),.q(_w_5036));
  bfr _b_3612(.a(_w_5037),.q(n209));
  bfr _b_4391(.a(_w_5816),.q(_w_5817));
  bfr _b_3613(.a(_w_5038),.q(_w_5039));
  spl3L g385_s_0(.a(n385),.q0(n385_0),.q1(n385_1),.q2(n385_2));
  bfr _b_3614(.a(_w_5039),.q(G160_16));
  bfr _b_4376(.a(_w_5801),.q(_w_5802));
  bfr _b_2692(.a(_w_4117),.q(n479_2));
  bfr _b_3615(.a(_w_5040),.q(_w_5041));
  bfr _b_3616(.a(_w_5041),.q(G160_17));
  bfr _b_3617(.a(_w_5042),.q(G160_18));
  bfr _b_6291(.a(_w_7716),.q(_w_7717));
  bfr _b_3624(.a(_w_5049),.q(_w_5050));
  spl4L G123_s_5(.a(G123_19),.q0(G123_20),.q1(G123_21),.q2(G123_22),.q3(G123_23));
  bfr _b_3868(.a(_w_5293),.q(_w_5294));
  bfr _b_4202(.a(_w_5627),.q(n1019));
  bfr _b_4934(.a(_w_6359),.q(_w_6360));
  bfr _b_3625(.a(_w_5050),.q(n257));
  bfr _b_6551(.a(_w_7976),.q(_w_7977));
  bfr _b_4074(.a(_w_5499),.q(_w_5500));
  bfr _b_6050(.a(_w_7475),.q(_w_7476));
  and_bi g1238(.a(n1236),.b(n1237),.q(n1238));
  bfr _b_3627(.a(_w_5052),.q(_w_5053));
  spl2 g678_s_0(.a(n678),.q0(n678_0),.q1(n678_1));
  bfr _b_3628(.a(_w_5053),.q(_w_5054));
  bfr _b_7177(.a(_w_8602),.q(_w_8569));
  bfr _b_3630(.a(_w_5055),.q(_w_5056));
  bfr _b_3636(.a(_w_5061),.q(_w_5062));
  bfr _b_2582(.a(_w_4007),.q(_w_4008));
  bfr _b_3637(.a(_w_5062),.q(n427_1));
  bfr _b_2671(.a(_w_4096),.q(_w_4097));
  bfr _b_3638(.a(_w_5063),.q(_w_5064));
  bfr _b_5112(.a(_w_6537),.q(_w_6535));
  bfr _b_2648(.a(_w_4073),.q(n403_0));
  and_bi g649(.a(n648),.b(n646),.q(n649));
  bfr _b_3641(.a(_w_5066),.q(_w_5067));
  bfr _b_5700(.a(_w_7125),.q(_w_7126));
  or_bb g685(.a(n456_4),.b(n469_6),.q(n685));
  bfr _b_3642(.a(_w_5067),.q(_w_5068));
  bfr _b_2865(.a(_w_4290),.q(_w_4291));
  bfr _b_3643(.a(_w_5068),.q(_w_5069));
  bfr _b_4373(.a(_w_5798),.q(_w_5799));
  bfr _b_3644(.a(_w_5069),.q(_w_5070));
  and_bi g468(.a(G114_0),.b(G123_11),.q(n468));
  bfr _b_3651(.a(_w_5076),.q(_w_5077));
  bfr _b_5795(.a(_w_7220),.q(_w_7221));
  bfr _b_3652(.a(_w_5077),.q(_w_5078));
  bfr _b_3658(.a(_w_5083),.q(_w_5084));
  bfr _b_6509(.a(_w_7934),.q(_w_7935));
  and_ii g1265(.a(n1263_0),.b(n1264),.q(_w_4761));
  bfr _b_3661(.a(_w_5086),.q(_w_5087));
  spl2 G76_s_0(.a(_w_8536),.q0(G76_0),.q1(G76_1));
  bfr _b_3663(.a(_w_5088),.q(_w_5089));
  bfr _b_5350(.a(_w_6775),.q(_w_6776));
  bfr _b_3668(.a(_w_5093),.q(_w_5094));
  and_ii g996(.a(n991),.b(n995),.q(_w_4860));
  bfr _b_3670(.a(_w_5095),.q(_w_5096));
  bfr _b_3751(.a(_w_5176),.q(_w_5177));
  bfr _b_7428(.a(_w_8853),.q(_w_8854));
  bfr _b_6794(.a(_w_8219),.q(_w_8220));
  bfr _b_3671(.a(_w_5096),.q(_w_5097));
  bfr _b_3403(.a(_w_4828),.q(_w_4829));
  or_bb g778(.a(n459_2),.b(n776_1),.q(n778));
  bfr _b_3672(.a(_w_5097),.q(_w_5098));
  spl4L g815_s_0(.a(n815),.q0(n815_0),.q1(n815_1),.q2(n815_2),.q3(n815_3));
  bfr _b_3794(.a(_w_5219),.q(_w_5220));
  bfr _b_6919(.a(_w_8344),.q(_w_8345));
  bfr _b_5576(.a(_w_7001),.q(_w_7002));
  bfr _b_3674(.a(_w_5099),.q(_w_5100));
  bfr _b_3675(.a(_w_5100),.q(_w_5101));
  bfr _b_4210(.a(_w_5635),.q(_w_5636));
  bfr _b_6917(.a(_w_8342),.q(_w_8343));
  bfr _b_4428(.a(_w_5853),.q(_w_5854));
  bfr _b_3677(.a(_w_5102),.q(_w_5103));
  bfr _b_3679(.a(_w_5104),.q(_w_5105));
  bfr _b_3686(.a(_w_5111),.q(_w_5112));
  spl2 G168_s_1(.a(G168_1),.q0(G168_4),.q1(G168_5));
  bfr _b_2762(.a(_w_4187),.q(_w_4188));
  bfr _b_3687(.a(_w_5112),.q(n433));
  and_bb g777(.a(n459_1),.b(n776_0),.q(n777));
  bfr _b_3688(.a(_w_5113),.q(_w_5114));
  bfr _b_5226(.a(_w_6651),.q(_w_6652));
  bfr _b_3691(.a(_w_5116),.q(n565));
  bfr _b_3693(.a(_w_5118),.q(_w_5119));
  spl2 g1395_s_0(.a(n1395),.q0(n1395_0),.q1(n1395_1));
  bfr _b_4476(.a(_w_5901),.q(n794));
  bfr _b_3695(.a(_w_5120),.q(_w_5121));
  bfr _b_3698(.a(_w_5123),.q(_w_5124));
  bfr _b_5868(.a(_w_7293),.q(_w_7294));
  bfr _b_3701(.a(_w_5126),.q(_w_5127));
  bfr _b_3703(.a(_w_5128),.q(_w_5129));
  bfr _b_3704(.a(_w_5129),.q(_w_5130));
  bfr _b_3706(.a(_w_5131),.q(_w_5132));
  bfr _b_3708(.a(_w_5133),.q(_w_5134));
  bfr _b_7449(.a(_w_8874),.q(_w_8841));
  bfr _b_4557(.a(_w_5982),.q(n831));
  and_bi g499(.a(G128_9),.b(G126_9),.q(n499));
  bfr _b_3478(.a(_w_4903),.q(_w_4904));
  bfr _b_3710(.a(_w_5135),.q(_w_5136));
  spl4L G177_s_2(.a(G177_1),.q0(G177_8),.q1(G177_9),.q2(G177_10),.q3(G177_11));
  bfr _b_3711(.a(_w_5136),.q(_w_5137));
  bfr _b_7012(.a(_w_8437),.q(_w_8438));
  bfr _b_4855(.a(_w_6280),.q(_w_6281));
  or_bb g348(.a(G103_0),.b(G169_13),.q(n348));
  bfr _b_5018(.a(G134),.q(_w_6444));
  bfr _b_3712(.a(_w_5137),.q(G5236));
  bfr _b_6877(.a(_w_8302),.q(_w_8303));
  bfr _b_5093(.a(_w_6518),.q(_w_6519));
  bfr _b_3714(.a(_w_5139),.q(_w_5140));
  bfr _b_3715(.a(_w_5140),.q(_w_5141));
  bfr _b_3717(.a(_w_5142),.q(_w_5143));
  bfr _b_7189(.a(_w_8614),.q(_w_8615));
  bfr _b_6838(.a(_w_8263),.q(_w_8264));
  bfr _b_4337(.a(_w_5762),.q(_w_5763));
  bfr _b_5762(.a(_w_7187),.q(_w_7188));
  bfr _b_3722(.a(_w_5147),.q(G160_0));
  bfr _b_3727(.a(_w_5152),.q(G5232));
  bfr _b_3731(.a(_w_5156),.q(_w_5157));
  spl4L G176_s_3(.a(G176_2),.q0(G176_12),.q1(_w_3405),.q2(_w_3409),.q3(G176_15));
  bfr _b_3732(.a(_w_5157),.q(_w_5158));
  and_bi g219(.a(G145_0),.b(n218),.q(n219));
  spl4L g185_s_0(.a(G5221_0),.q0(_w_5159),.q1(G5221_1),.q2(G5221_2),.q3(G5221_3));
  bfr _b_3733(.a(_w_5158),.q(n722));
  bfr _b_3734(.a(_w_5159),.q(_w_5160));
  bfr _b_4264(.a(_w_5689),.q(_w_5690));
  bfr _b_3735(.a(_w_5160),.q(_w_5161));
  bfr _b_2299(.a(_w_3724),.q(G173_16));
  bfr _b_4171(.a(_w_5596),.q(_w_5597));
  bfr _b_6390(.a(_w_7815),.q(_w_7816));
  bfr _b_3602(.a(_w_5027),.q(_w_5028));
  bfr _b_3736(.a(_w_5161),.q(_w_5162));
  bfr _b_5601(.a(_w_7026),.q(_w_7027));
  bfr _b_4614(.a(_w_6039),.q(_w_6040));
  bfr _b_3740(.a(_w_5165),.q(_w_5166));
  or_bb g1326(.a(n1312),.b(n1325),.q(n1326));
  bfr _b_4721(.a(_w_6146),.q(_w_6147));
  bfr _b_3742(.a(_w_5167),.q(_w_5168));
  bfr _b_3745(.a(_w_5170),.q(_w_5171));
  and_bb g548(.a(n408_1),.b(n547_0),.q(n548));
  bfr _b_4300(.a(_w_5725),.q(n409_1));
  bfr _b_3746(.a(_w_5171),.q(_w_5172));
  bfr _b_3747(.a(_w_5172),.q(_w_5173));
  bfr _b_3750(.a(_w_5175),.q(_w_5176));
  bfr _b_3752(.a(_w_5177),.q(_w_5178));
  bfr _b_3755(.a(_w_5180),.q(_w_5181));
  bfr _b_3758(.a(_w_5183),.q(_w_5184));
  bfr _b_3759(.a(_w_5184),.q(_w_5185));
  bfr _b_3899(.a(_w_5324),.q(_w_5325));
  bfr _b_3760(.a(_w_5185),.q(_w_5186));
  bfr _b_4197(.a(_w_5622),.q(_w_5623));
  bfr _b_3761(.a(_w_5186),.q(_w_5187));
  bfr _b_3161(.a(_w_4586),.q(_w_4587));
  bfr _b_5058(.a(_w_6483),.q(_w_6481));
  bfr _b_3664(.a(_w_5089),.q(_w_5090));
  bfr _b_3762(.a(_w_5187),.q(_w_5188));
  bfr _b_4267(.a(_w_5692),.q(G156_1));
  bfr _b_3768(.a(_w_5193),.q(_w_5194));
  bfr _b_3770(.a(_w_5195),.q(G5221));
  bfr _b_3771(.a(_w_5196),.q(_w_5197));
  bfr _b_3775(.a(_w_5200),.q(_w_5201));
  bfr _b_3773(.a(_w_5198),.q(_w_5199));
  bfr _b_3776(.a(_w_5201),.q(_w_5202));
  bfr _b_7384(.a(_w_8809),.q(_w_8810));
  bfr _b_2414(.a(_w_3839),.q(_w_3840));
  bfr _b_3780(.a(_w_5205),.q(_w_5206));
  bfr _b_4056(.a(_w_5481),.q(n218));
  bfr _b_3781(.a(_w_5206),.q(_w_5207));
  and_bi g574(.a(n573),.b(n572_0),.q(_w_4663));
  bfr _b_3157(.a(_w_4582),.q(_w_4583));
  bfr _b_3782(.a(_w_5207),.q(_w_5208));
  bfr _b_3785(.a(_w_5210),.q(_w_5211));
  bfr _b_2629(.a(_w_4054),.q(_w_4055));
  bfr _b_3787(.a(_w_5212),.q(_w_5213));
  bfr _b_1965(.a(_w_3390),.q(_w_3391));
  bfr _b_2733(.a(_w_4158),.q(_w_4159));
  bfr _b_4232(.a(_w_5657),.q(_w_5658));
  bfr _b_2901(.a(_w_4326),.q(_w_4327));
  bfr _b_4591(.a(_w_6016),.q(_w_6017));
  bfr _b_5910(.a(_w_7335),.q(_w_7336));
  or_bb g1350(.a(n1345),.b(n1349),.q(n1350));
  bfr _b_3788(.a(_w_5213),.q(_w_5214));
  and_bi g821(.a(G173_23),.b(G5253_1),.q(n821));
  bfr _b_3792(.a(_w_5217),.q(_w_5218));
  bfr _b_3623(.a(_w_5048),.q(_w_5049));
  bfr _b_3798(.a(_w_5223),.q(_w_5224));
  bfr _b_3799(.a(_w_5224),.q(_w_5225));
  bfr _b_3085(.a(_w_4510),.q(_w_4511));
  bfr _b_3800(.a(_w_5225),.q(_w_5226));
  bfr _b_3801(.a(_w_5226),.q(_w_5227));
  bfr _b_5842(.a(_w_7267),.q(_w_7268));
  spl4L G117_s_0(.a(_w_6417),.q0(G117_0),.q1(G117_1),.q2(G117_2),.q3(G117_3));
  bfr _b_3802(.a(_w_5227),.q(_w_5228));
  bfr _b_5882(.a(_w_7307),.q(_w_7308));
  spl2 G94_s_1(.a(G94_1),.q0(G94_4),.q1(G94_5));
  bfr _b_4020(.a(_w_5445),.q(_w_5446));
  bfr _b_4360(.a(_w_5785),.q(_w_5786));
  bfr _b_3804(.a(_w_5229),.q(_w_5230));
  and_bb g1196(.a(n1192_0),.b(n1195_0),.q(n1196));
  bfr _b_3810(.a(_w_5235),.q(_w_5236));
  bfr _b_3811(.a(_w_5236),.q(_w_5237));
  bfr _b_5403(.a(_w_6828),.q(_w_6829));
  bfr _b_4134(.a(_w_5559),.q(_w_5560));
  bfr _b_3812(.a(_w_5237),.q(_w_5238));
  bfr _b_6087(.a(_w_7512),.q(_w_7513));
  bfr _b_2200(.a(_w_3625),.q(_w_3626));
  bfr _b_3813(.a(_w_5238),.q(_w_5239));
  bfr _b_2974(.a(_w_4399),.q(n629));
  bfr _b_2358(.a(_w_3783),.q(_w_3784));
  bfr _b_3816(.a(_w_5241),.q(_w_5242));
  bfr _b_2355(.a(_w_3780),.q(_w_3781));
  bfr _b_3817(.a(_w_5242),.q(_w_5243));
  bfr _b_5928(.a(_w_7353),.q(_w_7354));
  or_bb g890(.a(n888),.b(n889),.q(n890));
  bfr _b_3818(.a(_w_5243),.q(_w_5244));
  bfr _b_3821(.a(_w_5246),.q(_w_5247));
  bfr _b_5981(.a(_w_7406),.q(_w_7407));
  bfr _b_3823(.a(_w_5248),.q(_w_5249));
  bfr _b_3825(.a(_w_5250),.q(_w_5251));
  or_bb g960(.a(G170_1),.b(n959_0),.q(n960));
  bfr _b_3826(.a(_w_5251),.q(G130_1));
  bfr _b_5070(.a(_w_6495),.q(_w_6496));
  bfr _b_3640(.a(_w_5065),.q(_w_5066));
  bfr _b_3833(.a(_w_5258),.q(_w_5259));
  bfr _b_3835(.a(_w_5260),.q(_w_5261));
  bfr _b_4059(.a(_w_5484),.q(G109_7));
  bfr _b_5313(.a(_w_6738),.q(_w_6739));
  bfr _b_5255(.a(_w_6680),.q(_w_6681));
  and_bi g349(.a(G103_4),.b(G168_12),.q(n349));
  bfr _b_4487(.a(_w_5912),.q(_w_5913));
  bfr _b_6901(.a(_w_8326),.q(_w_8327));
  bfr _b_4304(.a(_w_5729),.q(_w_5730));
  bfr _b_3836(.a(_w_5261),.q(_w_5262));
  bfr _b_4679(.a(_w_6104),.q(G107_7));
  bfr _b_2066(.a(_w_3491),.q(_w_3492));
  and_bi g930(.a(G160_21),.b(G5249_5),.q(n930));
  bfr _b_3839(.a(_w_5264),.q(_w_5265));
  bfr _b_7330(.a(_w_8755),.q(_w_8756));
  bfr _b_3840(.a(_w_5265),.q(_w_5266));
  bfr _b_7375(.a(_w_8800),.q(_w_8801));
  spl2 g769_s_0(.a(n769),.q0(n769_0),.q1(n769_1));
  bfr _b_3779(.a(_w_5204),.q(_w_5205));
  bfr _b_3842(.a(_w_5267),.q(_w_5268));
  bfr _b_3844(.a(_w_5269),.q(_w_5270));
  bfr _b_3847(.a(_w_5272),.q(_w_5273));
  bfr _b_3854(.a(_w_5279),.q(_w_5280));
  bfr _b_3855(.a(_w_5280),.q(_w_5281));
  bfr _b_3856(.a(_w_5281),.q(_w_5282));
  bfr _b_4346(.a(_w_5771),.q(_w_5772));
  or_bb g1187(.a(n1185),.b(n1186),.q(_w_6318));
  bfr _b_4593(.a(_w_6018),.q(_w_6019));
  bfr _b_4836(.a(_w_6261),.q(_w_6262));
  bfr _b_5089(.a(_w_6514),.q(_w_6515));
  bfr _b_3859(.a(_w_5284),.q(_w_5285));
  bfr _b_4848(.a(_w_6273),.q(_w_6274));
  bfr _b_3863(.a(_w_5288),.q(_w_5289));
  bfr _b_3864(.a(_w_5289),.q(_w_5290));
  spl2 g746_s_0(.a(n746),.q0(n746_0),.q1(n746_1));
  bfr _b_3867(.a(_w_5292),.q(_w_5293));
  bfr _b_4434(.a(_w_5859),.q(_w_5860));
  bfr _b_3871(.a(_w_5296),.q(n731));
  bfr _b_2506(.a(_w_3931),.q(G123_10));
  bfr _b_3873(.a(_w_5298),.q(_w_5299));
  bfr _b_7204(.a(_w_8629),.q(_w_8630));
  bfr _b_3880(.a(_w_5305),.q(_w_5306));
  bfr _b_5062(.a(G138),.q(_w_6488));
  bfr _b_6134(.a(_w_7559),.q(_w_7560));
  and_bi g865(.a(G6_1),.b(n632_4),.q(n865));
  bfr _b_4016(.a(_w_5441),.q(n614));
  bfr _b_4660(.a(_w_6085),.q(_w_6086));
  bfr _b_3881(.a(_w_5306),.q(_w_5307));
  bfr _b_3882(.a(_w_5307),.q(_w_5308));
  bfr _b_7184(.a(_w_8609),.q(_w_8610));
  bfr _b_3885(.a(_w_5310),.q(_w_5311));
  and_bi g1415(.a(n1414),.b(G135_6),.q(n1415));
  bfr _b_2979(.a(_w_4404),.q(n398_1));
  bfr _b_2700(.a(_w_4125),.q(n407_1));
  bfr _b_3886(.a(_w_5311),.q(_w_5312));
  bfr _b_4940(.a(_w_6365),.q(_w_6366));
  or_bb g299(.a(G169_9),.b(G92_0),.q(n299));
  bfr _b_3887(.a(_w_5312),.q(_w_5313));
  bfr _b_6242(.a(_w_7667),.q(_w_7668));
  bfr _b_3892(.a(_w_5317),.q(_w_5318));
  bfr _b_3895(.a(_w_5320),.q(_w_5321));
  bfr _b_2054(.a(_w_3479),.q(_w_3480));
  bfr _b_3900(.a(_w_5325),.q(_w_5326));
  bfr _b_2295(.a(_w_3720),.q(_w_3721));
  bfr _b_2461(.a(_w_3886),.q(_w_3887));
  bfr _b_3901(.a(_w_5326),.q(_w_5327));
  bfr _b_3902(.a(_w_5327),.q(_w_5328));
  bfr _b_5527(.a(_w_6952),.q(_w_6953));
  bfr _b_3907(.a(_w_5332),.q(_w_5333));
  bfr _b_3908(.a(_w_5333),.q(_w_5334));
  bfr _b_3909(.a(_w_5334),.q(n289_1));
  bfr _b_5181(.a(_w_6606),.q(_w_6607));
  bfr _b_4382(.a(_w_5807),.q(_w_5808));
  bfr _b_2850(.a(_w_4275),.q(_w_4276));
  bfr _b_3910(.a(_w_5335),.q(_w_5336));
  spl4L G96_s_3(.a(G96_3),.q0(G96_10),.q1(G96_11),.q2(G96_12),.q3(G96_13));
  bfr _b_3130(.a(_w_4555),.q(G174_1));
  bfr _b_4502(.a(_w_5927),.q(_w_5928));
  bfr _b_3911(.a(_w_5336),.q(n673));
  bfr _b_6406(.a(_w_7831),.q(_w_7832));
  bfr _b_3173(.a(_w_4598),.q(_w_4599));
  bfr _b_3913(.a(_w_5338),.q(G96_0));
  bfr _b_3914(.a(_w_5339),.q(G96_3));
  bfr _b_3915(.a(_w_5340),.q(_w_5341));
  and_bi g642(.a(n375_4),.b(n640_1),.q(n642));
  bfr _b_2667(.a(_w_4092),.q(n256_1));
  bfr _b_4604(.a(_w_6029),.q(_w_6030));
  bfr _b_3917(.a(_w_5342),.q(_w_5343));
  bfr _b_7526(.a(_w_8951),.q(_w_8950));
  bfr _b_5177(.a(G152),.q(_w_6603));
  bfr _b_4364(.a(_w_5789),.q(_w_5790));
  bfr _b_4540(.a(_w_5965),.q(_w_5966));
  bfr _b_3918(.a(_w_5343),.q(_w_5344));
  bfr _b_3922(.a(_w_5347),.q(_w_5348));
  bfr _b_3923(.a(_w_5348),.q(_w_5349));
  bfr _b_3924(.a(_w_5349),.q(_w_5350));
  bfr _b_3928(.a(_w_5353),.q(_w_5354));
  bfr _b_3930(.a(_w_5355),.q(_w_5356));
  bfr _b_5195(.a(_w_6620),.q(_w_6621));
  bfr _b_3932(.a(_w_5357),.q(_w_5358));
  spl2 g1164_s_0(.a(n1164),.q0(n1164_0),.q1(n1164_1));
  bfr _b_4107(.a(_w_5532),.q(_w_5533));
  bfr _b_7439(.a(_w_8864),.q(_w_8865));
  bfr _b_4471(.a(_w_5896),.q(G128_3));
  bfr _b_7053(.a(_w_8478),.q(_w_8479));
  bfr _b_4545(.a(_w_5970),.q(_w_5971));
  bfr _b_2727(.a(_w_4152),.q(_w_4153));
  bfr _b_3933(.a(_w_5358),.q(_w_5359));
  bfr _b_3939(.a(_w_5364),.q(_w_5365));
  spl2 g393_s_0(.a(n393),.q0(n393_0),.q1(_w_3513));
  bfr _b_4576(.a(_w_6001),.q(_w_6002));
  bfr _b_3941(.a(_w_5366),.q(_w_5367));
  bfr _b_3942(.a(_w_5367),.q(_w_5368));
  bfr _b_3946(.a(_w_5371),.q(_w_5372));
  bfr _b_2658(.a(_w_4083),.q(_w_4084));
  bfr _b_5074(.a(_w_6499),.q(_w_6500));
  bfr _b_3944(.a(_w_5369),.q(_w_5370));
  bfr _b_3947(.a(_w_5372),.q(_w_5373));
  bfr _b_6012(.a(_w_7437),.q(_w_7438));
  bfr _b_3949(.a(_w_5374),.q(_w_5375));
  bfr _b_3950(.a(_w_5375),.q(G129_1));
  bfr _b_7287(.a(_w_8712),.q(_w_8713));
  bfr _b_3952(.a(_w_5377),.q(_w_5378));
  bfr _b_4816(.a(_w_6241),.q(_w_6242));
  or_bb g338(.a(G101_8),.b(G88_0),.q(n338));
  bfr _b_3954(.a(_w_5379),.q(G5271));
  bfr _b_6032(.a(_w_7457),.q(_w_7456));
  bfr _b_4403(.a(_w_5828),.q(n471));
  bfr _b_3955(.a(_w_5380),.q(_w_5381));
  bfr _b_3957(.a(_w_5382),.q(_w_5383));
  bfr _b_4806(.a(_w_6231),.q(_w_6232));
  bfr _b_3958(.a(_w_5383),.q(_w_5384));
  spl2 g409_s_1(.a(n409_3),.q0(n409_4),.q1(n409_5));
  bfr _b_3959(.a(_w_5384),.q(_w_5385));
  or_bb g1469(.a(n1467),.b(n1468),.q(_w_4255));
  and_bb g342(.a(G88_2),.b(G98_7),.q(n342));
  bfr _b_3963(.a(_w_5388),.q(_w_5389));
  bfr _b_3214(.a(_w_4639),.q(_w_4640));
  bfr _b_4950(.a(_w_6375),.q(_w_6376));
  bfr _b_4149(.a(_w_5574),.q(_w_5575));
  bfr _b_3969(.a(_w_5394),.q(_w_5395));
  bfr _b_3970(.a(_w_5395),.q(n710));
  and_bb g1160(.a(G83_1),.b(n815_10),.q(n1160));
  bfr _b_3971(.a(_w_5396),.q(_w_5397));
  bfr _b_3972(.a(_w_5397),.q(_w_5398));
  bfr _b_6395(.a(_w_7820),.q(_w_7799));
  bfr _b_3975(.a(_w_5400),.q(_w_5401));
  bfr _b_4394(.a(_w_5819),.q(_w_5820));
  bfr _b_3979(.a(_w_5404),.q(_w_5405));
  bfr _b_5066(.a(_w_6491),.q(_w_6492));
  bfr _b_3980(.a(_w_5405),.q(_w_5406));
  bfr _b_6154(.a(_w_7579),.q(_w_7580));
  bfr _b_3981(.a(_w_5406),.q(n231));
  bfr _b_7070(.a(_w_8495),.q(_w_8496));
  bfr _b_3982(.a(_w_5407),.q(n374_0));
  bfr _b_3987(.a(_w_5412),.q(_w_5413));
  bfr _b_6515(.a(_w_7940),.q(_w_7941));
  bfr _b_3992(.a(_w_5417),.q(_w_5418));
  bfr _b_4829(.a(_w_6254),.q(_w_6255));
  bfr _b_5040(.a(_w_6465),.q(_w_6466));
  bfr _b_3995(.a(_w_5420),.q(_w_5421));
  bfr _b_3996(.a(_w_5421),.q(_w_5422));
  bfr _b_3997(.a(_w_5422),.q(_w_5423));
  bfr _b_4651(.a(_w_6076),.q(_w_6077));
  bfr _b_4001(.a(_w_5426),.q(_w_5427));
  bfr _b_5908(.a(_w_7333),.q(_w_7334));
  bfr _b_4005(.a(_w_5430),.q(_w_5431));
  bfr _b_4011(.a(_w_5436),.q(_w_5437));
  bfr _b_4014(.a(_w_5439),.q(n1303_1));
  bfr _b_3416(.a(_w_4841),.q(n1446));
  bfr _b_2936(.a(_w_4361),.q(_w_4362));
  bfr _b_4019(.a(_w_5444),.q(_w_5445));
  bfr _b_2050(.a(_w_3475),.q(n462_2));
  bfr _b_4021(.a(_w_5446),.q(_w_5447));
  bfr _b_4026(.a(_w_5451),.q(_w_5452));
  bfr _b_7424(.a(_w_8849),.q(_w_8850));
  bfr _b_5498(.a(_w_6923),.q(_w_6924));
  bfr _b_4028(.a(_w_5453),.q(_w_5454));
  bfr _b_4029(.a(_w_5454),.q(G5252));
  bfr _b_3477(.a(_w_4902),.q(n994));
  bfr _b_4030(.a(_w_5455),.q(n390));
  bfr _b_4472(.a(_w_5897),.q(n1182));
  bfr _b_4386(.a(_w_5811),.q(_w_5812));
  bfr _b_2845(.a(_w_4270),.q(_w_4271));
  bfr _b_4032(.a(_w_5457),.q(_w_5458));
  spl4L G92_s_0(.a(G92),.q0(_w_3944),.q1(G92_1),.q2(G92_2),.q3(_w_3945));
  bfr _b_4033(.a(_w_5458),.q(_w_5459));
  bfr _b_4034(.a(_w_5459),.q(G5267));
  and_bb g578(.a(n575),.b(n577),.q(_w_4427));
  bfr _b_2254(.a(_w_3679),.q(_w_3680));
  bfr _b_4036(.a(_w_5461),.q(_w_5462));
  bfr _b_4037(.a(_w_5462),.q(n478));
  bfr _b_4038(.a(_w_5463),.q(G174_5));
  bfr _b_7205(.a(_w_8630),.q(_w_8631));
  bfr _b_4043(.a(_w_5468),.q(_w_5469));
  and_bb g1287(.a(n1268_2),.b(n375_6),.q(n1287));
  bfr _b_4843(.a(_w_6268),.q(_w_6269));
  and_bb g1450(.a(n1445),.b(n1449),.q(n1450));
  bfr _b_4044(.a(_w_5469),.q(G5215));
  bfr _b_2911(.a(_w_4336),.q(_w_4337));
  bfr _b_4047(.a(_w_5472),.q(n434));
  bfr _b_4048(.a(_w_5473),.q(_w_5474));
  bfr _b_5013(.a(G131),.q(_w_6439));
  bfr _b_4051(.a(_w_5476),.q(n211));
  bfr _b_6302(.a(_w_7727),.q(_w_7728));
  bfr _b_3031(.a(_w_4456),.q(_w_4457));
  bfr _b_4055(.a(_w_5480),.q(_w_5481));
  bfr _b_4058(.a(_w_5483),.q(n603));
  bfr _b_4070(.a(_w_5495),.q(G177_0));
  bfr _b_4075(.a(_w_5500),.q(G177_1));
  bfr _b_6174(.a(_w_7599),.q(_w_7600));
  bfr _b_3292(.a(_w_4717),.q(_w_4718));
  bfr _b_5025(.a(_w_6450),.q(_w_6451));
  bfr _b_4076(.a(_w_5501),.q(G177_2));
  bfr _b_4077(.a(_w_5502),.q(_w_5503));
  bfr _b_4081(.a(_w_5506),.q(_w_5507));
  bfr _b_4082(.a(_w_5507),.q(_w_5508));
  bfr _b_3976(.a(_w_5401),.q(_w_5402));
  bfr _b_5033(.a(_w_6458),.q(_w_6459));
  bfr _b_4084(.a(_w_5509),.q(_w_5510));
  bfr _b_4086(.a(_w_5511),.q(_w_5512));
  bfr _b_4087(.a(_w_5512),.q(_w_5513));
  bfr _b_4349(.a(_w_5774),.q(_w_5775));
  bfr _b_4089(.a(_w_5514),.q(_w_5515));
  bfr _b_4090(.a(_w_5515),.q(_w_5516));
  bfr _b_4093(.a(_w_5518),.q(_w_5519));
  bfr _b_4096(.a(_w_5521),.q(_w_5522));
  and_bi g1029(.a(G174_13),.b(G5285_1),.q(n1029));
  bfr _b_4097(.a(_w_5522),.q(_w_5523));
  bfr _b_4099(.a(_w_5524),.q(_w_5525));
  spl4L G98_s_3(.a(G98_2),.q0(G98_12),.q1(G98_13),.q2(G98_14),.q3(G98_15));
  bfr _b_4102(.a(_w_5527),.q(_w_5528));
  bfr _b_4103(.a(_w_5528),.q(_w_5529));
  bfr _b_4104(.a(_w_5529),.q(_w_5530));
  bfr _b_4112(.a(_w_5537),.q(_w_5538));
  bfr _b_3830(.a(_w_5255),.q(n268_1));
  bfr _b_3241(.a(_w_4666),.q(n574));
  bfr _b_4117(.a(_w_5542),.q(_w_5543));
  bfr _b_2142(.a(_w_3567),.q(_w_3568));
  bfr _b_4118(.a(_w_5543),.q(_w_5544));
  bfr _b_5301(.a(_w_6726),.q(_w_6727));
  bfr _b_4119(.a(_w_5544),.q(_w_5545));
  bfr _b_7219(.a(_w_8644),.q(_w_8645));
  bfr _b_3778(.a(_w_5203),.q(_w_5204));
  bfr _b_4122(.a(_w_5547),.q(_w_5548));
  and_bi g317(.a(n316),.b(G135_1),.q(n317));
  bfr _b_5042(.a(_w_6467),.q(_w_6468));
  spl2 G127_s_0(.a(_w_6433),.q0(G127_0),.q1(_w_4026));
  bfr _b_2964(.a(_w_4389),.q(_w_4390));
  bfr _b_4125(.a(_w_5550),.q(_w_5551));
  bfr _b_6000(.a(_w_7425),.q(_w_7426));
  and_bi g1047(.a(n1046),.b(n1044),.q(_w_6052));
  bfr _b_4129(.a(_w_5554),.q(_w_5555));
  bfr _b_4931(.a(_w_6356),.q(_w_6357));
  bfr _b_4131(.a(_w_5556),.q(_w_5557));
  bfr _b_4132(.a(_w_5557),.q(_w_5558));
  bfr _b_4138(.a(_w_5563),.q(_w_5564));
  or_bb g1147(.a(G160_9),.b(G5291_5),.q(n1147));
  bfr _b_4142(.a(_w_5567),.q(_w_5568));
  and_bb g333(.a(G107_5),.b(G167_11),.q(n333));
  bfr _b_4143(.a(_w_5568),.q(_w_5569));
  bfr _b_4144(.a(_w_5569),.q(_w_5570));
  bfr _b_4145(.a(_w_5570),.q(_w_5571));
  bfr _b_3986(.a(_w_5411),.q(_w_5412));
  bfr _b_4147(.a(_w_5572),.q(_w_5573));
  bfr _b_4151(.a(_w_5576),.q(_w_5577));
  bfr _b_4785(.a(_w_6210),.q(G5294));
  bfr _b_4152(.a(_w_5577),.q(G5211));
  bfr _b_4154(.a(_w_5579),.q(_w_5580));
  bfr _b_4587(.a(_w_6012),.q(n1060));
  bfr _b_4155(.a(_w_5580),.q(_w_5581));
  bfr _b_5236(.a(_w_6661),.q(_w_6662));
  bfr _b_4157(.a(_w_5582),.q(_w_5583));
  bfr _b_4158(.a(_w_5583),.q(n224_1));
  bfr _b_4160(.a(_w_5585),.q(n1055));
  bfr _b_4416(.a(_w_5841),.q(_w_5842));
  bfr _b_4162(.a(_w_5587),.q(_w_5588));
  spl2 g374_s_0(.a(n374),.q0(_w_5407),.q1(n374_1));
  bfr _b_4163(.a(_w_5588),.q(_w_5589));
  bfr _b_4283(.a(_w_5708),.q(_w_5709));
  bfr _b_6476(.a(_w_7901),.q(_w_7902));
  bfr _b_4164(.a(_w_5589),.q(_w_5590));
  spl2 G153_s_0(.a(_w_6640),.q0(G153_0),.q1(_w_3917));
  bfr _b_4166(.a(_w_5591),.q(_w_5592));
  bfr _b_4541(.a(_w_5966),.q(_w_5967));
  spl3L g459_s_0(.a(n459),.q0(n459_0),.q1(_w_3478),.q2(_w_3483));
  or_bb g944(.a(n942),.b(n943),.q(n944));
  bfr _b_3697(.a(_w_5122),.q(_w_5123));
  bfr _b_4564(.a(_w_5989),.q(n1266));
  bfr _b_4167(.a(_w_5592),.q(_w_5593));
  bfr _b_2695(.a(_w_4120),.q(_w_4121));
  bfr _b_4661(.a(_w_6086),.q(_w_6087));
  bfr _b_4168(.a(_w_5593),.q(_w_5594));
  and_bi g1438(.a(n1437),.b(n1435),.q(n1438));
  bfr _b_4869(.a(_w_6294),.q(n1131));
  bfr _b_4172(.a(_w_5597),.q(_w_5598));
  bfr _b_4173(.a(_w_5598),.q(_w_5599));
  bfr _b_4175(.a(_w_5600),.q(_w_5601));
  bfr _b_4176(.a(_w_5601),.q(_w_5602));
  bfr _b_4177(.a(_w_5602),.q(_w_5603));
  bfr _b_4786(.a(_w_6211),.q(n1036));
  bfr _b_4182(.a(_w_5607),.q(_w_5608));
  bfr _b_7462(.a(_w_8887),.q(_w_8888));
  bfr _b_2335(.a(_w_3760),.q(_w_3761));
  bfr _b_4225(.a(_w_5650),.q(_w_5651));
  bfr _b_4186(.a(_w_5611),.q(_w_5612));
  or_bb g1387(.a(G100_8),.b(G105_10),.q(n1387));
  bfr _b_4427(.a(_w_5852),.q(_w_5853));
  bfr _b_6022(.a(G31),.q(_w_7448));
  bfr _b_2030(.a(_w_3455),.q(_w_3456));
  bfr _b_3728(.a(_w_5153),.q(n235));
  and_ii g990(.a(n985),.b(n989),.q(_w_6307));
  bfr _b_4187(.a(_w_5612),.q(_w_5613));
  bfr _b_7358(.a(_w_8783),.q(_w_8784));
  bfr _b_4188(.a(_w_5613),.q(G5237));
  bfr _b_4190(.a(_w_5615),.q(n1288));
  or_bb g1434(.a(n1432),.b(n1433),.q(n1434));
  bfr _b_4192(.a(_w_5617),.q(_w_5618));
  or_bb g363(.a(n361),.b(n362),.q(n363));
  bfr _b_4809(.a(_w_6234),.q(n243_1));
  bfr _b_4193(.a(_w_5618),.q(_w_5619));
  bfr _b_4194(.a(_w_5619),.q(_w_5620));
  bfr _b_4195(.a(_w_5620),.q(_w_5621));
  bfr _b_4199(.a(_w_5624),.q(_w_5625));
  bfr _b_4130(.a(_w_5555),.q(_w_5556));
  bfr _b_4512(.a(_w_5937),.q(_w_5938));
  bfr _b_4984(.a(G113),.q(_w_6410));
  bfr _b_3235(.a(_w_4660),.q(_w_4661));
  bfr _b_2636(.a(_w_4061),.q(_w_4062));
  bfr _b_4201(.a(_w_5626),.q(_w_5627));
  bfr _b_4849(.a(_w_6274),.q(G5300));
  spl2 g1252_s_0(.a(n1252),.q0(n1252_0),.q1(n1252_1));
  bfr _b_4205(.a(_w_5630),.q(_w_5631));
  bfr _b_1984(.a(_w_3409),.q(_w_3410));
  bfr _b_4206(.a(_w_5631),.q(_w_5632));
  spl2 G100_s_5(.a(G100_19),.q0(G100_20),.q1(G100_21));
  bfr _b_4209(.a(_w_5634),.q(_w_5635));
  bfr _b_4212(.a(_w_5637),.q(_w_5638));
  bfr _b_6779(.a(_w_8204),.q(_w_8205));
  bfr _b_5420(.a(_w_6845),.q(_w_6846));
  bfr _b_4213(.a(_w_5638),.q(_w_5639));
  bfr _b_4219(.a(_w_5644),.q(_w_5645));
  bfr _b_6929(.a(_w_8354),.q(_w_8355));
  bfr _b_4220(.a(_w_5645),.q(_w_5646));
  bfr _b_4221(.a(_w_5646),.q(_w_5647));
  bfr _b_4222(.a(_w_5647),.q(_w_5648));
  bfr _b_4224(.a(_w_5649),.q(_w_5650));
  and_bi g1230(.a(G150_5),.b(n1229),.q(n1230));
  bfr _b_4227(.a(_w_5652),.q(_w_5653));
  bfr _b_4231(.a(_w_5656),.q(_w_5657));
  bfr _b_4233(.a(_w_5658),.q(_w_5659));
  bfr _b_4235(.a(_w_5660),.q(_w_5661));
  bfr _b_5984(.a(G28),.q(_w_7410));
  bfr _b_4390(.a(_w_5815),.q(_w_5816));
  or_bb g374(.a(G141_4),.b(n372_1),.q(n374));
  bfr _b_4240(.a(_w_5665),.q(_w_5666));
  bfr _b_4241(.a(_w_5666),.q(G148_2));
  bfr _b_4242(.a(_w_5667),.q(_w_5668));
  bfr _b_4385(.a(_w_5810),.q(_w_5811));
  bfr _b_4243(.a(_w_5668),.q(n375));
  bfr _b_6577(.a(_w_8002),.q(_w_8003));
  bfr _b_3973(.a(_w_5398),.q(_w_5399));
  bfr _b_3494(.a(_w_4919),.q(_w_4920));
  bfr _b_4244(.a(_w_5669),.q(_w_5670));
  bfr _b_5864(.a(_w_7289),.q(_w_7290));
  bfr _b_4245(.a(_w_5670),.q(_w_5671));
  bfr _b_4456(.a(_w_5881),.q(G88_4));
  bfr _b_4246(.a(_w_5671),.q(_w_5672));
  and_bi g795(.a(n794),.b(n789_0),.q(_w_5902));
  bfr _b_4247(.a(_w_5672),.q(_w_5673));
  bfr _b_4248(.a(_w_5673),.q(n413_1));
  bfr _b_2721(.a(_w_4146),.q(_w_4147));
  bfr _b_4249(.a(_w_5674),.q(_w_5675));
  bfr _b_4251(.a(_w_5676),.q(_w_5677));
  bfr _b_4254(.a(_w_5679),.q(_w_5680));
  spl4L g804_s_0(.a(n804),.q0(n804_0),.q1(n804_1),.q2(n804_2),.q3(n804_3));
  bfr _b_4257(.a(_w_5682),.q(_w_5683));
  bfr _b_5097(.a(_w_6522),.q(_w_6523));
  bfr _b_4258(.a(_w_5683),.q(_w_5684));
  bfr _b_4320(.a(_w_5745),.q(_w_5746));
  bfr _b_4262(.a(_w_5687),.q(_w_5688));
  bfr _b_5132(.a(_w_6557),.q(_w_6558));
  spl4L G174_s_5(.a(G174_18),.q0(_w_3735),.q1(G174_21),.q2(G174_22),.q3(G174_23));
  bfr _b_2345(.a(_w_3770),.q(_w_3771));
  bfr _b_4265(.a(_w_5690),.q(_w_5691));
  bfr _b_5935(.a(_w_7360),.q(_w_7361));
  bfr _b_4268(.a(_w_5693),.q(_w_5694));
  bfr _b_3301(.a(_w_4726),.q(_w_4727));
  or_bb g1453(.a(n1451),.b(n1452),.q(_w_6298));
  bfr _b_4270(.a(_w_5695),.q(_w_5696));
  bfr _b_2009(.a(_w_3434),.q(_w_3435));
  bfr _b_4701(.a(_w_6126),.q(_w_6127));
  bfr _b_4271(.a(_w_5696),.q(_w_5697));
  bfr _b_4272(.a(_w_5697),.q(_w_5698));
  bfr _b_4274(.a(_w_5699),.q(n812));
  bfr _b_6048(.a(_w_7473),.q(_w_7474));
  bfr _b_4751(.a(_w_6176),.q(n1013));
  bfr _b_7261(.a(_w_8686),.q(_w_8687));
  or_bb g635(.a(n629),.b(n634),.q(_w_4614));
  bfr _b_2077(.a(_w_3502),.q(_w_3503));
  bfr _b_4277(.a(_w_5702),.q(n1110));
  bfr _b_4384(.a(_w_5809),.q(_w_5810));
  bfr _b_4281(.a(_w_5706),.q(G5297));
  bfr _b_4282(.a(_w_5707),.q(n677));
  bfr _b_2056(.a(_w_3481),.q(_w_3482));
  bfr _b_3639(.a(_w_5064),.q(_w_5065));
  bfr _b_4944(.a(_w_6369),.q(_w_6370));
  bfr _b_6383(.a(_w_7808),.q(_w_7809));
  bfr _b_4198(.a(_w_5623),.q(G5285_0));
  bfr _b_4290(.a(_w_5715),.q(_w_5716));
  bfr _b_4291(.a(_w_5716),.q(_w_5717));
  bfr _b_5550(.a(G172),.q(_w_6976));
  bfr _b_4292(.a(_w_5717),.q(_w_5718));
  bfr _b_5716(.a(_w_7141),.q(_w_7142));
  bfr _b_4294(.a(_w_5719),.q(_w_5720));
  bfr _b_4297(.a(_w_5722),.q(_w_5723));
  bfr _b_4299(.a(_w_5724),.q(_w_5725));
  and_bb g997(.a(G155_0),.b(G99_0),.q(n997));
  bfr _b_4301(.a(_w_5726),.q(_w_5727));
  and_bb g543(.a(n430_1),.b(n542_0),.q(n543));
  bfr _b_5049(.a(_w_6474),.q(_w_6475));
  bfr _b_3202(.a(_w_4627),.q(_w_4628));
  bfr _b_4302(.a(_w_5727),.q(_w_5728));
  bfr _b_5745(.a(_w_7170),.q(_w_7171));
  bfr _b_4306(.a(_w_5731),.q(_w_5732));
  bfr _b_4350(.a(_w_5775),.q(_w_5776));
  bfr _b_4307(.a(_w_5732),.q(_w_5733));
  bfr _b_4913(.a(_w_6338),.q(_w_6339));
  bfr _b_4309(.a(_w_5734),.q(_w_5735));
  bfr _b_6818(.a(_w_8243),.q(_w_8244));
  bfr _b_6570(.a(_w_7995),.q(_w_7996));
  bfr _b_5147(.a(_w_6572),.q(_w_6573));
  and_bb g898(.a(G82_0),.b(n804_4),.q(n898));
  bfr _b_2785(.a(_w_4210),.q(_w_4211));
  bfr _b_2559(.a(_w_3984),.q(_w_3985));
  bfr _b_4311(.a(_w_5736),.q(_w_5737));
  and_bb g403(.a(n375_0),.b(n402_0),.q(n403));
  bfr _b_3586(.a(_w_5011),.q(_w_5012));
  bfr _b_4688(.a(_w_6113),.q(G5281));
  bfr _b_4314(.a(_w_5739),.q(_w_5740));
  bfr _b_7249(.a(_w_8674),.q(_w_8675));
  bfr _b_3595(.a(_w_5020),.q(_w_5021));
  bfr _b_4554(.a(_w_5979),.q(_w_5980));
  and_bi g1456(.a(G174_5),.b(n1447_1),.q(n1456));
  bfr _b_4641(.a(_w_6066),.q(_w_6067));
  bfr _b_4316(.a(_w_5741),.q(_w_5742));
  bfr _b_6116(.a(_w_7541),.q(_w_7542));
  bfr _b_4318(.a(_w_5743),.q(n643_1));
  bfr _b_2565(.a(_w_3990),.q(_w_3991));
  bfr _b_4319(.a(_w_5744),.q(n643_2));
  bfr _b_4322(.a(_w_5747),.q(n527));
  and_bi g1264(.a(n552_6),.b(_w_7897),.q(_w_5884));
  and_bi g646(.a(n645_0),.b(G176_47),.q(n646));
  bfr _b_4326(.a(_w_5751),.q(n664));
  bfr _b_4329(.a(_w_5754),.q(_w_5755));
  bfr _b_3014(.a(_w_4439),.q(_w_4440));
  bfr _b_4333(.a(_w_5758),.q(G5306));
  bfr _b_4334(.a(_w_5759),.q(_w_5760));
  bfr _b_4336(.a(_w_5761),.q(_w_5762));
  bfr _b_3279(.a(_w_4704),.q(n458_2));
  bfr _b_4338(.a(_w_5763),.q(_w_5764));
  bfr _b_7185(.a(_w_8610),.q(_w_8611));
  bfr _b_3786(.a(_w_5211),.q(_w_5212));
  bfr _b_4340(.a(_w_5765),.q(n985));
  bfr _b_4315(.a(_w_5740),.q(_w_5741));
  bfr _b_4341(.a(_w_5766),.q(n414));
  bfr _b_7377(.a(_w_8802),.q(_w_8803));
  bfr _b_6752(.a(_w_8177),.q(_w_8178));
  spl4L G119_s_1(.a(G119_3),.q0(G119_4),.q1(G119_5),.q2(G119_6),.q3(G119_7));
  bfr _b_4342(.a(_w_5767),.q(_w_5768));
  spl4L G102_s_3(.a(G102_2),.q0(G102_11),.q1(G102_12),.q2(G102_13),.q3(G102_14));
  bfr _b_4343(.a(_w_5768),.q(_w_5769));
  bfr _b_4344(.a(_w_5769),.q(n1436));
  bfr _b_5858(.a(_w_7283),.q(_w_7284));
  bfr _b_4348(.a(_w_5773),.q(_w_5774));
  bfr _b_6644(.a(_w_8069),.q(_w_8070));
  bfr _b_4352(.a(_w_5777),.q(_w_5778));
  spl2 g415_s_1(.a(n415_3),.q0(n415_4),.q1(n415_5));
  bfr _b_4388(.a(_w_5813),.q(_w_5814));
  bfr _b_4668(.a(_w_6093),.q(_w_6094));
  and_bb g612(.a(G176_34),.b(n256_1),.q(n612));
  bfr _b_4354(.a(_w_5779),.q(_w_5780));
  bfr _b_4632(.a(_w_6057),.q(_w_6058));
  bfr _b_4356(.a(_w_5781),.q(_w_5782));
  bfr _b_4358(.a(_w_5783),.q(_w_5784));
  bfr _b_6445(.a(_w_7870),.q(_w_7871));
  spl2 g740_s_0(.a(n740),.q0(n740_0),.q1(n740_1));
  bfr _b_3709(.a(_w_5134),.q(_w_5135));
  bfr _b_4280(.a(_w_5705),.q(_w_5706));
  bfr _b_4359(.a(_w_5784),.q(_w_5785));
  bfr _b_4413(.a(_w_5838),.q(_w_5839));
  bfr _b_2793(.a(_w_4218),.q(_w_4219));
  bfr _b_4161(.a(_w_5586),.q(n974));
  bfr _b_4362(.a(_w_5787),.q(_w_5788));
  bfr _b_6855(.a(_w_8280),.q(_w_8281));
  bfr _b_4363(.a(_w_5788),.q(_w_5789));
  or_bb g1297(.a(n1279),.b(n1296),.q(_w_4316));
  bfr _b_4365(.a(_w_5790),.q(_w_5791));
  bfr _b_6880(.a(_w_8305),.q(_w_8306));
  bfr _b_6617(.a(_w_8042),.q(_w_8043));
  bfr _b_2194(.a(_w_3619),.q(_w_3620));
  bfr _b_3225(.a(_w_4650),.q(_w_4651));
  bfr _b_4367(.a(_w_5792),.q(_w_5793));
  bfr _b_3361(.a(_w_4786),.q(_w_4787));
  bfr _b_4370(.a(_w_5795),.q(_w_5796));
  bfr _b_2169(.a(_w_3594),.q(G125_2));
  bfr _b_4372(.a(_w_5797),.q(_w_5798));
  bfr _b_6167(.a(_w_7592),.q(_w_7593));
  bfr _b_4375(.a(_w_5800),.q(_w_5801));
  bfr _b_3136(.a(_w_4561),.q(n596));
  bfr _b_4695(.a(_w_6120),.q(_w_6121));
  bfr _b_2919(.a(_w_4344),.q(n1205));
  bfr _b_4379(.a(_w_5804),.q(G5228));
  bfr _b_4387(.a(_w_5812),.q(_w_5813));
  bfr _b_4393(.a(_w_5818),.q(_w_5819));
  bfr _b_4964(.a(_w_6389),.q(_w_6390));
  bfr _b_4398(.a(_w_5823),.q(_w_5824));
  and_bi g1398(.a(n1397),.b(n1396),.q(_w_6021));
  bfr _b_4400(.a(_w_5825),.q(G5238_0));
  bfr _b_4139(.a(_w_5564),.q(_w_5565));
  bfr _b_4404(.a(_w_5829),.q(_w_5830));
  bfr _b_4127(.a(_w_5552),.q(_w_5553));
  bfr _b_2286(.a(_w_3711),.q(_w_3712));
  bfr _b_3631(.a(_w_5056),.q(_w_5057));
  bfr _b_4405(.a(_w_5830),.q(_w_5831));
  bfr _b_7540(.a(_w_8965),.q(_w_8966));
  bfr _b_6816(.a(_w_8241),.q(_w_8242));
  bfr _b_4408(.a(_w_5833),.q(_w_5834));
  bfr _b_6963(.a(_w_8388),.q(_w_8389));
  spl2 g431_s_0(.a(G5238_0),.q0(G5238),.q1(G5241));
  bfr _b_4411(.a(_w_5836),.q(G166_0));
  bfr _b_6730(.a(_w_8155),.q(_w_8156));
  bfr _b_4415(.a(_w_5840),.q(_w_5841));
  bfr _b_2803(.a(_w_4228),.q(n435_1));
  bfr _b_4002(.a(_w_5427),.q(_w_5428));
  bfr _b_4859(.a(_w_6284),.q(n1092));
  or_bb g256(.a(n254),.b(n255),.q(_w_6283));
  bfr _b_4417(.a(_w_5842),.q(_w_5843));
  spl3L G163_s_1(.a(G163_1),.q0(G163_4),.q1(G163_5),.q2(G163_6));
  bfr _b_4419(.a(_w_5844),.q(G5259));
  or_bb g1278(.a(G157_0),.b(n1277),.q(n1278));
  bfr _b_4685(.a(_w_6110),.q(_w_6111));
  bfr _b_4420(.a(_w_5845),.q(_w_5846));
  bfr _b_4988(.a(G115),.q(_w_6414));
  and_bb g1309(.a(n1300_0),.b(n1308_0),.q(n1309));
  bfr _b_4423(.a(_w_5848),.q(_w_5849));
  bfr _b_4425(.a(_w_5850),.q(_w_5851));
  bfr _b_4429(.a(_w_5854),.q(_w_5855));
  bfr _b_4435(.a(_w_5860),.q(_w_5861));
  bfr _b_4436(.a(_w_5861),.q(_w_5862));
  bfr _b_4438(.a(_w_5863),.q(_w_5864));
  bfr _b_2661(.a(_w_4086),.q(_w_4087));
  bfr _b_4439(.a(_w_5864),.q(_w_5865));
  bfr _b_5026(.a(_w_6451),.q(_w_6452));
  bfr _b_4443(.a(_w_5868),.q(n475));
  bfr _b_6830(.a(_w_8255),.q(_w_8256));
  bfr _b_4444(.a(_w_5869),.q(_w_5870));
  bfr _b_5539(.a(_w_6964),.q(_w_6965));
  bfr _b_4445(.a(_w_5870),.q(_w_5871));
  bfr _b_4446(.a(_w_5871),.q(_w_5872));
  bfr _b_6266(.a(_w_7691),.q(_w_7692));
  bfr _b_4448(.a(_w_5873),.q(_w_5874));
  bfr _b_6924(.a(_w_8349),.q(_w_8350));
  bfr _b_4450(.a(_w_5875),.q(n463_1));
  bfr _b_4454(.a(_w_5879),.q(n977));
  bfr _b_4203(.a(_w_5628),.q(n682));
  bfr _b_4457(.a(_w_5882),.q(n758));
  bfr _b_4459(.a(_w_5884),.q(_w_5885));
  bfr _b_4461(.a(_w_5886),.q(_w_5887));
  bfr _b_5242(.a(_w_6667),.q(_w_6668));
  bfr _b_4462(.a(_w_5887),.q(_w_5888));
  bfr _b_6990(.a(_w_8415),.q(_w_8416));
  bfr _b_6646(.a(_w_8071),.q(_w_8072));
  bfr _b_6041(.a(_w_7466),.q(_w_7467));
  bfr _b_4467(.a(_w_5892),.q(n1264));
  bfr _b_4468(.a(_w_5893),.q(_w_5894));
  bfr _b_2897(.a(_w_4322),.q(_w_4323));
  bfr _b_4469(.a(_w_5894),.q(_w_5895));
  spl2 G82_s_0(.a(_w_8739),.q0(G82_0),.q1(G82_1));
  bfr _b_4473(.a(_w_5898),.q(n1076));
  bfr _b_7283(.a(_w_8708),.q(_w_8709));
  bfr _b_5450(.a(_w_6875),.q(_w_6876));
  bfr _b_2319(.a(_w_3744),.q(G148_4));
  bfr _b_4477(.a(_w_5902),.q(n795));
  bfr _b_4481(.a(_w_5906),.q(G173_1));
  bfr _b_2068(.a(_w_3493),.q(_w_3494));
  bfr _b_4482(.a(_w_5907),.q(_w_5908));
  bfr _b_4484(.a(_w_5909),.q(_w_5910));
  bfr _b_4491(.a(_w_5916),.q(_w_5917));
  bfr _b_4495(.a(_w_5920),.q(n1071));
  spl2 G11_s_0(.a(G11),.q0(G11_0),.q1(G11_1));
  bfr _b_4496(.a(_w_5921),.q(n801));
  bfr _b_4498(.a(_w_5923),.q(_w_5924));
  bfr _b_2497(.a(_w_3922),.q(G153_1));
  bfr _b_4012(.a(_w_5437),.q(n1303_0));
  bfr _b_4501(.a(_w_5926),.q(n451_2));
  bfr _b_4504(.a(_w_5929),.q(_w_5930));
  bfr _b_3398(.a(_w_4823),.q(_w_4824));
  bfr _b_4505(.a(_w_5930),.q(_w_5931));
  bfr _b_4507(.a(_w_5932),.q(_w_5933));
  bfr _b_6433(.a(_w_7858),.q(_w_7859));
  bfr _b_3016(.a(_w_4441),.q(_w_4442));
  bfr _b_4638(.a(_w_6063),.q(_w_6064));
  bfr _b_4511(.a(_w_5936),.q(_w_5937));
  bfr _b_4514(.a(_w_5939),.q(_w_5940));
  bfr _b_2426(.a(_w_3851),.q(_w_3852));
  bfr _b_3271(.a(_w_4696),.q(_w_4697));
  bfr _b_4515(.a(_w_5940),.q(_w_5941));
  bfr _b_3421(.a(_w_4846),.q(_w_4847));
  bfr _b_4516(.a(_w_5941),.q(_w_5942));
  bfr _b_4521(.a(_w_5946),.q(n637_0));
  bfr _b_4522(.a(_w_5947),.q(_w_5948));
  spl4L G158_s_0(.a(_w_6757),.q0(_w_3671),.q1(_w_3673),.q2(_w_3675),.q3(G158_3));
  bfr _b_4527(.a(_w_5952),.q(_w_5953));
  bfr _b_5911(.a(_w_7336),.q(_w_7337));
  bfr _b_2316(.a(_w_3741),.q(G174_18));
  bfr _b_4656(.a(_w_6081),.q(_w_6082));
  bfr _b_4528(.a(_w_5953),.q(_w_5954));
  bfr _b_3676(.a(_w_5101),.q(_w_5102));
  bfr _b_4530(.a(_w_5955),.q(_w_5956));
  and_bb g179(.a(G153_0),.b(G156_0),.q(G5199_0));
  bfr _b_4918(.a(_w_6343),.q(_w_6344));
  bfr _b_4534(.a(_w_5959),.q(_w_5960));
  bfr _b_4536(.a(_w_5961),.q(_w_5962));
  bfr _b_2868(.a(_w_4293),.q(_w_4294));
  bfr _b_4563(.a(_w_5988),.q(_w_5989));
  bfr _b_4537(.a(_w_5962),.q(_w_5963));
  bfr _b_4538(.a(_w_5963),.q(_w_5964));
  bfr _b_4542(.a(_w_5967),.q(_w_5968));
  bfr _b_4548(.a(_w_5973),.q(_w_5974));
  bfr _b_4549(.a(_w_5974),.q(_w_5975));
  bfr _b_4955(.a(_w_6380),.q(_w_6381));
  bfr _b_7250(.a(_w_8675),.q(_w_8676));
  bfr _b_3738(.a(_w_5163),.q(_w_5164));
  bfr _b_4289(.a(_w_5714),.q(_w_5715));
  bfr _b_4550(.a(_w_5975),.q(_w_5976));
  bfr _b_2657(.a(_w_4082),.q(_w_4083));
  bfr _b_4552(.a(_w_5977),.q(_w_5978));
  bfr _b_4553(.a(_w_5978),.q(_w_5979));
  bfr _b_4555(.a(_w_5980),.q(n199));
  bfr _b_4558(.a(_w_5983),.q(n839));
  bfr _b_4569(.a(_w_5994),.q(_w_5995));
  bfr _b_2866(.a(_w_4291),.q(_w_4292));
  bfr _b_4645(.a(_w_6070),.q(_w_6071));
  spl2 g1362_s_0(.a(n1362),.q0(n1362_0),.q1(n1362_1));
  bfr _b_4570(.a(_w_5995),.q(_w_5996));
  bfr _b_4667(.a(_w_6092),.q(_w_6093));
  bfr _b_4575(.a(_w_6000),.q(_w_6001));
  bfr _b_4579(.a(_w_6004),.q(_w_6005));
  bfr _b_4582(.a(_w_6007),.q(_w_6008));
  bfr _b_3196(.a(_w_4621),.q(_w_4622));
  bfr _b_4586(.a(_w_6011),.q(n1253));
  bfr _b_5170(.a(_w_6595),.q(_w_6596));
  bfr _b_4588(.a(_w_6013),.q(_w_6014));
  bfr _b_4590(.a(_w_6015),.q(_w_6016));
  bfr _b_4592(.a(_w_6017),.q(_w_6018));
  bfr _b_4596(.a(_w_6021),.q(_w_6022));
  bfr _b_4805(.a(_w_6230),.q(_w_6231));
  bfr _b_4597(.a(_w_6022),.q(_w_6023));
  bfr _b_4598(.a(_w_6023),.q(n1398));
  bfr _b_4599(.a(_w_6024),.q(_w_6025));
  bfr _b_4973(.a(G106),.q(_w_6399));
  bfr _b_4602(.a(_w_6027),.q(G146_3));
  bfr _b_4605(.a(_w_6030),.q(G5272));
  bfr _b_4610(.a(_w_6035),.q(_w_6036));
  bfr _b_6842(.a(_w_8267),.q(_w_8268));
  spl4L G128_s_2(.a(G128_2),.q0(G128_6),.q1(_w_3905),.q2(G128_8),.q3(G128_9));
  bfr _b_4613(.a(_w_6038),.q(_w_6039));
  bfr _b_4615(.a(_w_6040),.q(G5286));
  bfr _b_2869(.a(_w_4294),.q(G138_2));
  bfr _b_4616(.a(_w_6041),.q(n556_0));
  bfr _b_6341(.a(_w_7766),.q(_w_7767));
  bfr _b_4120(.a(_w_5545),.q(_w_5546));
  bfr _b_4784(.a(_w_6209),.q(_w_6210));
  bfr _b_5213(.a(_w_6638),.q(_w_6639));
  bfr _b_4619(.a(_w_6044),.q(n648));
  or_bb g473(.a(n469_0),.b(n472_0),.q(n473));
  bfr _b_4621(.a(_w_6046),.q(n891));
  bfr _b_4519(.a(_w_5944),.q(n545_1));
  bfr _b_4629(.a(_w_6054),.q(_w_6055));
  bfr _b_4631(.a(_w_6056),.q(_w_6057));
  bfr _b_4633(.a(_w_6058),.q(_w_6059));
  bfr _b_5625(.a(_w_7050),.q(_w_7051));
  bfr _b_4634(.a(_w_6059),.q(_w_6060));
  bfr _b_5160(.a(_w_6585),.q(_w_6586));
  bfr _b_4635(.a(_w_6060),.q(_w_6061));
  bfr _b_7378(.a(_w_8803),.q(_w_8804));
  bfr _b_3207(.a(_w_4632),.q(_w_4633));
  bfr _b_4636(.a(_w_6061),.q(_w_6062));
  bfr _b_4639(.a(_w_6064),.q(G5263));
  bfr _b_5924(.a(_w_7349),.q(_w_7350));
  bfr _b_4640(.a(_w_6065),.q(n573));
  bfr _b_3079(.a(_w_4504),.q(_w_4505));
  bfr _b_4642(.a(_w_6067),.q(n927));
  bfr _b_4643(.a(_w_6068),.q(n932));
  bfr _b_4650(.a(_w_6075),.q(_w_6076));
  and_bi g1149(.a(n1148),.b(n1146),.q(_w_4354));
  bfr _b_2688(.a(_w_4113),.q(_w_4114));
  bfr _b_4655(.a(_w_6080),.q(_w_6081));
  bfr _b_7248(.a(G80),.q(_w_8674));
  bfr _b_4658(.a(_w_6083),.q(n1443));
  bfr _b_4664(.a(_w_6089),.q(_w_6090));
  bfr _b_4666(.a(_w_6091),.q(_w_6092));
  bfr _b_5312(.a(_w_6737),.q(_w_6738));
  and_bi g295(.a(G166_8),.b(G90_6),.q(n295));
  bfr _b_4670(.a(_w_6095),.q(_w_6096));
  bfr _b_4673(.a(_w_6098),.q(n963));
  bfr _b_2775(.a(_w_4200),.q(_w_4201));
  bfr _b_4674(.a(_w_6099),.q(G5280));
  bfr _b_4676(.a(_w_6101),.q(_w_6102));
  bfr _b_2466(.a(_w_3891),.q(_w_3892));
  bfr _b_4677(.a(_w_6102),.q(G5295));
  bfr _b_4900(.a(_w_6325),.q(_w_6326));
  bfr _b_4678(.a(_w_6103),.q(n941));
  bfr _b_4851(.a(_w_6276),.q(n1084));
  bfr _b_4680(.a(_w_6105),.q(_w_6106));
  bfr _b_2190(.a(_w_3615),.q(_w_3616));
  bfr _b_4683(.a(_w_6108),.q(_w_6109));
  bfr _b_4687(.a(_w_6112),.q(G5250));
  bfr _b_6894(.a(_w_8319),.q(_w_8320));
  bfr _b_4689(.a(_w_6114),.q(G149_4));
  bfr _b_4690(.a(_w_6115),.q(n1087));
  bfr _b_4693(.a(_w_6118),.q(_w_6119));
  bfr _b_4702(.a(_w_6127),.q(_w_6128));
  bfr _b_6286(.a(_w_7711),.q(_w_7712));
  bfr _b_4749(.a(_w_6174),.q(_w_6175));
  spl2 G167_s_1(.a(G167_1),.q0(G167_4),.q1(G167_5));
  bfr _b_4857(.a(_w_6282),.q(G5301));
  bfr _b_4706(.a(_w_6131),.q(_w_6132));
  bfr _b_4713(.a(_w_6138),.q(n379_3));
  bfr _b_4716(.a(_w_6141),.q(_w_6142));
  bfr _b_4722(.a(_w_6147),.q(_w_6148));
  bfr _b_4724(.a(_w_6149),.q(_w_6150));
  or_bb g1455(.a(G174_6),.b(n1444_1),.q(n1455));
  bfr _b_4729(.a(_w_6154),.q(_w_6155));
  bfr _b_2644(.a(_w_4069),.q(_w_4070));
  bfr _b_4705(.a(_w_6130),.q(_w_6131));
  bfr _b_4731(.a(_w_6156),.q(n556));
  and_bi g377(.a(_w_6403),.b(G124_23),.q(n377));
  bfr _b_4732(.a(_w_6157),.q(_w_6158));
  bfr _b_5520(.a(_w_6945),.q(_w_6946));
  and_bi g611(.a(n610_0),.b(G176_43),.q(n611));
  bfr _b_4733(.a(_w_6158),.q(_w_6159));
  or_bb g867(.a(n863),.b(n866),.q(_w_6028));
  bfr _b_4735(.a(_w_6160),.q(_w_6161));
  bfr _b_3563(.a(_w_4988),.q(_w_4989));
  bfr _b_4736(.a(_w_6161),.q(_w_6162));
  bfr _b_5221(.a(_w_6646),.q(_w_6647));
  bfr _b_2972(.a(_w_4397),.q(_w_4398));
  bfr _b_4022(.a(_w_5447),.q(_w_5448));
  bfr _b_4737(.a(_w_6162),.q(_w_6163));
  or_bb g936(.a(n932),.b(n935),.q(n936));
  bfr _b_4738(.a(_w_6163),.q(n1010));
  bfr _b_4739(.a(_w_6164),.q(_w_6165));
  bfr _b_4740(.a(_w_6165),.q(n624));
  bfr _b_4741(.a(_w_6166),.q(_w_6167));
  and_ii g675(.a(n664),.b(n674),.q(_w_5443));
  bfr _b_4744(.a(_w_6169),.q(_w_6170));
  bfr _b_3669(.a(_w_5094),.q(_w_5095));
  bfr _b_3730(.a(_w_5155),.q(n212));
  bfr _b_4746(.a(_w_6171),.q(n1012));
  bfr _b_4752(.a(_w_6177),.q(_w_6178));
  bfr _b_4757(.a(_w_6182),.q(_w_6183));
  bfr _b_4759(.a(_w_6184),.q(_w_6185));
  bfr _b_4959(.a(_w_6384),.q(_w_6385));
  bfr _b_4765(.a(_w_6190),.q(G5292_0));
  bfr _b_3848(.a(_w_5273),.q(_w_5274));
  bfr _b_2797(.a(_w_4222),.q(_w_4223));
  bfr _b_4768(.a(_w_6193),.q(_w_6194));
  spl2 g984_s_1(.a(G5286_3),.q0(G5286_4),.q1(G5286_5));
  bfr _b_2524(.a(_w_3949),.q(_w_3950));
  bfr _b_4769(.a(_w_6194),.q(_w_6195));
  bfr _b_2478(.a(_w_3903),.q(_w_3904));
  bfr _b_4772(.a(_w_6197),.q(_w_6198));
  bfr _b_4773(.a(_w_6198),.q(G5273));
  bfr _b_4691(.a(_w_6116),.q(_w_6117));
  bfr _b_4775(.a(_w_6200),.q(_w_6201));
  bfr _b_2516(.a(_w_3941),.q(G88_1));
  bfr _b_4787(.a(_w_6212),.q(_w_6213));
  bfr _b_6768(.a(_w_8193),.q(_w_8194));
  spl4L g372_s_0(.a(n372),.q0(n372_0),.q1(n372_1),.q2(n372_2),.q3(n372_3));
  and_bi g716(.a(n715),.b(n714),.q(n716));
  spl2 G14_s_0(.a(_w_6493),.q0(G14_0),.q1(G14_1));
  bfr _b_4791(.a(_w_6216),.q(_w_6217));
  bfr _b_4793(.a(_w_6218),.q(_w_6219));
  bfr _b_4797(.a(_w_6222),.q(n1313));
  bfr _b_4798(.a(_w_6223),.q(_w_6224));
  bfr _b_4799(.a(_w_6224),.q(_w_6225));
  bfr _b_7304(.a(_w_8729),.q(_w_8730));
  bfr _b_3875(.a(_w_5300),.q(_w_5301));
  bfr _b_5039(.a(_w_6464),.q(_w_6465));
  bfr _b_5746(.a(_w_7171),.q(_w_7172));
  bfr _b_4800(.a(_w_6225),.q(G5296));
  bfr _b_2417(.a(_w_3842),.q(_w_3843));
  bfr _b_4801(.a(_w_6226),.q(n1052));
  bfr _b_6233(.a(_w_7658),.q(_w_7659));
  bfr _b_5595(.a(_w_7020),.q(_w_7021));
  and_bi g1433(.a(n1398_1),.b(n1431_1),.q(n1433));
  bfr _b_4802(.a(_w_6227),.q(n187));
  bfr _b_4804(.a(_w_6229),.q(n1165));
  bfr _b_5522(.a(_w_6947),.q(_w_6948));
  bfr _b_4807(.a(_w_6232),.q(G5298));
  bfr _b_4808(.a(_w_6233),.q(_w_6234));
  bfr _b_5023(.a(_w_6448),.q(_w_6449));
  bfr _b_4811(.a(_w_6236),.q(_w_6237));
  bfr _b_4814(.a(_w_6239),.q(_w_6240));
  bfr _b_4815(.a(_w_6240),.q(_w_6241));
  bfr _b_6846(.a(_w_8271),.q(_w_8272));
  bfr _b_4818(.a(_w_6243),.q(_w_6244));
  bfr _b_5773(.a(_w_7198),.q(_w_7199));
  bfr _b_4819(.a(_w_6244),.q(_w_6245));
  bfr _b_4825(.a(_w_6250),.q(_w_6251));
  bfr _b_5966(.a(_w_7391),.q(_w_7392));
  bfr _b_5001(.a(_w_6426),.q(_w_6427));
  bfr _b_4826(.a(_w_6251),.q(_w_6252));
  bfr _b_2224(.a(_w_3649),.q(_w_3650));
  bfr _b_4828(.a(_w_6253),.q(_w_6254));
  spl2 g579_s_1(.a(G5250_3),.q0(G5250_4),.q1(G5250_5));
  bfr _b_4830(.a(_w_6255),.q(_w_6256));
  bfr _b_5047(.a(_w_6472),.q(_w_6473));
  and_bi g837(.a(G173_17),.b(G5255_1),.q(n837));
  bfr _b_4285(.a(_w_5710),.q(_w_5711));
  bfr _b_4832(.a(_w_6257),.q(_w_6258));
  bfr _b_7366(.a(_w_8791),.q(_w_8792));
  bfr _b_4841(.a(_w_6266),.q(_w_6267));
  and_bi g232(.a(n231),.b(G146_1),.q(n232));
  bfr _b_4842(.a(_w_6267),.q(G5213_0));
  bfr _b_4846(.a(_w_6271),.q(n1079));
  bfr _b_4853(.a(_w_6278),.q(_w_6279));
  bfr _b_2747(.a(_w_4172),.q(_w_4173));
  bfr _b_2502(.a(_w_3927),.q(_w_3928));
  bfr _b_4861(.a(_w_6286),.q(n1104));
  bfr _b_4865(.a(_w_6290),.q(G5304));
  bfr _b_3919(.a(_w_5344),.q(_w_5345));
  bfr _b_4867(.a(_w_6292),.q(n1039));
  and_bb g914(.a(n911),.b(n913),.q(_w_6053));
  bfr _b_4870(.a(_w_6295),.q(n661));
  bfr _b_4873(.a(_w_6298),.q(_w_6299));
  bfr _b_4874(.a(_w_6299),.q(n1453));
  bfr _b_4882(.a(_w_6307),.q(G5287_0));
  bfr _b_4883(.a(_w_6308),.q(n1162));
  bfr _b_4884(.a(_w_6309),.q(n1179));
  bfr _b_6832(.a(_w_8257),.q(_w_8258));
  and_bi g1464(.a(G158_5),.b(n1447_2),.q(n1464));
  spl4L G177_s_4(.a(G177_3),.q0(G177_16),.q1(G177_17),.q2(G177_18),.q3(G177_19));
  bfr _b_2908(.a(_w_4333),.q(n337_1));
  bfr _b_4885(.a(_w_6310),.q(_w_6311));
  bfr _b_4890(.a(_w_6315),.q(_w_6316));
  bfr _b_6464(.a(_w_7889),.q(_w_7890));
  bfr _b_4441(.a(_w_5866),.q(_w_5867));
  bfr _b_4893(.a(_w_6318),.q(_w_6319));
  bfr _b_4895(.a(_w_6320),.q(_w_6321));
  bfr _b_4899(.a(_w_6324),.q(_w_6325));
  bfr _b_4901(.a(_w_6326),.q(n686));
  spl4L g465_s_0(.a(n465),.q0(_w_3452),.q1(_w_3455),.q2(_w_3461),.q3(n465_3));
  bfr _b_4902(.a(_w_6327),.q(n1223));
  bfr _b_4903(.a(_w_6328),.q(n1119));
  bfr _b_4904(.a(_w_6329),.q(n1258));
  bfr _b_4906(.a(_w_6331),.q(_w_6332));
  bfr _b_4909(.a(_w_6334),.q(G177_7));
  bfr _b_4910(.a(_w_6335),.q(_w_6336));
  bfr _b_4823(.a(_w_6248),.q(_w_6249));
  bfr _b_4911(.a(_w_6336),.q(_w_6337));
  bfr _b_4981(.a(G111),.q(_w_6406));
  bfr _b_4812(.a(_w_6237),.q(_w_6238));
  bfr _b_4914(.a(_w_6339),.q(n1250));
  bfr _b_2794(.a(_w_4219),.q(n415_2));
  bfr _b_4916(.a(_w_6341),.q(_w_6342));
  bfr _b_6166(.a(_w_7591),.q(_w_7592));
  bfr _b_4917(.a(_w_6342),.q(_w_6343));
  bfr _b_6903(.a(_w_8328),.q(_w_8329));
  bfr _b_4919(.a(_w_6344),.q(_w_6345));
  bfr _b_3409(.a(_w_4834),.q(_w_4835));
  bfr _b_4924(.a(_w_6349),.q(n1324_0));
  bfr _b_4926(.a(_w_6351),.q(_w_6352));
  bfr _b_4928(.a(_w_6353),.q(n1280));
  and_bi g854(.a(G175_6),.b(n853),.q(n854));
  bfr _b_4930(.a(_w_6355),.q(_w_6356));
  bfr _b_3741(.a(_w_5166),.q(_w_5167));
  bfr _b_4932(.a(_w_6357),.q(_w_6358));
  spl4L g545_s_0(.a(n545),.q0(n545_0),.q1(_w_5934),.q2(n545_2),.q3(n545_3));
  bfr _b_5081(.a(_w_6506),.q(_w_6507));
  bfr _b_6442(.a(_w_7867),.q(_w_7868));
  bfr _b_4935(.a(_w_6360),.q(_w_6361));
  bfr _b_4933(.a(_w_6358),.q(_w_6359));
  bfr _b_4938(.a(_w_6363),.q(_w_6364));
  bfr _b_4941(.a(_w_6366),.q(_w_6367));
  bfr _b_4942(.a(_w_6367),.q(_w_6368));
  bfr _b_6066(.a(G37),.q(_w_7492));
  bfr _b_4945(.a(_w_6370),.q(_w_6371));
  bfr _b_7317(.a(_w_8742),.q(_w_8743));
  bfr _b_4758(.a(_w_6183),.q(_w_6184));
  bfr _b_4946(.a(_w_6371),.q(_w_6372));
  spl3L g433_s_0(.a(n433),.q0(n433_0),.q1(n433_1),.q2(_w_4220));
  and_bb g392(.a(G138_2),.b(n391_0),.q(n392));
  bfr _b_4948(.a(_w_6373),.q(_w_6374));
  bfr _b_4952(.a(_w_6377),.q(_w_6378));
  bfr _b_4954(.a(_w_6379),.q(_w_6380));
  or_bb g809(.a(G160_15),.b(G5250_5),.q(n809));
  bfr _b_4960(.a(_w_6385),.q(_w_6386));
  bfr _b_5484(.a(_w_6909),.q(_w_6910));
  bfr _b_5306(.a(_w_6731),.q(_w_6732));
  bfr _b_4961(.a(_w_6386),.q(_w_6387));
  spl4L G173_s_5(.a(G173_18),.q0(_w_4306),.q1(G173_21),.q2(G173_22),.q3(G173_23));
  bfr _b_4963(.a(_w_6388),.q(_w_6389));
  bfr _b_4967(.a(_w_6392),.q(_w_6391));
  bfr _b_4968(.a(G100),.q(_w_6393));
  bfr _b_4970(.a(G102),.q(_w_6395));
  bfr _b_4971(.a(G104),.q(_w_6397));
  bfr _b_4972(.a(_w_6397),.q(_w_6396));
  bfr _b_2652(.a(_w_4077),.q(_w_4078));
  bfr _b_4975(.a(G108),.q(_w_6401));
  bfr _b_4976(.a(_w_6401),.q(_w_6402));
  bfr _b_2823(.a(_w_4248),.q(_w_4249));
  bfr _b_4977(.a(_w_6402),.q(_w_6400));
  bfr _b_4979(.a(_w_6404),.q(_w_6405));
  bfr _b_4980(.a(_w_6405),.q(_w_6403));
  and_bi g1040(.a(G41_1),.b(n588_7),.q(n1040));
  bfr _b_2375(.a(_w_3800),.q(_w_3801));
  bfr _b_4983(.a(_w_6408),.q(_w_6407));
  bfr _b_4990(.a(G116),.q(_w_6416));
  bfr _b_4998(.a(_w_6423),.q(_w_6422));
  bfr _b_3270(.a(_w_4695),.q(_w_4696));
  bfr _b_5003(.a(G122),.q(_w_6429));
  bfr _b_6563(.a(_w_7988),.q(_w_7989));
  bfr _b_5154(.a(_w_6579),.q(_w_6580));
  bfr _b_5005(.a(G125),.q(_w_6431));
  bfr _b_2234(.a(_w_3659),.q(_w_3660));
  bfr _b_4630(.a(_w_6055),.q(_w_6056));
  bfr _b_5006(.a(_w_6431),.q(_w_6432));
  bfr _b_5007(.a(_w_6432),.q(_w_6430));
  bfr _b_5008(.a(G127),.q(_w_6433));
  bfr _b_2141(.a(_w_3566),.q(_w_3567));
  bfr _b_5009(.a(G129),.q(_w_6435));
  bfr _b_5011(.a(G13),.q(_w_6437));
  and_bb g896(.a(n893),.b(n895),.q(_w_4830));
  and_bb g864(.a(G27_1),.b(n630_4),.q(n864));
  bfr _b_5012(.a(_w_6437),.q(_w_6436));
  bfr _b_2273(.a(_w_3698),.q(_w_3699));
  bfr _b_5016(.a(G133),.q(_w_6442));
  bfr _b_4694(.a(_w_6119),.q(_w_6120));
  bfr _b_5031(.a(_w_6456),.q(_w_6457));
  bfr _b_2180(.a(_w_3605),.q(_w_3606));
  bfr _b_5032(.a(_w_6457),.q(_w_6458));
  bfr _b_5073(.a(_w_6498),.q(_w_6499));
  bfr _b_2343(.a(_w_3768),.q(_w_3769));
  bfr _b_5035(.a(_w_6460),.q(_w_6461));
  bfr _b_5080(.a(_w_6505),.q(_w_6506));
  bfr _b_5036(.a(_w_6461),.q(_w_6462));
  bfr _b_6084(.a(_w_7509),.q(_w_7491));
  bfr _b_5038(.a(_w_6463),.q(_w_6464));
  bfr _b_5041(.a(_w_6466),.q(_w_6467));
  bfr _b_6340(.a(_w_7765),.q(_w_7766));
  bfr _b_5048(.a(_w_6473),.q(_w_6474));
  bfr _b_5705(.a(_w_7130),.q(_w_7131));
  bfr _b_5051(.a(_w_6476),.q(_w_6477));
  and_bb g477(.a(G147_2),.b(n476_0),.q(_w_4645));
  bfr _b_5053(.a(_w_6478),.q(_w_6479));
  bfr _b_6099(.a(_w_7524),.q(_w_7525));
  bfr _b_5055(.a(_w_6480),.q(_w_6443));
  bfr _b_3084(.a(_w_4509),.q(_w_4510));
  bfr _b_5056(.a(G135),.q(_w_6482));
  bfr _b_5057(.a(_w_6482),.q(_w_6483));
  bfr _b_2241(.a(_w_3666),.q(_w_3667));
  bfr _b_5059(.a(G137),.q(_w_6485));
  bfr _b_6669(.a(_w_8094),.q(_w_8095));
  bfr _b_5063(.a(_w_6488),.q(_w_6489));
  spl4L g984_s_0(.a(G5286_0),.q0(_w_6033),.q1(G5286_1),.q2(G5286_2),.q3(G5286_3));
  bfr _b_5065(.a(G139),.q(_w_6491));
  bfr _b_5130(.a(_w_6555),.q(_w_6556));
  bfr _b_5069(.a(_w_6494),.q(_w_6495));
  bfr _b_5077(.a(_w_6502),.q(_w_6503));
  spl4L G176_s_7(.a(G176_13),.q0(_w_3399),.q1(G176_27),.q2(_w_3404),.q3(G176_29));
  bfr _b_5079(.a(_w_6504),.q(_w_6505));
  spl4L G157_s_0(.a(_w_6736),.q0(G157_0),.q1(G157_1),.q2(G157_2),.q3(G157_3));
  bfr _b_5086(.a(_w_6511),.q(_w_6512));
endmodule
