module c6288 (N1,N103,N120,N137,N154,N171,N18,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N35,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N52,N528,N69,N86,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N545,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288);
  input N1,N103,N120,N137,N154,N171,N18,N188,N205,N222,N239,N256,N273,N290,N307,N324,N341,N35,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N52,N528,N69,N86;
  output N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N545,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288;
  wire _w_16288,_w_16286,_w_16285,_w_16283,_w_16281,_w_16279,_w_16278,_w_16276,_w_16275,_w_16274,_w_16273,_w_16269,_w_16268,_w_16263,_w_16260,_w_16259,_w_16255,_w_16247,_w_16244,_w_16240,_w_16236,_w_16235,_w_16234,_w_16233,_w_16231,_w_16229,_w_16227,_w_16224,_w_16223,_w_16220,_w_16219,_w_16218,_w_16213,_w_16207,_w_16203,_w_16201,_w_16198,_w_16197,_w_16194,_w_16191,_w_16190,_w_16189,_w_16188,_w_16187,_w_16185,_w_16182,_w_16179,_w_16178,_w_16177,_w_16175,_w_16165,_w_16163,_w_16161,_w_16159,_w_16151,_w_16150,_w_16149,_w_16148,_w_16146,_w_16144,_w_16142,_w_16136,_w_16135,_w_16134,_w_16133,_w_16125,_w_16123,_w_16122,_w_16116,_w_16111,_w_16109,_w_16107,_w_16105,_w_16104,_w_16102,_w_16097,_w_16096,_w_16093,_w_16092,_w_16089,_w_16088,_w_16087,_w_16256,_w_16086,_w_16084,_w_16082,_w_16080,_w_16077,_w_16074,_w_16072,_w_16070,_w_16068,_w_16067,_w_16066,_w_16065,_w_16064,_w_16063,_w_16060,_w_16057,_w_16056,_w_16054,_w_16052,_w_16051,_w_16050,_w_16047,_w_16039,_w_16038,_w_16036,_w_16035,_w_16033,_w_16032,_w_16027,_w_16025,_w_16023,_w_16022,_w_16020,_w_16019,_w_16013,_w_16009,_w_16008,_w_16007,_w_16005,_w_16003,_w_16000,_w_15999,_w_15998,_w_15994,_w_15992,_w_15991,_w_16121,_w_15990,_w_15989,_w_15986,_w_15984,_w_15983,_w_15982,_w_15981,_w_15978,_w_15977,_w_15976,_w_15974,_w_15973,_w_15972,_w_15971,_w_15969,_w_15965,_w_15960,_w_15958,_w_15957,_w_15956,_w_15955,_w_15954,_w_15949,_w_15948,_w_15946,_w_15945,_w_15944,_w_15943,_w_15941,_w_15935,_w_15924,_w_15920,_w_15919,_w_15916,_w_15915,_w_15914,_w_15913,_w_15910,_w_15907,_w_15906,_w_15905,_w_15903,_w_15902,_w_15901,_w_15898,_w_15897,_w_15895,_w_15890,_w_15886,_w_15882,_w_15877,_w_15874,_w_15873,_w_15872,_w_15868,_w_15866,_w_15863,_w_15862,_w_15858,_w_15857,_w_15849,_w_15844,_w_15843,_w_15840,_w_15835,_w_15830,_w_15828,_w_15826,_w_15825,_w_15823,_w_15822,_w_15821,_w_15820,_w_15816,_w_15815,_w_15814,_w_15810,_w_15808,_w_15807,_w_15805,_w_15804,_w_15803,_w_15802,_w_15800,_w_15799,_w_15798,_w_15795,_w_15789,_w_15788,_w_15780,_w_15779,_w_15778,_w_16001,_w_15777,_w_15776,_w_15775,_w_15774,_w_15772,_w_15768,_w_15766,_w_15765,_w_15764,_w_15763,_w_15761,_w_15760,_w_15757,_w_15756,_w_15755,_w_15754,_w_15753,_w_15752,_w_15741,_w_15740,_w_15739,_w_15738,_w_15730,_w_15723,_w_15722,_w_15721,_w_15719,_w_15715,_w_15713,_w_15710,_w_15709,_w_15707,_w_15702,_w_15699,_w_15697,_w_15691,_w_15687,_w_15682,_w_15676,_w_15673,_w_15668,_w_15666,_w_15665,_w_15664,_w_15662,_w_15661,_w_15660,_w_15659,_w_15658,_w_15657,_w_15654,_w_15650,_w_15649,_w_15648,_w_15642,_w_15641,_w_15640,_w_15639,_w_15638,_w_16258,_w_15636,_w_15632,_w_15631,_w_15629,_w_15628,_w_15627,_w_15626,_w_15624,_w_15620,_w_15617,_w_15610,_w_15609,_w_15605,_w_15603,_w_15601,_w_16204,_w_15600,_w_15599,_w_15598,_w_15596,_w_15594,_w_15635,_w_15593,_w_15592,_w_15591,_w_15590,_w_15586,_w_15583,_w_15581,_w_15578,_w_15576,_w_15571,_w_15567,_w_15566,_w_15562,_w_15561,_w_15558,_w_15557,_w_15554,_w_15553,_w_15552,_w_15550,_w_15549,_w_15548,_w_15547,_w_15790,_w_15546,_w_15545,_w_15544,_w_15541,_w_15540,_w_15539,_w_15536,_w_15533,_w_15531,_w_15529,_w_15527,_w_16004,_w_15526,_w_15525,_w_15521,_w_15519,_w_15518,_w_15516,_w_15511,_w_15509,_w_15497,_w_15494,_w_15492,_w_15491,_w_15490,_w_15489,_w_15488,_w_15483,_w_15482,_w_15481,_w_15479,_w_15475,_w_15474,_w_15801,_w_15472,_w_15468,_w_15467,_w_15466,_w_15463,_w_15462,_w_15461,_w_15459,_w_15457,_w_15456,_w_15453,_w_15452,_w_15450,_w_15449,_w_15448,_w_15447,_w_15446,_w_15445,_w_15444,_w_15443,_w_15442,_w_15441,_w_15440,_w_15437,_w_15434,_w_15742,_w_15433,_w_15431,_w_15430,_w_15425,_w_15423,_w_15422,_w_15421,_w_15419,_w_15415,_w_15412,_w_15408,_w_15407,_w_15403,_w_15401,_w_15398,_w_15396,_w_15395,_w_15394,_w_15393,_w_15392,_w_15390,_w_15389,_w_15385,_w_15542,_w_15383,_w_15380,_w_15379,_w_15377,_w_15376,_w_15375,_w_15369,_w_15368,_w_15367,_w_15366,_w_15881,_w_15359,_w_15356,_w_15353,_w_16140,_w_15352,_w_15346,_w_15343,_w_15339,_w_15337,_w_15331,_w_15329,_w_15327,_w_15326,_w_15324,_w_15646,_w_15319,_w_15317,_w_15314,_w_15313,_w_16059,_w_15311,_w_15310,_w_15309,_w_15308,_w_15307,_w_15306,_w_15305,_w_15304,_w_15302,_w_15301,_w_15299,_w_15298,_w_15926,_w_15297,_w_15294,_w_15287,_w_15286,_w_15284,_w_15283,_w_15281,_w_15279,_w_15277,_w_15276,_w_15275,_w_15273,_w_15272,_w_15271,_w_15267,_w_15265,_w_15262,_w_15260,_w_15259,_w_15256,_w_15255,_w_15250,_w_15244,_w_15242,_w_15438,_w_15240,_w_15238,_w_15237,_w_15230,_w_15228,_w_15226,_w_15225,_w_15224,_w_15221,_w_15218,_w_15217,_w_15216,_w_15211,_w_15210,_w_15209,_w_15208,_w_15207,_w_15206,_w_15204,_w_15414,_w_15202,_w_15201,_w_15200,_w_15199,_w_15198,_w_15195,_w_15194,_w_15193,_w_15191,_w_15190,_w_15189,_w_15186,_w_15181,_w_15179,_w_15177,_w_15176,_w_15172,_w_15170,_w_15168,_w_15165,_w_15164,_w_15162,_w_15161,_w_15160,_w_15157,_w_15156,_w_15155,_w_15153,_w_15152,_w_15151,_w_15149,_w_15147,_w_15145,_w_15143,_w_15140,_w_15137,_w_15136,_w_16280,_w_15135,_w_15130,_w_15129,_w_15127,_w_15120,_w_15117,_w_15115,_w_15111,_w_15110,_w_15109,_w_15188,_w_15108,_w_15107,_w_15106,_w_15105,_w_15102,_w_15093,_w_15092,_w_15091,_w_15084,_w_15083,_w_15082,_w_15282,_w_15080,_w_15079,_w_15078,_w_15077,_w_15076,_w_15073,_w_15072,_w_15070,_w_15067,_w_15063,_w_15062,_w_15060,_w_15058,_w_15056,_w_15054,_w_15053,_w_15050,_w_15049,_w_15043,_w_15042,_w_15041,_w_15039,_w_15038,_w_15034,_w_15033,_w_16195,_w_15028,_w_15027,_w_15023,_w_15022,_w_16091,_w_15020,_w_15016,_w_15015,_w_15013,_w_16073,_w_15621,_w_15012,_w_15010,_w_15007,_w_15006,_w_15005,_w_15003,_w_15000,_w_14998,_w_14996,_w_14995,_w_14991,_w_15025,_w_14987,_w_14983,_w_14982,_w_14981,_w_14980,_w_14979,_w_14978,_w_14977,_w_14974,_w_14973,_w_14972,_w_14969,_w_14968,_w_14965,_w_14955,_w_14952,_w_14951,_w_14949,_w_14948,_w_14945,_w_14944,_w_14941,_w_14940,_w_14938,_w_14934,_w_14931,_w_14930,_w_14928,_w_14924,_w_14923,_w_14919,_w_14913,_w_14912,_w_14911,_w_14910,_w_14908,_w_14904,_w_14902,_w_14901,_w_14900,_w_16226,_w_14898,_w_14897,_w_14896,_w_14895,_w_14894,_w_14891,_w_14890,_w_14889,_w_14886,_w_14884,_w_14881,_w_14877,_w_14874,_w_14873,_w_14869,_w_14868,_w_14865,_w_14862,_w_14860,_w_14857,_w_14853,_w_14850,_w_14849,_w_14848,_w_14847,_w_14846,_w_14843,_w_14838,_w_14837,_w_14835,_w_15134,_w_14834,_w_14832,_w_14831,_w_14830,_w_14828,_w_15506,_w_14827,_w_14826,_w_14825,_w_14824,_w_14821,_w_14816,_w_14812,_w_14809,_w_14807,_w_14801,_w_14798,_w_14797,_w_14794,_w_14793,_w_14792,_w_14789,_w_14788,_w_14786,_w_14785,_w_14783,_w_14781,_w_14778,_w_14777,_w_14773,_w_14771,_w_14767,_w_14765,_w_14764,_w_14763,_w_14762,_w_14761,_w_14760,_w_14759,_w_14756,_w_16284,_w_16209,_w_14750,_w_14749,_w_14748,_w_14744,_w_14742,_w_16221,_w_14741,_w_14739,_w_14738,_w_14735,_w_14732,_w_14730,_w_14729,_w_14726,_w_15663,_w_14725,_w_14723,_w_14722,_w_15066,_w_14712,_w_14817,_w_14710,_w_14709,_w_14708,_w_14703,_w_14702,_w_14700,_w_14697,_w_14925,_w_14694,_w_14692,_w_14691,_w_14689,_w_14688,_w_14684,_w_14683,_w_14682,_w_14681,_w_15300,_w_15030,_w_14680,_w_14678,_w_14676,_w_14671,_w_14670,_w_14669,_w_14668,_w_14667,_w_14665,_w_14664,_w_14662,_w_14660,_w_14657,_w_15980,_w_14656,_w_14655,_w_14654,_w_14650,_w_14649,_w_14647,_w_14645,_w_14643,_w_14639,_w_14638,_w_14637,_w_14636,_w_14635,_w_14634,_w_14633,_w_14632,_w_14629,_w_14626,_w_14623,_w_14620,_w_14619,_w_14618,_w_14617,_w_14613,_w_14610,_w_14609,_w_14608,_w_14607,_w_14604,_w_14598,_w_14597,_w_14594,_w_14591,_w_14587,_w_14586,_w_15370,_w_14582,_w_14580,_w_15796,_w_14576,_w_14575,_w_14573,_w_14572,_w_14571,_w_14570,_w_14568,_w_14567,_w_14566,_w_14564,_w_15680,_w_14561,_w_14560,_w_16085,_w_14559,_w_14558,_w_14557,_w_14554,_w_14552,_w_14551,_w_14612,_w_14549,_w_15734,_w_14546,_w_14545,_w_14544,_w_14543,_w_14540,_w_14539,_w_14536,_w_14534,_w_14533,_w_14531,_w_14530,_w_14526,_w_14524,_w_16114,_w_14522,_w_14518,_w_14517,_w_14515,_w_14512,_w_14509,_w_14508,_w_14507,_w_14505,_w_14501,_w_14499,_w_14498,_w_14497,_w_14496,_w_14495,_w_14489,_w_15126,_w_14488,_w_14486,_w_14485,_w_14484,_w_14483,_w_14481,_w_14479,_w_14478,_w_14960,_w_14477,_w_14476,_w_14472,_w_14471,_w_14469,_w_14468,_w_14466,_w_14465,_w_14464,_w_15773,_w_14461,_w_14456,_w_14455,_w_15829,_w_14454,_w_14453,_w_14452,_w_14451,_w_14450,_w_14448,_w_15047,_w_14447,_w_14441,_w_14440,_w_14439,_w_14436,_w_14434,_w_14430,_w_14429,_w_14428,_w_14425,_w_14424,_w_14421,_w_14420,_w_14418,_w_14416,_w_16271,_w_16192,_w_14414,_w_15724,_w_14411,_w_14410,_w_14409,_w_14408,_w_14407,_w_14406,_w_14405,_w_14399,_w_14398,_w_14397,_w_14396,_w_14393,_w_14392,_w_14390,_w_14389,_w_14386,_w_15988,_w_14382,_w_14381,_w_14380,_w_14378,_w_14374,_w_14373,_w_14372,_w_14371,_w_14370,_w_14369,_w_14368,_w_14365,_w_14363,_w_14360,_w_14359,_w_14357,_w_14354,_w_14351,_w_14349,_w_14343,_w_14342,_w_14340,_w_15787,_w_14335,_w_14332,_w_14331,_w_14330,_w_14328,_w_14326,_w_14324,_w_14323,_w_14321,_w_14318,_w_14317,_w_14315,_w_14312,_w_14311,_w_14310,_w_14309,_w_15720,_w_14308,_w_14305,_w_14299,_w_14296,_w_14290,_w_14289,_w_14285,_w_14284,_w_14282,_w_14281,_w_14279,_w_15880,_w_14278,_w_14277,_w_14275,_w_14274,_w_14273,_w_14272,_w_14569,_w_14269,_w_14268,_w_14266,_w_14265,_w_14260,_w_14257,_w_14256,_w_14255,_w_14253,_w_14250,_w_14248,_w_14247,_w_14244,_w_14242,_w_14239,_w_14238,_w_14233,_w_14230,_w_14227,_w_14225,_w_14219,_w_14218,_w_14217,_w_14216,_w_14261,_w_14214,_w_14213,_w_14210,_w_14209,_w_14208,_w_14206,_w_14204,_w_15962,_w_14201,_w_14200,_w_14199,_w_14197,_w_14196,_w_14193,_w_14192,_w_14191,_w_14190,_w_14183,_w_14181,_w_14180,_w_14179,_w_14178,_w_14176,_w_14173,_w_14172,_w_14171,_w_14169,_w_14166,_w_14165,_w_14164,_w_14163,_w_14161,_w_14160,_w_14158,_w_14491,_w_14155,_w_14153,_w_14152,_w_14151,_w_14150,_w_14149,_w_14148,_w_14147,_w_14145,_w_14144,_w_14143,_w_14142,_w_14140,_w_14135,_w_14134,_w_14133,_w_14132,_w_14131,_w_14129,_w_14916,_w_14128,_w_14121,_w_14119,_w_14116,_w_14115,_w_14113,_w_14112,_w_14111,_w_14110,_w_14108,_w_14107,_w_14105,_w_15436,_w_14103,_w_16115,_w_14102,_w_14100,_w_14099,_w_14098,_w_14096,_w_14095,_w_14094,_w_14093,_w_14953,_w_14090,_w_14085,_w_14080,_w_14603,_w_14077,_w_14072,_w_14071,_w_14584,_w_14069,_w_14066,_w_14063,_w_14061,_w_14060,_w_14058,_w_14056,_w_14054,_w_14053,_w_14052,_w_14049,_w_14048,_w_14047,_w_14038,_w_14037,_w_14036,_w_14035,_w_14033,_w_14032,_w_14031,_w_14027,_w_15683,_w_14026,_w_14024,_w_14023,_w_14020,_w_14019,_w_14018,_w_14017,_w_14014,_w_14013,_w_14012,_w_14008,_w_14006,_w_14005,_w_16124,_w_14622,_w_14003,_w_14000,_w_13998,_w_13996,_w_13992,_w_13991,_w_13990,_w_13987,_w_13986,_w_13985,_w_13984,_w_13975,_w_13974,_w_13973,_w_13971,_w_15185,_w_13967,_w_13965,_w_13964,_w_13963,_w_13960,_w_13959,_w_13958,_w_14646,_w_13957,_w_16026,_w_15325,_w_13955,_w_13954,_w_13953,_w_13952,_w_13951,_w_13947,_w_13946,_w_15358,_w_13945,_w_13944,_w_13943,_w_13942,_w_13936,_w_13930,_w_13928,_w_13927,_w_15505,_w_13926,_w_13925,_w_13922,_w_13921,_w_13920,_w_13919,_w_13909,_w_13908,_w_13907,_w_13906,_w_13905,_w_14858,_w_13904,_w_13899,_w_15360,_w_13898,_w_15770,_w_13896,_w_16046,_w_13893,_w_15524,_w_13890,_w_13889,_w_14458,_w_13888,_w_14384,_w_13887,_w_13884,_w_13883,_w_13877,_w_13876,_w_13875,_w_13874,_w_13873,_w_13872,_w_13871,_w_13866,_w_13863,_w_13862,_w_13861,_w_13860,_w_13859,_w_13856,_w_13854,_w_13852,_w_13849,_w_13847,_w_13844,_w_13843,_w_13842,_w_13840,_w_13839,_w_13838,_w_13836,_w_13835,_w_13833,_w_13832,_w_13831,_w_13830,_w_13829,_w_13827,_w_13826,_w_13823,_w_13822,_w_13819,_w_13815,_w_13813,_w_13808,_w_13806,_w_13804,_w_13803,_w_13796,_w_13795,_w_13791,_w_13786,_w_13785,_w_13784,_w_16103,_w_13777,_w_13775,_w_15341,_w_13773,_w_13772,_w_13770,_w_13768,_w_13767,_w_13766,_w_14659,_w_13764,_w_13761,_w_13759,_w_13756,_w_13755,_w_13754,_w_13753,_w_16037,_w_13752,_w_13747,_w_13745,_w_13744,_w_13743,_w_13794,_w_13742,_w_13740,_w_13799,_w_13739,_w_13738,_w_13736,_w_13735,_w_13733,_w_13732,_w_13729,_w_13728,_w_13721,_w_13720,_w_13716,_w_13715,_w_13713,_w_13712,_w_13711,_w_13710,_w_15675,_w_13705,_w_13704,_w_13703,_w_13701,_w_15667,_w_13700,_w_13698,_w_13696,_w_14125,_w_13695,_w_13691,_w_13689,_w_13687,_w_14743,_w_13685,_w_13682,_w_13681,_w_13678,_w_13677,_w_13676,_w_13674,_w_13673,_w_13672,_w_15993,_w_13671,_w_13669,_w_13667,_w_13665,_w_13664,_w_13663,_w_13661,_w_13658,_w_13657,_w_13655,_w_13654,_w_13652,_w_13650,_w_13649,_w_13648,_w_13646,_w_13645,_w_13643,_w_13641,_w_13640,_w_13639,_w_13636,_w_13635,_w_13634,_w_13633,_w_13630,_w_13629,_w_13628,_w_13627,_w_15296,_w_13626,_w_13820,_w_13623,_w_13622,_w_13620,_w_13619,_w_13618,_w_13616,_w_13615,_w_13613,_w_13612,_w_13611,_w_14078,_w_13608,_w_13607,_w_13606,_w_13605,_w_13604,_w_13602,_w_13601,_w_13599,_w_13597,_w_15685,_w_13596,_w_13595,_w_14755,_w_13592,_w_13591,_w_13590,_w_13586,_w_13585,_w_13583,_w_13582,_w_13580,_w_13579,_w_13578,_w_13577,_w_13574,_w_13573,_w_13572,_w_13571,_w_13570,_w_13567,_w_13566,_w_15212,_w_13564,_w_13563,_w_13562,_w_14907,_w_13561,_w_13559,_w_13558,_w_13557,_w_13556,_w_15114,_w_13553,_w_13551,_w_13547,_w_13545,_w_13543,_w_13542,_w_13539,_w_13538,_w_13535,_w_13533,_w_13532,_w_14839,_w_13530,_w_13529,_w_13528,_w_13526,_w_13525,_w_16217,_w_13997,_w_13524,_w_13521,_w_13520,_w_13519,_w_13517,_w_13516,_w_14387,_w_13511,_w_13509,_w_13506,_w_13505,_w_13503,_w_15911,_w_13502,_w_13501,_w_13500,_w_15952,_w_13497,_w_13496,_w_13495,_w_13494,_w_13493,_w_13492,_w_13486,_w_13485,_w_13484,_w_13480,_w_13478,_w_13477,_w_13475,_w_13471,_w_13470,_w_13464,_w_13463,_w_13461,_w_13458,_w_13457,_w_13456,_w_13455,_w_13450,_w_13449,_w_13445,_w_13444,_w_13442,_w_15900,_w_13441,_w_13439,_w_13435,_w_13432,_w_13428,_w_13425,_w_13424,_w_13423,_w_13421,_w_13420,_w_13419,_w_13418,_w_15909,_w_13417,_w_13413,_w_13479,_w_13411,_w_13410,_w_13409,_w_15879,_w_13408,_w_13406,_w_13405,_w_13404,_w_13402,_w_13401,_w_13400,_w_13399,_w_13398,_w_13397,_w_13394,_w_13392,_w_13391,_w_14040,_w_13390,_w_13387,_w_13386,_w_13378,_w_13377,_w_13374,_w_13372,_w_13370,_w_13365,_w_13362,_w_13361,_w_13360,_w_13359,_w_13356,_w_13354,_w_14880,_w_13351,_w_13350,_w_13349,_w_13348,_w_13345,_w_13340,_w_13339,_w_13338,_w_13336,_w_13332,_w_13331,_w_13330,_w_13328,_w_13324,_w_13321,_w_13320,_w_13319,_w_13950,_w_13318,_w_13317,_w_13316,_w_13311,_w_13307,_w_13306,_w_13305,_w_13301,_w_15595,_w_13300,_w_13299,_w_15859,_w_14055,_w_13296,_w_13294,_w_13293,_w_13292,_w_13291,_w_13287,_w_13284,_w_13283,_w_15767,_w_13282,_w_13281,_w_13279,_w_13273,_w_13662,_w_13272,_w_13269,_w_13267,_w_13266,_w_13265,_w_13261,_w_13260,_w_15930,_w_13259,_w_13256,_w_14927,_w_13252,_w_13251,_w_13249,_w_13247,_w_13243,_w_13242,_w_13240,_w_13238,_w_13232,_w_13229,_w_13227,_w_13225,_w_15528,_w_13223,_w_13222,_w_13217,_w_13389,_w_13215,_w_13213,_w_13212,_w_13209,_w_13207,_w_13204,_w_13203,_w_13202,_w_13200,_w_13198,_w_13196,_w_13193,_w_13185,_w_13183,_w_13182,_w_13181,_w_13178,_w_13177,_w_14235,_w_13176,_w_15087,_w_13175,_w_13970,_w_13174,_w_13172,_w_13171,_w_13165,_w_13161,_w_13160,_w_13159,_w_13155,_w_13153,_w_13152,_w_13151,_w_15559,_w_13149,_w_13148,_w_13147,_w_13145,_w_13140,_w_13139,_w_13138,_w_13137,_w_13136,_w_13135,_w_13132,_w_13131,_w_13129,_w_13128,_w_13124,_w_13123,_w_13122,_w_13120,_w_13119,_w_15112,_w_13117,_w_13116,_w_13112,_w_13110,_w_13108,_w_13107,_w_13105,_w_13102,_w_13101,_w_13099,_w_13098,_w_13097,_w_13094,_w_15182,_w_13093,_w_15321,_w_13092,_w_16028,_w_13088,_w_13087,_w_13086,_w_13084,_w_13083,_w_13077,_w_15409,_w_13076,_w_13075,_w_13071,_w_13069,_w_13066,_w_13064,_w_13061,_w_13059,_w_13058,_w_13089,_w_13054,_w_13050,_w_13048,_w_13047,_w_13043,_w_15700,_w_13038,_w_13037,_w_13033,_w_13032,_w_13027,_w_13025,_w_13024,_w_13019,_w_13018,_w_13314,_w_13017,_w_13016,_w_13015,_w_13013,_w_13011,_w_14075,_w_13653,_w_13008,_w_13581,_w_13007,_w_14769,_w_13005,_w_13002,_w_13001,_w_13000,_w_12997,_w_15750,_w_12996,_w_12995,_w_12992,_w_12991,_w_12989,_w_12988,_w_12987,_w_12986,_w_12984,_w_15892,_w_12983,_w_15036,_w_14295,_w_12982,_w_12981,_w_13383,_w_12976,_w_12974,_w_12972,_w_12971,_w_12969,_w_14768,_w_12967,_w_12960,_w_12959,_w_12956,_w_15328,_w_12951,_w_12950,_w_12949,_w_12948,_w_12947,_w_12946,_w_15004,_w_12944,_w_12940,_w_12938,_w_12933,_w_13624,_w_12931,_w_12930,_w_12928,_w_12927,_w_12926,_w_14802,_w_12925,_w_12923,_w_12922,_w_12921,_w_12920,_w_15051,_w_12918,_w_12917,_w_12915,_w_12914,_w_12913,_w_12912,_w_12910,_w_12909,_w_12908,_w_12907,_w_12906,_w_12905,_w_12903,_w_12902,_w_12900,_w_12898,_w_12897,_w_12894,_w_12893,_w_12892,_w_16239,_w_12891,_w_14993,_w_12889,_w_12886,_w_12885,_w_12884,_w_12883,_w_12882,_w_12879,_w_12878,_w_12877,_w_12876,_w_12875,_w_12873,_w_12872,_w_12871,_w_12965,_w_12868,_w_12866,_w_12865,_w_12863,_w_12862,_w_12861,_w_12860,_w_12854,_w_12853,_w_12852,_w_12850,_w_12849,_w_12845,_w_12844,_w_12842,_w_12840,_w_14715,_w_12838,_w_15852,_w_12837,_w_12833,_w_12832,_w_12831,_w_12829,_w_12828,_w_12825,_w_12824,_w_12823,_w_15579,_w_12821,_w_12820,_w_12818,_w_12817,_w_12835,_w_12816,_w_12815,_w_12812,_w_12809,_w_12806,_w_12804,_w_12802,_w_12799,_w_12797,_w_12796,_w_12795,_w_12792,_w_12791,_w_13157,_w_12790,_w_12787,_w_12786,_w_12785,_w_12782,_w_12780,_w_13885,_w_12779,_w_12778,_w_12775,_w_12773,_w_12770,_w_12769,_w_12767,_w_12766,_w_15243,_w_12760,_w_12754,_w_12750,_w_12746,_w_15861,_w_14412,_w_12745,_w_12743,_w_12739,_w_12738,_w_12735,_w_12734,_w_12732,_w_16021,_w_12730,_w_12726,_w_12725,_w_12723,_w_12718,_w_12716,_w_12715,_w_12712,_w_12711,_w_12710,_w_12709,_w_15887,_w_12708,_w_12707,_w_12706,_w_12705,_w_12703,_w_12702,_w_12698,_w_12697,_w_12696,_w_13205,_w_12695,_w_12694,_w_12691,_w_15809,_w_13286,_w_12690,_w_12687,_w_12683,_w_12681,_w_12680,_w_12675,_w_12674,_w_12673,_w_12672,_w_12667,_w_12665,_w_12664,_w_12663,_w_12660,_w_12658,_w_12656,_w_12654,_w_12652,_w_12650,_w_12649,_w_12648,_w_12646,_w_12645,_w_12642,_w_12641,_w_14353,_w_13385,_w_12637,_w_12911,_w_12636,_w_12634,_w_12633,_w_12632,_w_12631,_w_12628,_w_12627,_w_15634,_w_12623,_w_12620,_w_12616,_w_12615,_w_12613,_w_12612,_w_14084,_w_12610,_w_12608,_w_12607,_w_12606,_w_12604,_w_12603,_w_13778,_w_12600,_w_12595,_w_12594,_w_12593,_w_16166,_w_12591,_w_12590,_w_14123,_w_12589,_w_12588,_w_13541,_w_12587,_w_12585,_w_12582,_w_12581,_w_12574,_w_12573,_w_12572,_w_12570,_w_12568,_w_12567,_w_13034,_w_12566,_w_12564,_w_14852,_w_12563,_w_12560,_w_12559,_w_12558,_w_12557,_w_14752,_w_12555,_w_12553,_w_12550,_w_12549,_w_15647,_w_12548,_w_12546,_w_12544,_w_14195,_w_12543,_w_12542,_w_12541,_w_12540,_w_12537,_w_12533,_w_12532,_w_12531,_w_12529,_w_12528,_w_12527,_w_12526,_w_12522,_w_12519,_w_12518,_w_12517,_w_12514,_w_13322,_w_12513,_w_15235,_w_13749,_w_12512,_w_12511,_w_12509,_w_12507,_w_14287,_w_12504,_w_12502,_w_12499,_w_12497,_w_12496,_w_12495,_w_16112,_w_12492,_w_12491,_w_12490,_w_12486,_w_12484,_w_12483,_w_15118,_w_12482,_w_12480,_w_12479,_w_12477,_w_12476,_w_12474,_w_12473,_w_12472,_w_12471,_w_12468,_w_12466,_w_15381,_w_12464,_w_12463,_w_12462,_w_12460,_w_12456,_w_12455,_w_12453,_w_12452,_w_12450,_w_12448,_w_12447,_w_12444,_w_12441,_w_12438,_w_12437,_w_12436,_w_12435,_w_12434,_w_13056,_w_12431,_w_12428,_w_12426,_w_12425,_w_12424,_w_12423,_w_12422,_w_12421,_w_12420,_w_12419,_w_12417,_w_12416,_w_12414,_w_12412,_w_12409,_w_12408,_w_14663,_w_12407,_w_12406,_w_16254,_w_12404,_w_12403,_w_12400,_w_12399,_w_12398,_w_12396,_w_12394,_w_15811,_w_12391,_w_12389,_w_12388,_w_12387,_w_12383,_w_15950,_w_12382,_w_12378,_w_12370,_w_12367,_w_12366,_w_15836,_w_12364,_w_12363,_w_14588,_w_12362,_w_12361,_w_12360,_w_12359,_w_12357,_w_12356,_w_12355,_w_12352,_w_12350,_w_12348,_w_12346,_w_12345,_w_12344,_w_12336,_w_12334,_w_12332,_w_15850,_w_12329,_w_12326,_w_12552,_w_12325,_w_12322,_w_12320,_w_12319,_w_12316,_w_12314,_w_12311,_w_12310,_w_12309,_w_12308,_w_12307,_w_12305,_w_12304,_w_12880,_w_12301,_w_12300,_w_12296,_w_12295,_w_14137,_w_12293,_w_12292,_w_12290,_w_12289,_w_12288,_w_12287,_w_12286,_w_12284,_w_12283,_w_12282,_w_13029,_w_12281,_w_12280,_w_12279,_w_16043,_w_12278,_w_12275,_w_12272,_w_12271,_w_12269,_w_12267,_w_12265,_w_12264,_w_12262,_w_12260,_w_12259,_w_12256,_w_12255,_w_12251,_w_12249,_w_12248,_w_12247,_w_15132,_w_14707,_w_14043,_w_12244,_w_15071,_w_12242,_w_12238,_w_12235,_w_14044,_w_12233,_w_12232,_w_12230,_w_12229,_w_12227,_w_12225,_w_12223,_w_12221,_w_12219,_w_12218,_w_12217,_w_14301,_w_12216,_w_12215,_w_12214,_w_12213,_w_12212,_w_12211,_w_12210,_w_12207,_w_12204,_w_13368,_w_12199,_w_15495,_w_12197,_w_12195,_w_12194,_w_12191,_w_12190,_w_12189,_w_12187,_w_12186,_w_15361,_w_14537,_w_12184,_w_12181,_w_12180,_w_12179,_w_12178,_w_12177,_w_12175,_w_12173,_w_12172,_w_12789,_w_12171,_w_12170,_w_12169,_w_13210,_w_12168,_w_12167,_w_12166,_w_12165,_w_12161,_w_15587,_w_12158,_w_12157,_w_12156,_w_12758,_w_12153,_w_12152,_w_12149,_w_12148,_w_12147,_w_12145,_w_12144,_w_12143,_w_12142,_w_12141,_w_12136,_w_12135,_w_12133,_w_12131,_w_12129,_w_12122,_w_14177,_w_12121,_w_12119,_w_12118,_w_12116,_w_12115,_w_13587,_w_12114,_w_15251,_w_12112,_w_12111,_w_12110,_w_12109,_w_12105,_w_12103,_w_12102,_w_12101,_w_12100,_w_12099,_w_14400,_w_12098,_w_12097,_w_12096,_w_12094,_w_15075,_w_12093,_w_12090,_w_12088,_w_12085,_w_12084,_w_15606,_w_12083,_w_12079,_w_12078,_w_13289,_w_12076,_w_12073,_w_12072,_w_12071,_w_12068,_w_12067,_w_12066,_w_12065,_w_12064,_w_12063,_w_12061,_w_12137,_w_12059,_w_12057,_w_12056,_w_12053,_w_12052,_w_12051,_w_12050,_w_12048,_w_12044,_w_16062,_w_12042,_w_12040,_w_12039,_w_12038,_w_12037,_w_12036,_w_12035,_w_12034,_w_12033,_w_12032,_w_12031,_w_12030,_w_12029,_w_12028,_w_12026,_w_15678,_w_12021,_w_12020,_w_12019,_w_12018,_w_12014,_w_12013,_w_12009,_w_13741,_w_12007,_w_12005,_w_11999,_w_14988,_w_12377,_w_11998,_w_11995,_w_11994,_w_13790,_w_11993,_w_11992,_w_11991,_w_11989,_w_11988,_w_11987,_w_11986,_w_11985,_w_11981,_w_11980,_w_11975,_w_11974,_w_11971,_w_11970,_w_13916,_w_11969,_w_11966,_w_11965,_w_11964,_w_11963,_w_11962,_w_11961,_w_11960,_w_12800,_w_11958,_w_16170,_w_11956,_w_14863,_w_11951,_w_14870,_w_11950,_w_11949,_w_11948,_w_15322,_w_11946,_w_11945,_w_11942,_w_11941,_w_11940,_w_11938,_w_11937,_w_11936,_w_11934,_w_11932,_w_11931,_w_11930,_w_11927,_w_15520,_w_11926,_w_11925,_w_11921,_w_11920,_w_11918,_w_11917,_w_11915,_w_11906,_w_11905,_w_11904,_w_11902,_w_11901,_w_11900,_w_11898,_w_11897,_w_11896,_w_11895,_w_11892,_w_11891,_w_11890,_w_11887,_w_11886,_w_11885,_w_13758,_w_11884,_w_11883,_w_11881,_w_11879,_w_11876,_w_11875,_w_11873,_w_11872,_w_11871,_w_11870,_w_14795,_w_11869,_w_11866,_w_11865,_w_11864,_w_11863,_w_11860,_w_15732,_w_11858,_w_11855,_w_11854,_w_15372,_w_11853,_w_11852,_w_15575,_w_11851,_w_11850,_w_11849,_w_12503,_w_11846,_w_11845,_w_11843,_w_11842,_w_11841,_w_11837,_w_11836,_w_11832,_w_11828,_w_11827,_w_12082,_w_11824,_w_15522,_w_11822,_w_11818,_w_13917,_w_11817,_w_11816,_w_11815,_w_11814,_w_11983,_w_11813,_w_13126,_w_11812,_w_11811,_w_11810,_w_11808,_w_11807,_w_11806,_w_11803,_w_11799,_w_11798,_w_13459,_w_11797,_w_13933,_w_11796,_w_11795,_w_11792,_w_11791,_w_11789,_w_11788,_w_11786,_w_14338,_w_11783,_w_14630,_w_11782,_w_11781,_w_11780,_w_11775,_w_12120,_w_11770,_w_11769,_w_11768,_w_16083,_w_11766,_w_13258,_w_11765,_w_11763,_w_14460,_w_11760,_w_11759,_w_11758,_w_15656,_w_11756,_w_11755,_w_11754,_w_15701,_w_15515,_w_11750,_w_11749,_w_11741,_w_11739,_w_11736,_w_11735,_w_11734,_w_11731,_w_11730,_w_11728,_w_11726,_w_11725,_w_11723,_w_11722,_w_11721,_w_11720,_w_11718,_w_11716,_w_11714,_w_11713,_w_15024,_w_11710,_w_13979,_w_11709,_w_11708,_w_11706,_w_11705,_w_11704,_w_11702,_w_11701,_w_11700,_w_11696,_w_11695,_w_11694,_w_15947,_w_11691,_w_11689,_w_11687,_w_11683,_w_14803,_w_11682,_w_11681,_w_11773,_w_11678,_w_11675,_w_11674,_w_11671,_w_11670,_w_11668,_w_11667,_w_11666,_w_11665,_w_11663,_w_11662,_w_14377,_w_11660,_w_11829,_w_11657,_w_11656,_w_11654,_w_11652,_w_11651,_w_11648,_w_11647,_w_11644,_w_11643,_w_11642,_w_11639,_w_11638,_w_11637,_w_11635,_w_15336,_w_11633,_w_11632,_w_12888,_w_11629,_w_11626,_w_11623,_w_11622,_w_11621,_w_11620,_w_11619,_w_11990,_w_11617,_w_11616,_w_11615,_w_11614,_w_11613,_w_11612,_w_11610,_w_12580,_w_11609,_w_11608,_w_14964,_w_11605,_w_11604,_w_11601,_w_11599,_w_11598,_w_11597,_w_11595,_w_11594,_w_15264,_w_14510,_w_11592,_w_11591,_w_11589,_w_11588,_w_11587,_w_11583,_w_11581,_w_11580,_w_11579,_w_11577,_w_11574,_w_11573,_w_11572,_w_11571,_w_11570,_w_11569,_w_11567,_w_11566,_w_11563,_w_11561,_w_16081,_w_11560,_w_14875,_w_11558,_w_13233,_w_11557,_w_11556,_w_11555,_w_11554,_w_11552,_w_11551,_w_13621,_w_11550,_w_13447,_w_11772,_w_11549,_w_11545,_w_14490,_w_11544,_w_11541,_w_11540,_w_11539,_w_11538,_w_11537,_w_11534,_w_13750,_w_11532,_w_11530,_w_11527,_w_11526,_w_11525,_w_12331,_w_11524,_w_11523,_w_11520,_w_11519,_w_11518,_w_11517,_w_11516,_w_15996,_w_11511,_w_11503,_w_11502,_w_15837,_w_11501,_w_11500,_w_11499,_w_11498,_w_11496,_w_13253,_w_11495,_w_11494,_w_11490,_w_11489,_w_11487,_w_11559,_w_11486,_w_11484,_w_11478,_w_14391,_w_11477,_w_12973,_w_11476,_w_11471,_w_11470,_w_11467,_w_11466,_w_11465,_w_11464,_w_11463,_w_11462,_w_11461,_w_14621,_w_11458,_w_11457,_w_11454,_w_11453,_w_11452,_w_11450,_w_11449,_w_15350,_w_11444,_w_11443,_w_13792,_w_11441,_w_11438,_w_11437,_w_11436,_w_11435,_w_11434,_w_14404,_w_11432,_w_11431,_w_11429,_w_11428,_w_11427,_w_11426,_w_11425,_w_11424,_w_11423,_w_12202,_w_11422,_w_11421,_w_11419,_w_11416,_w_11414,_w_11893,_w_11413,_w_11406,_w_11405,_w_11403,_w_11401,_w_11399,_w_15146,_w_11398,_w_11397,_w_11394,_w_11393,_w_11390,_w_12443,_w_11387,_w_11386,_w_11385,_w_11384,_w_11383,_w_14800,_w_11380,_w_13600,_w_11378,_w_11377,_w_11376,_w_12662,_w_11373,_w_11372,_w_14985,_w_11369,_w_11368,_w_14842,_w_11522,_w_11365,_w_11364,_w_11363,_w_11362,_w_11361,_w_11360,_w_11359,_w_11357,_w_13290,_w_11356,_w_11353,_w_11352,_w_11351,_w_11349,_w_11536,_w_11347,_w_11345,_w_11342,_w_11341,_w_11339,_w_11338,_w_11337,_w_11335,_w_11334,_w_11333,_w_11331,_w_11330,_w_11327,_w_11326,_w_15391,_w_11325,_w_11323,_w_11321,_w_11319,_w_11318,_w_11315,_w_11313,_w_11311,_w_11309,_w_11308,_w_15424,_w_11839,_w_11305,_w_11304,_w_11302,_w_11300,_w_11297,_w_15037,_w_11295,_w_11292,_w_11547,_w_11291,_w_11290,_w_11289,_w_11287,_w_11285,_w_11284,_w_11283,_w_11282,_w_11280,_w_11279,_w_14467,_w_13162,_w_11277,_w_11757,_w_11276,_w_11275,_w_11273,_w_11272,_w_11270,_w_11268,_w_11266,_w_11260,_w_11259,_w_11258,_w_15896,_w_11257,_w_11256,_w_11719,_w_11255,_w_11254,_w_11253,_w_11252,_w_11251,_w_11388,_w_11248,_w_11247,_w_11244,_w_11241,_w_11237,_w_11235,_w_11233,_w_11479,_w_11232,_w_11230,_w_11229,_w_11228,_w_14139,_w_11226,_w_11223,_w_11222,_w_11221,_w_12150,_w_11219,_w_11217,_w_11216,_w_11214,_w_11213,_w_15382,_w_11212,_w_11210,_w_11209,_w_11207,_w_11206,_w_11204,_w_11202,_w_11201,_w_11200,_w_11199,_w_14779,_w_11198,_w_11197,_w_11195,_w_11194,_w_11192,_w_11191,_w_11190,_w_11189,_w_11187,_w_11185,_w_11183,_w_11181,_w_11178,_w_12859,_w_11177,_w_11515,_w_11173,_w_13074,_w_11172,_w_11168,_w_11166,_w_11164,_w_11417,_w_11163,_w_11161,_w_11160,_w_11159,_w_11158,_w_11157,_w_11156,_w_11155,_w_11153,_w_11151,_w_11149,_w_11148,_w_12763,_w_11147,_w_11145,_w_11143,_w_11142,_w_11141,_w_11139,_w_11137,_w_11134,_w_11132,_w_11131,_w_11130,_w_11129,_w_11127,_w_11125,_w_11123,_w_13395,_w_11122,_w_11121,_w_11119,_w_11117,_w_11116,_w_11115,_w_11110,_w_11109,_w_16006,_w_15248,_w_11107,_w_11105,_w_11104,_w_11102,_w_11098,_w_11096,_w_11095,_w_11094,_w_11091,_w_11090,_w_11089,_w_11088,_w_15693,_w_11087,_w_15008,_w_11080,_w_16183,_w_11079,_w_11077,_w_11075,_w_11074,_w_12055,_w_11073,_w_11072,_w_11070,_w_11069,_w_11068,_w_12478,_w_11066,_w_11065,_w_11064,_w_12298,_w_11061,_w_11057,_w_11056,_w_11054,_w_11053,_w_11052,_w_14699,_w_12222,_w_11051,_w_11048,_w_11047,_w_15538,_w_11046,_w_11475,_w_11045,_w_11044,_w_11042,_w_11039,_w_11844,_w_11036,_w_11034,_w_14130,_w_11032,_w_11038,_w_11031,_w_11029,_w_11028,_w_12554,_w_11027,_w_15340,_w_11025,_w_11023,_w_11022,_w_11021,_w_15295,_w_11020,_w_11019,_w_11018,_w_11017,_w_11016,_w_11014,_w_11013,_w_11011,_w_11086,_w_11010,_w_11008,_w_11007,_w_11006,_w_11005,_w_11004,_w_11003,_w_10999,_w_10998,_w_11692,_w_10997,_w_12736,_w_10996,_w_13430,_w_10991,_w_10989,_w_10988,_w_10986,_w_10984,_w_10983,_w_10982,_w_10981,_w_10980,_w_10978,_w_14882,_w_10977,_w_13679,_w_10976,_w_10975,_w_10973,_w_10970,_w_11188,_w_10969,_w_10968,_w_10965,_w_10964,_w_10963,_w_10961,_w_10960,_w_10959,_w_10957,_w_14766,_w_10956,_w_10955,_w_10954,_w_10953,_w_10950,_w_10948,_w_10944,_w_13144,_w_10943,_w_10942,_w_13552,_w_10941,_w_10940,_w_10939,_w_10937,_w_10936,_w_15934,_w_10935,_w_11618,_w_10933,_w_10932,_w_11348,_w_10931,_w_10928,_w_10927,_w_10924,_w_10923,_w_15413,_w_10922,_w_10920,_w_10917,_w_10916,_w_10911,_w_10910,_w_10909,_w_13431,_w_10906,_w_10903,_w_15234,_w_10901,_w_10897,_w_10896,_w_16012,_w_11381,_w_10895,_w_10894,_w_10893,_w_10892,_w_10890,_w_10888,_w_10886,_w_14480,_w_10885,_w_11389,_w_10882,_w_10881,_w_10880,_w_10879,_w_10876,_w_10873,_w_10871,_w_11973,_w_10870,_w_10866,_w_10865,_w_10863,_w_15908,_w_14675,_w_13376,_w_10862,_w_10861,_w_14221,_w_10859,_w_10857,_w_10856,_w_10854,_w_11856,_w_10853,_w_14961,_w_10849,_w_10845,_w_10843,_w_10842,_w_12644,_w_10841,_w_10839,_w_10838,_w_10835,_w_10833,_w_10832,_w_10831,_w_16261,_w_13845,_w_10829,_w_10824,_w_10820,_w_16174,_w_10819,_w_15633,_w_10817,_w_10858,_w_10816,_w_10815,_w_10814,_w_10813,_w_12813,_w_10812,_w_10811,_w_10809,_w_10808,_w_11627,_w_10972,_w_10806,_w_10802,_w_10801,_w_10800,_w_10797,_w_10796,_w_12668,_w_10795,_w_10793,_w_10790,_w_14909,_w_10786,_w_10785,_w_10782,_w_12127,_w_10780,_w_10779,_w_10778,_w_10777,_w_10776,_w_10775,_w_10773,_w_10772,_w_15068,_w_10771,_w_10769,_w_11224,_w_10766,_w_10764,_w_10763,_w_10762,_w_10760,_w_10759,_w_10757,_w_10756,_w_10754,_w_15009,_w_10752,_w_10751,_w_13568,_w_10749,_w_16264,_w_10747,_w_10746,_w_10742,_w_11261,_w_10740,_w_10739,_w_10737,_w_13780,_w_10736,_w_10734,_w_10732,_w_10729,_w_11778,_w_10728,_w_10727,_w_10725,_w_10723,_w_10722,_w_10719,_w_10718,_w_10716,_w_13995,_w_10715,_w_10714,_w_10713,_w_10712,_w_10710,_w_10708,_w_10704,_w_10703,_w_10702,_w_10701,_w_10700,_w_10699,_w_10698,_w_10695,_w_14459,_w_10693,_w_14188,_w_10692,_w_10689,_w_10688,_w_12001,_w_10687,_w_10686,_w_10685,_w_10684,_w_10683,_w_10682,_w_10681,_w_12245,_w_10679,_w_10678,_w_10674,_w_10673,_w_10672,_w_10671,_w_15312,_w_10670,_w_10669,_w_12505,_w_10668,_w_10667,_w_10666,_w_10694,_w_10663,_w_10661,_w_10659,_w_10657,_w_12390,_w_10654,_w_10653,_w_10652,_w_10650,_w_10649,_w_10646,_w_11584,_w_10645,_w_10643,_w_10642,_w_10638,_w_10637,_w_15485,_w_10629,_w_10626,_w_10625,_w_10624,_w_10620,_w_10619,_w_10617,_w_10612,_w_10611,_w_10609,_w_10607,_w_10605,_w_15142,_w_10604,_w_10601,_w_10598,_w_10597,_w_11602,_w_10595,_w_15384,_w_10593,_w_10591,_w_10587,_w_13028,_w_10586,_w_13065,_w_10584,_w_16251,_w_10583,_w_10582,_w_10741,_w_10581,_w_10580,_w_10579,_w_10578,_w_12881,_w_10577,_w_10574,_w_12410,_w_10573,_w_10572,_w_13403,_w_10571,_w_10570,_w_10565,_w_10564,_w_14519,_w_10563,_w_10562,_w_10561,_w_10560,_w_10558,_w_10557,_w_12764,_w_10555,_w_10553,_w_10552,_w_14118,_w_10550,_w_11774,_w_10548,_w_10545,_w_10544,_w_10543,_w_10541,_w_10540,_w_10538,_w_10537,_w_10535,_w_10534,_w_10533,_w_10532,_w_10531,_w_10530,_w_10525,_w_10523,_w_10522,_w_10519,_w_10518,_w_10516,_w_10515,_w_13527,_w_10966,_w_10514,_w_10512,_w_10510,_w_10508,_w_10505,_w_11358,_w_10504,_w_10503,_w_10502,_w_16169,_w_10501,_w_10499,_w_10498,_w_14625,_w_10497,_w_10495,_w_10492,_w_10491,_w_10490,_w_10489,_w_10488,_w_10487,_w_10486,_w_15616,_w_13130,_w_11293,_w_10483,_w_10482,_w_10477,_w_10475,_w_12228,_w_10474,_w_10473,_w_15288,_w_12626,_w_10470,_w_12597,_w_10469,_w_10468,_w_10467,_w_11332,_w_10464,_w_10463,_w_10461,_w_10457,_w_10455,_w_10453,_w_10452,_w_14236,_w_10450,_w_15786,_w_10449,_w_10447,_w_10636,_w_10445,_w_10443,_w_10441,_w_10440,_w_10439,_w_10438,_w_15215,_w_11699,_w_10437,_w_10434,_w_14698,_w_10432,_w_10430,_w_11354,_w_10427,_w_10426,_w_10424,_w_10423,_w_10421,_w_10420,_w_10416,_w_10415,_w_15150,_w_11888,_w_10414,_w_11679,_w_10413,_w_12576,_w_10412,_w_10411,_w_10410,_w_10409,_w_10406,_w_11676,_w_10405,_w_10403,_w_10402,_w_10401,_w_10400,_w_10399,_w_10398,_w_12935,_w_11953,_w_10396,_w_10395,_w_13326,_w_13295,_w_10394,_w_10392,_w_10390,_w_10389,_w_10705,_w_10387,_w_10381,_w_10380,_w_12347,_w_10378,_w_10377,_w_10375,_w_10720,_w_10372,_w_10371,_w_11497,_w_10369,_w_10368,_w_14504,_w_10364,_w_11298,_w_10363,_w_10361,_w_10359,_w_10357,_w_10356,_w_11507,_w_10354,_w_10352,_w_10351,_w_10664,_w_10349,_w_10348,_w_10347,_w_10341,_w_10339,_w_10337,_w_10333,_w_10331,_w_14433,_w_10328,_w_10327,_w_10326,_w_10323,_w_10321,_w_10320,_w_10319,_w_16030,_w_10448,_w_10318,_w_10317,_w_10316,_w_10315,_w_10314,_w_15040,_w_10311,_w_14578,_w_10310,_w_10309,_w_10307,_w_10305,_w_10303,_w_14592,_w_10302,_w_11903,_w_10301,_w_16016,_w_10297,_w_13730,_w_10296,_w_10295,_w_10294,_w_10293,_w_10292,_w_10291,_w_10289,_w_10288,_w_10287,_w_10286,_w_10284,_w_10283,_w_10282,_w_10279,_w_10278,_w_12196,_w_10276,_w_13727,_w_10275,n954_0,N511_16,_w_6227,n946_0,_w_11727,n941_0,_w_7445,_w_13237,n1054_1,_w_8216,_w_15717,n938_0,_w_13544,n1412_1,n935_0,_w_15577,_w_12506,n1695_1,n578_1,n926_0,_w_7419,n1194_1,n1269,n947_1,n1074_1,n732_0,_w_6848,n220_1,_w_9981,n919_1,n919_0,_w_14810,_w_11761,n916_1,_w_15104,_w_12469,n825_1,_w_8261,_w_11834,n916_0,n741_0,n905_1,_w_12751,n1295,N239_18,_w_12772,N239_16,n1190,_w_9402,_w_8488,_w_12205,_w_9397,N239_11,_w_12811,n770,N239_2,N239_0,_w_15069,n1779_0,_w_14791,_w_6214,_w_7757,n884_1,_w_7845,_w_14711,_w_10651,_w_8097,n1512_1,n860_0,_w_11059,_w_5914,_w_9407,_w_5967,_w_13938,n883,_w_12006,_w_6085,n211,n1403,_w_9150,n844_1,_w_10878,n247_1,_w_9348,_w_12385,n1063_1,_w_9440,n1039_0,n829_1,_w_15997,_w_11400,n716_0,_w_10147,n816_1,_w_8332,_w_5887,n816_0,_w_13035,_w_12349,n460_0,n237_1,_w_14322,_w_9220,n1244_1,n995_0,_w_12523,N35_17,n808_1,_w_16171,n877_1,n1708,n807_0,n137_0,n804_0,n802_0,n1652_1,_w_9683,n1779_1,_w_14333,n1652_0,n1873_1,n267,_w_12285,n383,_w_12937,_w_11528,N171_15,n1631,_w_11485,_w_10913,_w_8931,_w_6144,N171_5,n238,n1523,_w_14346,_w_6485,N171_3,n1057,n1686_1,_w_15894,n1686_0,n874_1,n324_1,n1177_1,n762_0,n253_1,_w_8246,_w_7548,_w_11576,n1783_1,_w_7874,n795_1,n1533_0,n787_0,_w_15021,n527_1,n1324_1,n970,_w_15477,_w_13878,_w_7907,n805_1,n1855_0,_w_12701,_w_10907,_w_10794,n822_0,n1046_2,_w_13275,n1010_0,_w_7842,_w_15602,_w_12351,n605_1,n605_0,n1229_0,N409_8,n364_0,_w_10804,n850,n1025_0,n810_0,_w_13918,_w_6966,_w_14212,_w_11410,_w_8430,n768_1,n634_1,_w_9951,n742_1,n742_0,_w_14887,_w_10528,n1437_0,n1839_1,n1839_0,n204_1,n204_0,n1409_1,_w_8781,n729_1,n300_0,n727_0,n803,n112_1,n1468_1,_w_10904,_w_7183,n1712_0,_w_9342,_w_14283,_w_12130,n725_1,_w_7130,n722_1,_w_14159,n632,_w_8785,n820_0,n1570_0,n718_1,n718_0,n1479_0,_w_14770,_w_5635,_w_9087,n717_0,n716_1,n1310,n1841_1,n715_1,n713_1,_w_8622,n300_1,n1816,_w_12774,_w_12303,n845_0,_w_15357,_w_6491,n709_1,_w_10419,n1332_1,N171_8,_w_14859,_w_8373,n295_1,_w_11469,n1297,_w_6270,_w_13355,_w_10252,n1709_0,n1278_1,_w_13514,N137_17,_w_12822,_w_9601,n590_0,_w_5899,n688_0,_w_6498,_w_7001,n687_0,n569,n1675_1,n1675_0,_w_14550,_w_14532,n1389,_w_8540,n997_1,n826_1,n54_1,n682_1,_w_10549,n681_0,_w_6773,_w_11823,n393_1,n673_0,n144_0,n93_0,_w_15018,n669_1,_w_13304,N120_16,n1421_1,n1331,_w_15847,n998_0,N120_15,N120_14,n345_1,_w_15762,_w_6295,_w_11825,_w_10103,N120_10,n517_1,_w_16075,_w_6301,_w_9771,N120_7,_w_5641,N120_5,_w_12945,N120_3,_w_9919,N120_2,_w_11100,n655_0,_w_15630,n1336_0,n1062_1,n1468_0,n640_1,n640_0,_w_6950,n532_1,n127_1,n1633,n127_0,n628_1,n327_1,n255_0,n696_0,_w_7090,n1302_1,_w_15573,n771_1,n832_0,_w_13352,n594_1,_w_12968,_w_9749,_w_10256,_w_7481,n174,_w_16024,_w_13384,_w_5495,n913_1,n1466,n620_0,n1426,_w_15933,n817_0,n618_0,n694_1,n1772,n1864_0,_w_8447,_w_13195,n616_1,n1329_1,_w_13787,n1060_0,n1202_0,n1030_1,n588_1,n585_1,n940_1,n931_1,n931_0,n626_0,n712_1,n1566_1,n781_0,_w_6746,_w_8669,n582_0,_w_12054,n132_1,n1806_0,_w_13487,_w_10345,_w_6159,n118,_w_10163,_w_10313,n1378_1,n1378_0,n1637_1,_w_8055,_w_8475,n660_1,n997_0,_w_12720,_w_12317,n944_1,_w_12539,n306_0,n566_1,n705,_w_15513,n566_0,n835_0,n648_1,_w_10945,n911_0,n560_0,_w_5532,n1306_1,N477_5,n1306_0,n877_0,_w_9906,_w_15940,n769_1,n223_0,n356,_w_14091,_w_7147,n549_1,n708_0,_w_11415,n368_1,n1672_1,n1672_0,n1848,_w_10260,n539_1,_w_6563,n1777_1,n753,_w_7672,_w_11840,n533_0,n1109_1,_w_5859,n531_1,_w_12598,_w_11909,n153_0,n811_1,n530_1,n956_1,_w_16242,_w_11680,n232_0,n998,_w_15758,_w_5762,n475_1,n1881_1,_w_10436,n225_1,_w_7512,_w_8088,n225_0,n1025_1,_w_10733,n976_1,_w_13924,n883_1,_w_12814,_w_11150,n1537_0,_w_11805,n1075_0,n652_1,_w_7857,n652_0,_w_14258,_w_11382,_w_9251,n1142,_w_6186,n606_1,_w_11819,n535_0,_w_7446,_w_15473,n213_1,N426_19,n1004_0,n778_0,_w_5313,n66_0,n97_0,n126_0,_w_6544,n811,_w_10273,_w_8150,n955_0,n108_2,n1428_0,_w_13809,_w_9676,n581_1,_w_6653,n108_1,n201_0,_w_8311,_w_7307,_w_16061,_w_13982,_w_8722,n373_1,n373_0,_w_6032,n1049_1,n914,n1049_0,_w_8531,_w_9494,n129_1,n191_0,_w_6176,n1028_0,n137,_w_12714,_w_8590,_w_8025,n183_1,n183_0,_w_15582,n1158_0,n307_1,_w_12788,n1191_1,_w_6482,n831_1,_w_7981,n831_0,n1530_0,n272,n730_1,n1179_0,_w_11703,n490_1,n567,_w_13381,n1113_1,n276_0,n1055,_w_7029,n1826_0,n1716_0,_w_9279,_w_9628,n727_1,n138_0,N528_12,_w_12953,n1741,_w_7020,N307_9,_w_14565,n1296_1,_w_9886,N443_9,_w_7316,n658_1,_w_11002,_w_7743,_w_13187,_w_8492,_w_6621,n663_0,n396_1,n1886_0,n1344,n184_1,_w_12756,_w_10594,n184_0,_w_10028,_w_11246,n1594_0,_w_5348,_w_7355,n1024_1,_w_6972,n1024_0,N154_17,_w_9084,n384_1,n150_1,n1227_0,_w_13045,n599_0,n722_0,_w_15785,n629_1,N358_17,_w_7182,N358_16,N358_10,_w_13762,_w_6293,_w_6586,n790_0,_w_12077,_w_6263,_w_10592,_w_7571,N358_3,_w_10020,N358_0,_w_11847,N528_11,n207_1,n1638_1,_w_7805,n596_1,_w_7960,n666_0,_w_8682,n1459_1,n1037_0,_w_13199,_w_8675,n158_0,n1206_1,_w_10547,n365,_w_8593,_w_10322,n139_0,n362_1,n1606_1,n454_0,n308_0,_w_5507,_w_9714,n693_1,_w_15174,_w_10235,n1717,_w_13274,n1540,n728_1,n1560_1,_w_6021,n1560_0,n1550_0,n118_0,n1457_1,n673_1,n177_1,_w_8817,_w_15141,n145_0,n1579_0,n960_1,n133_0,_w_16048,n451_1,_w_10373,n1176_1,N52_8,N392_8,n1787_0,_w_15967,n1485_1,n1070_0,n1348_0,_w_11392,_w_10640,n1186_1,_w_5892,n784_1,_w_15261,n107_0,n420_0,n757_0,n731_0,_w_11878,_w_5513,_w_10887,n124_0,n117_1,n94_1,N222_1,n377_0,n436_1,n651_1,_w_11328,n1698,n247,n1131,_w_15095,n255_1,_w_14168,_w_8570,_w_15622,n374_0,_w_12896,n1410_1,_w_10493,n105_0,_w_13375,n65_0,_w_9864,n1065_1,_w_14716,_w_12381,n860_1,n982,n848_0,n859_1,_w_15378,_w_10675,n859_0,n869_0,n1505_0,n738_1,_w_9254,n101_1,n898_0,_w_16011,_w_13932,n1533,_w_14303,N528_19,_w_8786,n690_1,N528_15,_w_16282,_w_10480,n667_1,_w_6024,_w_10787,_w_6229,N528_9,n787,N528_8,n1679_0,_w_15239,N528_7,n1068_0,N528_5,_w_15899,n719_1,_w_5554,_w_11211,_w_8898,N528_1,_w_9838,n190_1,_w_7841,_w_14644,n190_0,_w_13869,n228_1,n964_1,n228_0,n1832,_w_7173,n1540_0,_w_15342,_w_6813,_w_15278,n141_1,n141_0,_w_13999,_w_7793,n612_1,n529,_w_15500,n45_1,n222_0,_w_11826,_w_10203,n1031,n1040_1,n256_0,_w_10616,n928_0,_w_5836,_w_14101,_w_12341,n909,n1614_1,N137_15,_w_12372,_w_5942,N137_13,_w_15029,n735_1,_w_9208,N137_11,N137_8,_w_10265,N256_18,n164_1,n385,_w_7327,_w_10662,_w_9487,n397_0,_w_14339,_w_7028,n1010_1,N154_19,_w_13250,_w_9408,n1836_1,n1641_0,N154_16,_w_14876,n822_1,_w_9571,N154_15,_w_10823,n1015,_w_10460,N154_9,n1736_0,_w_15348,n1259_1,n543_1,_w_15061,_w_10527,n942_0,_w_10081,n1780_1,n187_1,_w_6951,_w_12449,N154_1,n1781_1,_w_14079,_w_10500,n1168_0,n471_1,_w_14138,n471_0,_w_13748,n329_0,N1_19,N188_8,_w_11521,N1_16,_w_8614,_w_15290,_w_11480,_w_10431,N1_11,n483_0,n1545_1,N1_9,_w_15486,N1_8,_w_6454,_w_6896,N1_6,N1_4,_w_10462,N1_3,_w_9306,_w_16055,N1_2,_w_11249,n1217_0,n1281_0,N1_1,_w_13699,n1256,_w_8098,_w_13091,_w_7030,n1621_1,n301_1,n951_1,n990,n951_0,N460_9,n1168_1,_w_6254,n908_1,n301,n56_2,n56_0,n1837,n500,_w_9134,n904_1,n1471,_w_15936,n747_0,n1037_1,n1287_0,_w_12457,_w_9835,n679_0,n96_0,n763_1,N239_17,n958_0,_w_7318,n498_1,_w_9216,_w_10952,n1883_1,n1876_1,_w_6512,n54_0,n48_1,N324_19,_w_16045,n844_0,_w_5714,n786_0,_w_6703,n195_1,N324_11,_w_14313,N324_9,n185_0,n182_0,N324_8,N324_5,n1012_0,N324_3,N324_2,n708_1,N324_1,_w_11630,n347_0,_w_14574,n1068_1,_w_8794,n462_1,n808_0,_w_14050,n974_0,_w_13631,n1694_1,_w_15231,n1694_0,n625,_w_10755,n180_0,_w_8333,n967_0,_w_15417,_w_10958,n294,_w_13095,n587_0,N341_18,N35_16,n543_0,n540_1,n841,n566,N341_16,n1448,N1_5,_w_12629,_w_11939,_w_8857,n657_1,n1199_1,n957_0,N341_10,N341_4,n441_0,n1194_0,_w_8911,_w_12489,_w_9572,n1628_1,N341_2,_w_15001,n733_1,_w_11562,n1818,N358_6,_w_7684,_w_16145,_w_12276,n983,_w_15502,N409_14,N409_13,n1563,_w_6928,n1376_0,n621,_w_10330,N409_5,_w_13722,_w_12584,N409_3,_w_7401,_w_11944,_w_10884,_w_9593,_w_8330,n866_0,n1555,_w_12621,n192_0,n1490_1,_w_11924,_w_10753,_w_9207,_w_14714,n801_0,_w_7698,n1533_1,_w_10038,n1224_1,n634_0,N426_14,_w_5704,_w_11101,n142_0,n749,_w_11186,n792_1,n143_0,_w_12498,n397,_w_11784,N426_11,_w_12174,_w_7515,_w_8126,_w_8395,_w_9222,N341_12,n1402,n1050,_w_15694,N426_9,_w_13241,_w_8443,N426_7,_w_13666,n1293_0,N460_17,n1370_0,_w_15688,n1549_0,n936_1,_w_6588,_w_11684,_w_9566,N460_16,_w_9142,_w_15619,n1819_0,N460_7,N460_5,n1009_1,_w_13737,_w_12315,_w_8668,_w_13049,n893_1,n613_1,N205_11,_w_10848,n421_1,n432_1,_w_14446,_w_9560,N477_18,n1862,_w_5693,N477_16,n80,_w_5989,_w_6821,_w_16139,N307_2,N341_5,_w_5783,_w_7722,N358_9,N477_0,N409_9,_w_5851,_w_8729,N154_7,N511_15,_w_13989,_w_7741,N511_14,n534_0,_w_8082,_w_6870,n60_0,_w_7378,_w_11265,n538_0,_w_11913,n1588_1,n895_1,n140_0,_w_10621,n361_1,n857,n79,_w_12239,_w_5803,_w_10005,_w_6356,N528_13,n817_1,n1257,_w_6036,_w_14872,_w_5608,_w_9106,n540_0,n766_0,n820_1,n1782_0,N103_17,N103_15,_w_15465,_w_7750,_w_8460,N103_7,n648,_w_15011,_w_8616,N103_5,n1871,_w_13194,_w_11473,_w_7957,n1878_0,_w_16099,N103_2,_w_6507,_w_8830,n720_0,_w_6374,_w_12075,n1606_0,n62_1,_w_7891,n326_0,_w_12198,_w_10192,N443_18,N443_16,_w_7350,N443_15,n1821_0,n379_0,_w_10342,_w_10182,_w_13073,_w_11698,_w_6111,N443_6,n1107_1,_w_10867,_w_8438,_w_13774,n567_0,n1553,_w_5334,_w_10343,_w_5742,_w_13818,_w_13515,n1715_0,n591_0,n1440_1,n208_0,_w_10758,n69_1,n286_0,n196_1,_w_10222,n636_1,n636_0,n896,n846_1,_w_5566,_w_16272,_w_15838,n161_0,_w_11344,_w_6399,N460_12,n85_1,n841_1,_w_16173,_w_16108,n1701,_w_5557,_w_8412,n85_0,_w_6690,_w_8638,n796_1,n1188_0,_w_14939,_w_7356,n796_0,_w_9653,n236_0,n1217,n886_0,n1873,N35_18,N358_12,n622_1,n53_1,_w_6438,n1134_0,_w_6502,n304_0,N35_13,_w_10556,N35_12,_w_9544,_w_6212,n78_1,n617_1,_w_8003,_w_11346,N35_9,_w_13482,N35_7,n661_0,_w_10631,_w_8061,n49_0,n1458_0,n1136_1,_w_7104,n1494_0,n438_1,n429_1,N86_7,n923_1,n429_0,_w_16199,n569_0,n1759_1,n1759_0,n1609,N443_0,_w_13143,_w_8052,_w_8066,_w_12545,_w_8966,n1609_0,n1731_1,n470,_w_9609,_w_6069,N307_18,N545_0,n905_0,_w_7906,N307_17,_w_10851,N426_3,n670_1,_w_6852,_w_10198,_w_9635,n121_1,N307_10,n259_0,_w_14442,N528_10,N307_8,_w_14403,N307_5,_w_9312,_w_6357,_w_11911,N307_3,_w_15246,N307_1,n1165_0,_w_10551,n799_0,n285_0,n1314,_w_11111,n1622,n153_1,n155_1,n1814_1,_w_12957,_w_7140,n1785,n504_0,n394_0,n1531,n493_0,N86_19,_w_14971,_w_11136,N86_17,_w_11923,n1122,n1655_1,_w_7007,_w_10765,N86_15,N86_13,_w_9324,n246_1,_w_13052,_w_10781,n1652,_w_13230,_w_7660,_w_13219,n1507,_w_15839,n1671,_w_14226,N86_4,_w_8331,N86_3,n842_0,_w_9463,N86_0,_w_7911,n1418_1,_w_12731,n281,_w_14124,_w_11009,n773,_w_9882,n267_0,n1092,_w_7405,_w_12430,n814_1,n1689,n1372_0,n152,n427_1,_w_14231,n640,_w_16098,_w_5928,_w_6674,n1731_0,n1239_1,n333_1,n1272_0,_w_6180,n487_1,n487_0,n35_2,n35_1,n588_0,_w_14010,n874_0,_w_11374,n35_0,_w_12874,_w_12538,n1031_1,n832_1,_w_7475,n130_1,_w_5525,N426_17,n68_1,_w_7064,n1800_1,n1323_0,_w_9997,n537_0,_w_12043,n41_0,n1619_1,_w_15196,n1619_0,_w_11001,_w_6331,_w_9122,N528_0,n82_1,_w_5545,n1721_1,n82_0,n792,n1854_0,n45_0,n1150,n1767_0,n1227_1,_w_16152,_w_12521,n1485_0,n308_1,_w_14358,n882,n726_1,n461,_w_5838,_w_15614,N69_15,_w_14042,_w_7846,_w_13197,_w_6153,n484_1,_w_5844,_w_13263,N69_10,n1315,N528_6,_w_7249,N69_6,n546,_w_16101,N69_3,n1413,_w_6322,N69_1,n1345_1,n262_0,_w_9161,_w_15651,_w_11113,_w_5962,n74_0,n1497_1,n530_0,n52_1,_w_5873,_w_13523,n712_0,_w_11838,n264_1,_w_7574,_w_6827,_w_6806,_w_15213,_w_11412,_w_8208,n526_0,_w_7480,_w_7995,n621_1,n734_1,_w_13469,n734_0,n366_1,_w_15759,n521_0,n576_1,_w_8833,n576_0,N494_18,n748_1,n1196_0,_w_9291,_w_12312,n1880_0,N494_17,N494_16,_w_15783,_w_14122,n1076_1,_w_5868,n241_1,n1000_0,n140_1,N494_12,_w_13221,n875_0,N494_9,n1773_1,n664_0,_w_11451,n514_1,n72,_w_7900,n1847_0,_w_8960,n664_1,_w_6623,_w_15961,n730_0,n144_1,n520_0,n763_0,n593_1,n1543_0,n620,n614_1,_w_12857,n388_1,_w_14068,n165,N69_4,n388_0,_w_12012,n1185_0,n1273_0,n75_0,_w_12619,n260,n1739_0,_w_12379,_w_9278,n400_1,n1602,n637_1,_w_14701,n213_0,_w_6248,_w_13769,n305_0,_w_14355,_w_8069,_w_9647,n240_0,n1016_0,N222_19,N358_15,N222_18,N341_6,_w_15833,_w_15263,_w_11411,n1399,_w_5694,_w_15175,n898,N222_14,_w_9563,_w_15335,n564_0,n536,_w_5442,N222_7,_w_14293,_w_6081,N273_18,N273_15,n1209_1,n1011,N273_2,_w_6832,N273_0,n1111,N137_18,n1174_1,_w_12123,n631_1,n1646,_w_12535,n1086_1,_w_15464,N103_9,N426_8,_w_6290,_w_6511,n1086_0,n81_0,_w_14203,n602_0,_w_16253,_w_10799,_w_9259,n1861_1,_w_13731,_w_5628,n280_0,n1750_1,n1704_0,n84_1,n1409_0,_w_6198,n288_1,_w_6475,n274_0,n502_0,n456_2,_w_5426,n456_1,N290_14,N290_8,n807_1,n945_1,n1703_0,N290_5,n959_0,_w_15751,_w_8164,_w_8739,n1802_1,n1802_0,_w_13911,_w_9797,_w_11037,N375_4,_w_5862,_w_7273,n235_1,n1829_0,_w_13507,_w_10644,n843_1,_w_13452,_w_5963,n342_0,n243_1,_w_9507,_w_10074,_w_15637,_w_14696,N137_9,_w_8007,_w_12162,_w_8923,_w_13901,n1198,_w_11954,n238_0,n378_1,_w_9143,n378_0,N409_18,_w_14292,n714_0,N188_19,N188_18,_w_12080,N188_17,n1711,_w_9137,N188_16,N188_15,_w_16034,_w_15791,_w_13841,_w_11833,N188_14,N188_13,_w_7819,N188_5,_w_11124,N188_3,n246_0,_w_6460,n1491_1,_w_6745,_w_14470,n250_1,n217_1,_w_5519,n834_1,n1392,_w_10383,n403_1,n1199_0,_w_12638,n705_1,n451,n403_0,_w_7610,n252_0,n481_0,n952_1,n1248,n737_2,N205_17,N205_14,N205_13,_w_8284,n921,_w_12516,_w_9436,_w_12994,N205_12,n1376,_w_7256,N205_10,n1341_0,_w_9008,n1107_0,N205_8,_w_10912,_w_7292,N205_6,n1043,N358_8,N341_7,N205_4,n608_0,_w_12602,_w_7589,_w_9549,_w_10034,n103,N205_1,_w_8112,n258_0,n384,_w_15604,n411_0,_w_12302,n73_0,_w_14871,_w_12870,_w_6118,_w_5329,n273_0,n274_1,_w_8632,n1154_1,_w_11322,n1193,_w_7799,n344_1,n103_1,n1430_1,n1076_0,n279_1,n302_0,n872_0,n305,_w_5542,_w_13022,n282_1,_w_6650,_w_9984,n192_2,n448_1,_w_14641,_w_6393,_w_13180,_w_8370,n579_0,n1221_1,_w_6133,n268_0,_w_8944,_w_9021,n283_0,_w_15733,n760_1,n265_0,_w_5616,_w_6547,_w_16287,_w_10271,n499_0,N341_13,n394_1,_w_15625,n1621_0,n226_0,N324_6,_w_6659,_w_13865,n489_0,_w_5435,n244_1,_w_5602,n1860_0,n1239,n452_0,n285_1,_w_15615,_w_15387,n1782_1,n294_1,_w_7866,n1094_0,_w_12240,n732_1,_w_9379,_w_5940,_w_8449,_w_8909,n1746_0,n371_0,_w_8527,n750_0,_w_6846,n372_1,n1432,_w_15670,N154_18,_w_5732,_w_6523,_w_12855,_w_7664,n297_1,_w_6073,_w_16143,N494_8,_w_11968,n1706_0,_w_9464,n417_1,n109_1,_w_10608,_w_7137,n1662_0,N511_17,_w_12661,n109_0,_w_12719,n635_0,n1067_1,_w_12998,n1036,_w_7389,n1067_0,N392_3,n950_0,n48_0,n303_0,_w_6555,n423_1,n341_1,_w_12759,n1165_1,n304_1,_w_11978,N392_19,_w_14556,_w_12393,n1033_0,N392_17,_w_10089,N392_16,n525,n270_0,_w_12713,n1097_1,N392_12,N392_4,N239_10,N477_14,n1344_1,_w_14528,n646_1,n360,n899_0,_w_9665,n646_0,_w_6501,n1055_1,n751_0,_w_11912,_w_7161,n466,n478_0,n943_1,_w_15588,n593,_w_11565,n320_1,N392_15,n97_1,n1172_1,N273_13,n783_1,_w_6404,_w_6382,n1838_1,n1838_0,n643_1,_w_10622,N375_12,_w_7967,n643_0,n1581_0,n1428,n1534_1,_w_13594,N35_6,_w_7420,n1534_0,_w_15797,n186_0,n330_1,_w_15158,n1878,n132,n669_0,_w_5550,_w_6873,_w_12729,n528_1,_w_8626,n330_0,_w_15096,n703_1,_w_8384,_w_15568,_w_9968,n1703_1,n966,_w_12092,_w_5817,n1140_1,_w_10224,n1140_0,n1879_1,_w_9424,n338_1,_w_5687,N273_7,n444,n983_0,n289_1,n420_1,n809,n508_1,_w_7804,_w_10458,n1063_0,_w_9976,n181_0,n656,_w_12243,n1389_1,n1389_0,_w_8659,_w_10744,_w_10324,n840_1,n348_1,n348_0,n171_1,_w_10263,_w_14184,n1692_1,_w_8220,n1612_1,n1869_1,_w_8451,n356_1,_w_9015,_w_12159,_w_11093,n1365_1,n97,_w_14473,_w_12081,n1215_1,_w_14064,_w_5842,_w_13448,n262_1,_w_13436,_w_7291,_w_10947,n1085_1,n1098_1,n1156,n366_0,n1700_1,_w_12901,N239_7,_w_6458,n1700_0,_w_11460,n675_1,_w_7194,n986_1,_w_10826,n1347_0,_w_10267,_w_16184,_w_13170,n418_0,n1324,_w_6769,_w_14529,n702_0,_w_6809,_w_7474,n100_0,_w_15386,n603_0,n1069_1,n1356_0,n376_0,n456,n381_1,n1215_0,_w_13353,n1241_1,_w_13030,_w_7605,_w_9821,n825_0,_w_8691,n475,_w_10132,n892_0,_w_14376,n1042,n1103_1,n1167_1,_w_14986,n1167_0,N35_11,n387_0,n865_1,_w_13719,n424_0,n1650,_w_9128,_w_8617,n1805_0,n557_1,n1876_0,n1073_0,n94_0,N18_16,_w_8918,_w_7444,_w_8877,N18_14,N18_13,_w_15871,_w_7814,n835_1,n1097_0,_w_8937,_w_13962,N18_10,n1178_1,N18_9,_w_11928,n1764,n415_0,_w_7358,N18_7,N494_11,n52_0,_w_7135,n856_1,n1470_0,N18_1,N18_0,n624_0,n1124_0,_w_9831,_w_10442,N511_2,_w_10542,N358_11,n88_1,_w_15968,n399_1,n437_0,_w_13325,n405_1,n546_1,n406_1,_w_12899,n1517_1,n406_0,_w_12942,n409_1,n514_0,_w_14222,_w_7797,N375_19,_w_9775,_w_12297,n239_1,N375_18,n830_0,n1021,_w_14579,_w_10590,n1159,N375_10,n1293_1,_w_6468,N375_9,_w_8006,N375_8,N375_6,_w_15891,_w_5339,N409_4,n754_1,_w_10844,n390_1,n177_0,_w_6764,N375_0,_w_9479,n1697_0,n970_1,_w_8497,n165_0,_w_13188,n697_0,n901_1,_w_8848,n901_0,n338_0,_w_10221,n1440_0,n1607_1,n994_1,_w_5570,n617_0,_w_6267,n426_0,n334,n1894,_w_16049,_w_5996,_w_12614,n1348_1,n769_0,n1467_1,_w_12494,n433_1,_w_12134,n1257_1,n1860,_w_8141,n1257_0,_w_11271,_w_7826,N86_16,n1181_1,n1028_1,n1750,_w_8790,n1181_0,n1251_1,_w_12856,n283,_w_16117,n1183_1,n146_2,n146_0,_w_12781,n217_0,_w_11138,_w_7213,_w_12268,n642_0,_w_11868,_w_6911,n440_1,_w_14746,_w_9953,n442_1,n442_0,_w_11395,n1018_0,n920_1,n472_1,n1518_0,n1808_0,_w_9432,n453_1,_w_10157,n453_0,_w_13714,n810_1,n57_0,n922_1,_w_11112,n1000_1,n922_0,_w_12062,n793_1,_w_10078,_w_6666,n1809_0,_w_6807,_w_11234,_w_7155,_w_12380,_w_7107,n961_0,_w_8814,n460_1,n548_0,n914_1,n914_0,N392_0,n1473_1,_w_6292,_w_12954,n887_0,_w_6239,n774_0,_w_7095,n1289_1,n466_1,n345,n335_1,n468_0,n1339,_w_13680,n189_1,_w_11771,n189_0,_w_12154,_w_6473,_w_10925,n196_0,n805_0,_w_14695,_w_5749,_w_10164,n1719_0,_w_5804,_w_11329,_w_9762,_w_9896,n1019_0,_w_8307,n492_0,n1684_1,n1859,_w_8758,_w_9288,_w_14523,n798_1,n897,_w_12534,n498_0,_w_5471,_w_5787,n1206_0,_w_10243,_w_10821,n1360_1,_w_7078,n455_1,n741_1,n1879,n507_1,_w_14270,n507_0,n1555_0,_w_10628,n292_1,_w_14753,_w_12226,n621_0,_w_11103,n805,n503,n1098_0,n881_0,n309_0,n214,_w_11672,n277_1,_w_7492,N290_19,n831,n1100_0,n910_0,n1371_1,_w_11575,n305_1,_w_14011,_w_13026,_w_12151,n1101_0,n150,_w_15159,n1104_1,n666,_w_5584,n1104_0,n625_0,n1796_0,_w_11231,n1311_1,n1303_0,n1106_1,n299_1,_w_15985,_w_14157,n96,N1_0,n1743_1,_w_6787,N443_14,n570,n42_0,n1119_1,n1122_0,n752,_w_14538,_w_6973,n1125_1,n583,n1127_1,_w_12270,n1132,_w_10883,n532_0,n1276,n111_1,n1841_0,n1127_0,_w_13692,_w_8132,_w_9126,n1856_1,_w_10822,N35_10,n872,N307_11,_w_6528,n1679_1,n1758_0,_w_11779,n862_0,_w_12164,_w_11625,n871_0,n1139_0,_w_8756,_w_9600,_w_6052,n757_1,n1142_0,_w_7635,_w_9664,_w_10119,n1612_0,_w_15831,n1658,_w_6259,_w_13489,_w_12113,n1148_0,_w_7975,_w_15257,n1155_1,_w_5346,n1734_0,_w_6339,_w_7753,_w_12445,_w_11509,n534_1,_w_8329,n1329,n1561_0,n1161_0,n475_0,N273_6,n261_1,n1163_1,n1065_0,n608_1,_w_15869,_w_8717,n1164_1,_w_10721,n821_0,_w_14724,_w_9783,_w_16040,_w_5356,n868_1,n1164_0,N137_6,_w_12091,n161_1,N426_16,n465_1,n1170_1,n1173_0,n1735_0,n1898_1,_w_11790,_w_5639,_w_6422,_w_14780,n1898_0,n1180_1,n1182_1,_w_12657,_w_8244,n240_1,_w_11848,n768_0,N273_17,_w_14733,n1818_1,_w_10101,_w_15867,_w_11180,n588,_w_15232,_w_6363,n1818_0,n1359,_w_6343,_w_9062,n1184_1,n351_0,n1215,n1187_1,_w_12470,_w_10418,_w_8322,n1115_0,_w_9044,_w_7520,_w_13023,n414_0,n746,_w_8673,n1190_0,n960_0,N86_6,n1193_0,n995_1,n1566,_w_10864,N375_17,n1421_0,_w_10655,_w_10002,n1203_1,N443_13,n1203_0,n1342_1,_w_6598,N137_0,n1342_0,n1205_1,_w_6344,n728_0,n1526,n501_0,n706_1,n250_0,_w_8806,_w_11677,N426_2,n1217_1,n1218_1,n1218_0,n1783_0,_w_7186,n1503_0,n430_0,n1578_1,_w_12686,_w_10589,n1653_1,n1578_0,_w_13270,n1581_1,n1822_1,n1815_1,n326,n1230_0,_w_7010,_w_11306,n1599_1,n754_0,n720_1,n295_0,_w_8760,n1232_1,n1797_0,n1232_0,n1235_1,n1236_0,_w_14819,_w_10524,_w_5667,_w_12008,n1238_1,n997,n1564_1,_w_13235,_w_7890,_w_14693,_w_11208,n1833,_w_9887,n1845_0,n1846,_w_7167,n1245_1,n911_1,n1245_0,N205_9,n1256_1,n1256_0,n527_0,n1625_1,n723,_w_11650,n258_1,_w_13708,_w_9650,n1262_0,n1263_0,n1126,_w_6065,_w_14280,n1270_1,n1270_0,_w_13127,n1278_0,_w_9860,n893_0,_w_11408,N375_16,_w_8855,n1266_0,n1765_0,n1267_1,_w_11867,n1268_1,_w_12139,_w_8912,_w_15679,n1271_1,_w_15841,_w_15510,_w_8004,n1273_1,_w_13981,n1274_1,_w_5657,_w_14344,_w_11553,n132_0,_w_9377,_w_13113,N35_4,n1275_1,n1279_1,n1268_0,n1280_1,n1003_0,_w_8134,_w_8305,_w_13668,_w_9656,n594_0,n1280_0,n1282_0,_w_13068,n1851_1,_w_12086,_w_10138,n1283_1,n385_1,n901,_w_15942,n1780_0,n1283_0,n890_0,n1284_1,N103_1,_w_7828,n1285_0,n685_0,n1572,_w_8671,n1866_1,_w_8482,n705_0,n1297_1,n1297_0,n1299_1,n1299_0,_w_8312,_w_6376,n1300_0,_w_10818,n1500_1,_w_16246,_w_11239,n1300_1,n1305_0,n1309_1,_w_9146,n1326_0,n388,n1104,_w_5961,n1309_0,_w_6912,_w_7479,n1483,n1312_0,n426_1,n1314_1,n1314_0,_w_6790,_w_9769,_w_6881,n1315_1,n312_1,n1401_1,N222_3,n1158_1,_w_14245,n1369_1,_w_13039,n1317_0,_w_12728,n1442_1,_w_10569,_w_6977,_w_14474,n1318_1,n869_1,n1430_0,n1318_0,n1201,n639_1,_w_8559,_w_10949,N86_12,n1320_1,n836_0,n1321_1,_w_13168,_w_12647,_w_9088,_w_10639,n1321_0,n1134_1,n1327_0,_w_16243,_w_13760,n1330_1,N69_0,n1333_1,n1143,n977_0,_w_6302,n1335_1,_w_5827,n168_0,n1082_0,_w_10234,n715_0,_w_7454,_w_8842,n1364_1,_w_6476,n1339_0,_w_8092,n1674_1,_w_9505,_w_10298,n1341_1,n1351_1,_w_9645,_w_9832,n1354_1,n840_0,n1673_1,_w_8805,n1673_0,n481_1,_w_7682,n78_2,_w_9451,n1359_0,n804,n1739_1,_w_5792,n79_0,_w_14653,_w_9853,_w_10889,n1145,n1370_1,_w_13280,n483_1,n1248_1,n1374_1,N358_14,n258,n1374_0,n642_1,n1062_0,n1375_0,n1584,_w_12183,_w_8193,n1254_1,_w_15399,n1793_0,n150_0,_w_9061,N290_4,n1379_0,_w_14754,N154_8,n1380_0,n878_0,n469_1,n293,n1382_1,_w_15672,_w_8173,N511_5,n1382_0,n1383_1,_w_8770,n767,_w_10788,n1453,_w_10600,n1208_1,_w_15044,_w_11697,n1385_1,n1386_1,_w_6795,_w_14167,_w_8881,_w_9791,_w_7121,n102_1,_w_13491,_w_9300,n107_1,n1392_1,_w_11506,n857_0,n1392_0,_w_11126,N86_5,_w_6068,n60,_w_12742,_w_12605,n543,_w_14861,n1394_1,n1338_1,_w_5502,n1394_0,n1395_0,_w_7649,n273_1,n1397_1,n91_0,n1093,_w_14109,_w_13895,n828_0,_w_9504,n1090,_w_6175,N239_9,n417_0,_w_7697,_w_6197,n1899,_w_6241,_w_9318,_w_11861,N171_2,n675_0,n1088,_w_15517,n1187_0,n848,_w_6709,n1124_1,n1064,n1773,_w_9358,N171_14,_w_9700,n120,n1529,n237_0,_w_11448,n510_0,_w_14234,n1460_1,_w_7375,n1558,N52_6,_w_15736,_w_6471,_w_13412,_w_7243,_w_14348,n194,n823_1,n1232,n1762,_w_16176,_w_10142,n1220,n73,_w_12740,_w_8288,_w_11831,n1058,n1051_0,_w_11673,n645_0,_w_5490,_w_5673,_w_8323,n1052,_w_14001,n1404,_w_5469,_w_12985,n949,_w_5945,_w_11084,_w_7495,n1041,_w_7849,_w_13476,_w_10852,n1550,_w_16042,N205_7,n1774_1,n1736_1,N103_8,n1115_1,n1388,n299,_w_10745,n315_1,_w_14086,_w_9800,n1733_0,n1768_0,_w_11776,_w_5672,n906,n1008,n1006,_w_11439,n1002,_w_6783,n1178_0,n1001,n739,_w_7103,N307_7,n938_1,_w_15806,n192_1,n1188,n806,_w_7913,_w_11793,n575_0,_w_13036,n1775,_w_13226,n86,_w_9255,n980,n976,n975,_w_9895,_w_14385,n971,_w_9223,_w_13125,n968,N426_12,_w_8564,_w_7185,n965,n516_0,N103_18,_w_7603,_w_8796,_w_10877,n896_1,_w_11800,_w_6710,n1465_0,_w_15703,n1377_1,n1527,N477_7,_w_5449,_w_15870,n1608_1,n352,n1197,n78,n959,n953,_w_8355,_w_12016,N341_19,n1152_0,_w_6195,n946,_w_13651,n1347_1,n941,n954,_w_9083,_w_8417,n938,_w_6687,_w_5321,_w_8701,n522,n1658_0,N273_9,n813_1,_w_11751,n1756_1,N426_10,n236_1,N290_1,n1231,_w_13683,n172,_w_10232,N324_0,n935,N86_9,N103_12,n578,_w_9236,n926,_w_9331,n1084,n1030,n1288_0,_w_5643,_w_10807,n1194,_w_8056,n732,n920,N1_18,_w_14997,n1185_1,n312_0,_w_9313,N477_8,n1403_0,n506,_w_13805,_w_6915,_w_8349,_w_13276,n104_1,n916,n1481_1,n1143_0,_w_6600,_w_14774,_w_7536,_w_14154,_w_7917,_w_8926,n1822_0,_w_5520,n905,n1068,_w_12465,_w_5376,n1755_1,n297_0,n895,_w_15851,_w_6936,n1225,N324_16,n402_0,_w_9038,_w_9369,N290_13,n1452_1,_w_15884,n772,n890,n1046,_w_10188,n885,n1781,_w_13934,n1494_1,n590_1,_w_6041,_w_8201,n1779,N205_5,_w_11396,_w_8828,_w_12017,n884,_w_10367,_w_7122,_w_9718,n880,N409_11,_w_16180,_w_9415,n828_1,_w_13632,_w_8108,_w_9185,_w_11894,N86_18,n1587,_w_15508,_w_8695,n1247_1,n1835_1,N205_3,n1272_1,_w_8394,_w_7978,n1471_1,n133_1,n765,n1512,n677,_w_8583,n1852_0,_w_6385,n853,n201_1,_w_7331,_w_12761,N103_11,n446_0,n846,n696,_w_15249,n136,n1511,n842,_w_8123,_w_14541,_w_8555,n1214_1,_w_10045,_w_11535,n836,n830,n490_0,n1865,_w_6801,n829,n828,_w_12432,n367_0,N528_4,_w_6557,_w_8892,n1646_0,n1438,_w_11314,N171_9,_w_6921,_w_12220,n827,_w_15671,N120_12,n1593_0,_w_7312,n121,n750_1,_w_16010,_w_6526,_w_14975,_w_11447,n824,n823,n422,n821,n1040,n1610,_w_11653,N375_1,n888,_w_11312,n612_0,n1269_1,_w_5665,_w_10056,n1784_0,n807,_w_15743,_w_6149,n1381_0,n1603_0,_w_12291,n855,n802,n1131_1,_w_7862,n332_0,_w_15233,n1116,n41_1,n795,n912,_w_9266,n293_1,_w_16160,_w_9176,n788,n136_0,n1863,_w_14205,n1287,_w_10840,_w_10266,n294_0,_w_8093,n542_0,N69_14,n1145_1,n211_0,n399,_w_11919,n758,n1017,n1783,n790,_w_13262,_w_6850,n147_1,n1081,_w_11859,N443_17,_w_11250,n1071,n548,_w_7763,_w_16262,_w_9663,n602_1,n302_1,_w_13549,n776,_w_14314,n775,n1449_0,_w_15878,_w_12547,n812,n1515_1,_w_6524,_w_16228,n1884,_w_13373,n1305_1,n762,_w_9748,_w_11908,n367,n379_1,n760,_w_15103,n969,_w_7051,_w_13379,n152_0,_w_8962,n1023,_w_10024,n173,n1615_0,_w_12459,_w_11947,n1010,n449_1,_w_6188,n149,n1373_0,_w_15432,_w_12440,_w_7884,n1025,n763,_w_6549,n824_0,n1856_0,_w_5327,n742,n210_1,_w_14437,n737,_w_14527,n1467_0,n731,N511_18,_w_5909,_w_13146,n1065,_w_7466,_w_14267,_w_7597,n112,n1641_1,n1712,n1356,_w_13588,n1312,_w_10433,n1089_1,N443_10,n632_0,_w_9553,n748,n1112,_w_11055,n466_0,_w_6916,n781,n817,n384_0,n684,N35_14,_w_6377,N103_16,_w_7301,n1196,n929,N392_11,n59_0,_w_5501,n1319,n1570,_w_7245,_w_10262,n718,n717,n1683,_w_14815,_w_14015,n222_1,n713,_w_9317,n119,_w_8114,n1732_1,n1808,_w_7116,_w_7879,n845,_w_8532,n738,_w_9490,_w_12771,n234_0,n484_0,n707,n706,n878_1,n467,n1793,_w_10446,_w_6048,_w_12993,_w_11548,_w_6335,_w_7744,n694,n995,n736,n1603,_w_11907,_w_5595,_w_12024,n446_1,n298_1,N460_2,n1083,n1641,_w_8435,n1175_1,n634,n692,_w_5949,n114_0,N120_1,n1799_0,n690,n936,_w_16095,_w_9520,N545_1,_w_12556,_w_9856,n1166,n683,n579,n688,n687,n459,_w_11135,n913,_w_12784,n682,n1209,n1526_0,_w_15564,n1551_0,_w_6462,_w_9211,n731_1,n399_0,_w_16018,_w_11628,n713_0,_w_10726,_w_6141,n675,_w_10658,n674,_w_16113,_w_15674,n1869,n1596_1,n102_0,n673,_w_14734,n144,_w_15618,n670,n1535_0,n1413_0,n1452_0,n81_1,n662,_w_8179,n1476_1,_w_9217,_w_5308,n655,n370_1,n463_0,n1536_0,_w_8509,N341_3,N392_2,_w_14661,n1724_1,_w_11243,n946_1,N137_1,_w_6193,n1308_1,_w_7467,n127,n943_0,n1387,_w_11512,_w_5447,_w_15695,n959_1,_w_14929,n253_0,n327,n1591_1,_w_12373,_w_11645,n800,_w_6400,n627,_w_11586,n907,_w_10080,n1737_1,N239_4,_w_9430,_w_7736,n365_1,_w_10730,n781_1,N273_16,n661,_w_16132,n846_0,n622,n747_1,_w_12200,n1191,n77_1,_w_6143,N443_7,_w_11264,_w_9881,_w_14721,n1543,_w_5897,_w_15689,n344_0,N86_10,n125,_w_11371,_w_9492,n1481_0,n1118_0,n780,N256_3,_w_13414,n618,_w_15584,_w_6011,n617,_w_7309,n542_1,n300,n1207,_w_10803,n1294,n616,_w_11717,n513_0,n1290_0,n1060,n615,_w_7868,n339,N69_8,n862,n1484,n608,_w_13466,n700,n607,n1709,n437_1,_w_7720,_w_11967,_w_7836,n67,_w_10027,_w_14833,_w_14070,n1542_0,_w_8057,_w_7843,_w_10987,_w_9261,_w_10417,n223_1,_w_6182,n1722_0,n368_0,_w_13422,n948_0,n597,_w_13190,_w_11071,_w_7168,_w_9472,_w_14679,n1251_0,n1045_0,n1475_0,n1778_1,n587,_w_15074,_w_10875,n542,n923,_w_9691,n586,N324_18,n1205_0,n1118_1,n333_0,n1732,_w_6479,_w_14799,_w_9933,_w_7148,n585,_w_6090,n1420,_w_9954,_w_13498,_w_8030,n624_1,_w_15885,n1789,n991_1,_w_5655,n1379,N137_16,n1242_0,n1281,n1657,_w_13510,n663_1,n1664_1,_w_14039,n455_0,n899,n541_1,_w_8076,_w_11446,n271_0,n1020,n626,_w_5751,n1246,_w_7081,n198_1,N35_19,n735,n1013,_w_12651,n712,n108,_w_14555,n191_1,n1178,_w_8281,n759,n1133_0,_w_11729,n448_0,n984,_w_12263,n1378,_w_8404,n541_0,n491,n96_1,_w_15291,_w_15220,n575,n1151,n567_1,_w_15794,_w_11402,_w_8519,n1289_0,_w_12864,_w_5631,n660,n944,_w_9419,n256,n834_0,n835,_w_16164,_w_5623,n1548_0,n565,n1031_0,n864,_w_8058,n1094,_w_12047,n554,n459_0,n234_1,_w_7409,n223,_w_13453,n107,n612,n1622_1,_w_10207,n549,_w_10990,n631,n547,n1718_1,_w_13106,n1843,_w_13309,_w_9943,n204,_w_15792,_w_6284,n629,_w_8733,n1643_1,_w_15856,_w_6280,N290_11,_w_15975,n1662,_w_10306,_w_5754,n1638_0,n540,n1640_1,_w_9194,_w_8010,_w_14718,_w_8829,_w_15781,n1107,_w_13560,_w_6096,n1311_0,n1502_1,n159_1,n1866,_w_6045,n1777,_w_15363,n1770_0,n478_1,n870,n915,n1841,n533,_w_12429,n182_1,_w_14935,n208,_w_6148,n410,n1820_0,_w_12000,n1212_0,n1335_0,_w_11922,n530,n528,n337,_w_10828,N290_0,_w_14229,_w_7580,n357_0,n777_0,_w_14435,_w_13465,_w_8228,n1332,n1075,n53_0,n553,_w_12765,n635,_w_10336,_w_8922,_w_14918,n219,_w_9069,_w_6308,n535,_w_12961,n744_0,_w_15769,n1591_0,_w_12583,n1374,_w_5359,n1697_1,_w_14883,n213,n999,n88,_w_12209,n1751,_w_11303,_w_9000,_w_9584,n1004,n1214,_w_13864,n741,n778,n679_1,_w_15918,_w_6428,n735_0,n209,n507,n66,n1186_0,n880_1,n939_0,_w_15247,_w_5791,_w_6487,n424_1,_w_5663,_w_7252,n490,n955,_w_16130,_w_11636,_w_11367,n709,n778_1,_w_8631,n201,_w_11762,n1323_1,_w_14302,n1853_0,n1680_0,_w_5383,n373,n801_1,n1615,n284,n1079_0,n1049,n571,_w_14146,n354_1,n1106,n129,_w_13096,n354_0,n115,_w_7278,_w_5632,_w_9730,n1315_0,n614_0,n36,_w_11753,_w_11661,_w_9874,N460_1,n1135,n1028,_w_13892,n616_0,_w_5347,n875,n229,n183,_w_11049,n1606,n1506_0,_w_7373,n1697,_w_10899,n844,n1806,_w_6283,_w_13388,n799_1,n972,_w_8879,n171,n354,_w_13834,_w_11787,_w_6814,_w_8832,_w_15725,N341_0,_w_13531,_w_5484,_w_15514,n789,_w_12805,n1460,_w_10647,_w_5990,_w_14822,n62,n160,n1113,n678,n136_1,n871,_w_9482,N154_10,n714_1,n668,N171_1,_w_6080,_w_13867,n723_1,_w_6154,n1401_0,_w_15726,_w_8326,n477,n62_0,n1602_0,n138,_w_6106,N222_0,n324_0,_w_15017,N375_13,n489,_w_11685,_w_10632,_w_7811,n638,_w_15192,_w_12025,n1243,_w_14271,n917_0,n458,n443,_w_15684,n1091,_w_10768,n159,n1747,_w_6728,N511_1,n415,n1499_0,n193,n1175,_w_15655,n1691,N426_13,n1259,n663,n1886_1,n42_2,_w_10340,n1762_0,_w_11505,n306_1,_w_7551,_w_13211,n772_0,_w_5902,_w_11899,_w_6171,n1039,_w_10254,n1024,_w_6958,n1598,_w_14600,_w_11481,n1085,_w_8959,_w_10456,n1544_1,n296_1,n76_0,_w_6416,n148,_w_13483,_w_12669,_w_11688,n1713_0,N171_13,n350,n652,_w_7734,N477_19,n896_0,n249_1,n419,n1466_0,_w_12841,n1300,n1611,n572,n207,n1695_0,_w_5927,n1459,n1628,N409_12,n104,n510,n580,n907_1,_w_7796,n1707_1,n1371_0,_w_11585,_w_8022,_w_12793,_w_11835,n1479,n1690,n1682_0,_w_8154,_w_11977,n484,N239_19,n43,_w_6582,n838_1,n941_1,n766,n681,n198,_w_11179,n1253_1,n454,n1808_1,n1548_1,N103_6,n1226,n1752_1,_w_6066,n693,n430,n185_1,n1832_0,_w_9801,n737_0,_w_8356,_w_10451,n216,n1730,n1419_1,n639_0,n1778_0,N511_3,n1880,n740,_w_9940,n676_0,_w_16079,n401,N477_1,n1579,_w_9149,n1782,n1173_1,n685,n641,_w_13285,_w_5625,n1182_0,n195_0,_w_6545,n245_1,n1756,n1077,n903,_w_12851,n1056,_w_8934,n374_1,_w_14820,n1715_1,_w_5378,_w_7231,n162_1,n1176,_w_7441,n1169,n1070,N409_19,_w_8878,N273_1,n170_0,n1186,n385_0,_w_8128,n851,n1087,_w_8658,n1275_0,_w_8749,_w_14198,n122,_w_8103,n757,_w_8961,_w_6122,n197,_w_9679,n1513,N222_11,n1665_0,n94,_w_12846,n1052_1,_w_15099,n111,n377,_w_11455,n1584_0,n42,n436,n1541,n651,n1506_1,n1233_0,N375_7,n374,_w_5682,_w_12446,_w_10623,n221,n59,_w_9545,_w_14286,_w_13968,n206,N477_2,_w_12415,n1137,_w_9580,n1177,n801,n859,_w_12433,_w_12313,N511_6,_w_7416,_w_14542,n815,_w_7933,n101,_w_8292,n1223,_w_9314,N171_19,n459_1,_w_8613,_w_11286,n944_0,_w_5696,_w_12525,n202,_w_7361,_w_8535,_w_8702,n1678_1,_w_12467,n1116_0,_w_6346,N494_13,_w_10926,n932_1,n710,n1634_1,_w_14141,_w_9969,_w_8232,n141,n585_0,n1541_0,_w_5915,n293_0,_w_5385,n1615_1,_w_6232,_w_7554,N18_18,_w_15532,n1809_1,_w_14288,_w_13949,n222,n1825_1,n1061_1,_w_7455,n200,_w_13675,n1647_0,n1071_0,_w_12266,_w_11430,_w_7792,n164,_w_6115,N18_6,n469_0,n1367,n1462_0,n654_1,_w_7274,n289,_w_9086,_w_16126,n102,n1130_1,_w_6671,_w_11889,_w_10635,n794,n471,n501_1,n329,N205_2,_w_11957,_w_6082,_w_5809,n951,n545,N256_14,n309,n225,_w_12963,n1836_0,n1422_0,_w_15589,n499_1,n1515_0,n312,_w_12941,n474_1,_w_8073,_w_13816,N188_1,n185,n1147,_w_7286,n1384,n402_1,n680,_w_13978,n679,n1519,N154_12,N154_11,n1685_0,_w_15252,_w_13688,n1508_1,n1355,n1230,_w_9500,n1083_1,_w_8168,n1209_0,n237,n691_1,_w_10476,_w_6100,n750,n1428_1,_w_14087,_w_5409,_w_8561,n1678,n1656,n421,n498,_w_7595,_w_7477,n1366_1,_w_7247,n1883,n852_1,N290_3,n232_1,n563_0,_w_14745,N69_9,_w_10061,n277,n575_1,n54,_w_14383,N324_13,_w_14808,n147_0,n1095_0,_w_14356,n550,n113,_w_5588,_w_8575,_w_15727,n1676_0,_w_5604,n138_1,N392_10,_w_16237,_w_10382,n48,_w_12323,n686,_w_11600,_w_5881,_w_6306,_w_6918,_w_13254,n392,_w_13812,_w_13776,_w_9096,_w_5414,_w_12237,_w_11631,_w_6943,_w_7058,_w_10567,n462,_w_9983,n787_1,N324_12,_w_16138,n1097,n1316,n1381,n1345_0,_w_10696,_w_9564,_w_14513,n332,n325,_w_16044,_w_15292,N120_8,_w_9813,n445,n1286_0,_w_7937,n145,_w_11809,N341_8,_w_15315,n1317_1,_w_13765,n1472,n581,_w_13347,_w_7037,_w_9880,n733,n978,_w_7218,_w_7545,n427_0,n1224_0,_w_13224,_w_10183,n1273,n1734,_w_5493,_w_5585,_w_6433,_w_11982,_w_8214,n866,n341_0,n1125_0,n1628_0,n501,_w_6018,_w_7275,n286,n839_0,n517_0,_w_7265,n1009,_w_10177,_w_7724,N290_15,_w_8917,_w_5540,_w_10397,n361,n493,n1765_1,n147,n1287_1,N256_19,n1555_1,n1815,n1653,n438,n1222,n318_0,n1072_1,_w_9900,_w_15469,_w_14337,n1398_1,n79_1,N205_19,_w_5946,_w_5621,_w_15388,n1629_0,_w_10634,n396,n1795,n356_0,_w_7152,N273_8,_w_12324,n1569_1,_w_5617,_w_15970,_w_8710,_w_8720,n1163_0,_w_6597,_w_14854,_w_14494,_w_10173,n1069,n188_1,n720,n316,_w_5789,n485,n1070_1,n1547_0,_w_8990,_w_13609,n364_1,_w_9605,N18_17,n290,_w_9587,N528_2,_w_9932,n1082,_w_12454,_w_11240,n599_1,n423_0,n827_0,n1715,n573_0,n863_0,n1827,n1069_0,n881_1,_w_11669,n1820_1,_w_6119,n1625,n623,_w_10459,n69,N256_2,n365_0,n259,_w_11083,_w_8847,n196,_w_9858,_w_8378,n77,n57,n531_0,_w_12046,_w_11546,N307_12,_w_8567,n522_1,n140,n176,N477_15,n1599_0,n1391_0,_w_9960,n161,n181,_w_13057,n85,_w_12601,_w_12045,_w_7117,n561,_w_12128,n1433,_w_12924,n1151_0,_w_9627,n549_0,n87,n174_1,_w_10974,n189,n960,n955_1,_w_6935,_w_14740,n236,_w_5706,n858,n1253_0,n104_0,n1320_0,_w_7460,_w_9815,N120_13,_w_13474,_w_10750,n599,n953_1,_w_5460,n212,_w_9537,_w_6505,n1459_0,n1675,_w_6329,N86_14,_w_7124,_w_12500,n886,n1095,N18_5,n1249,n1687,n317_1,_w_5988,_w_9596,n1755_0,n1377,n368,n1489,_w_13707,_w_5968,n1613_1,n1793_1,n1494,_w_13063,n1614_0,_w_6946,_w_7598,n1654,_w_9307,n1281_1,n700_0,n931,_w_8379,_w_9644,_w_11433,_w_6630,N307_16,n315,_w_15748,_w_9712,n417,_w_7284,N477_12,n1879_0,_w_13880,N375_2,n799,_w_16265,_w_8880,_w_9552,n36_1,n539,n335,n738_0,n95,n398,n958,_w_7190,N392_9,n619_1,n1085_0,_w_12867,n1761,n1854,_w_13660,n170_1,_w_9441,_w_9536,n833,_w_14413,_w_13103,n275,n1409,n642,_w_10465,_w_6099,_w_16186,_w_14057,n974_1,n394,_w_14758,_w_6723,n431,_w_12679,n1686,_w_8678,n1479_1,n1229,_w_12955,_w_10900,n1338,_w_12182,_w_7614,n814,_w_10810,n81,_w_14596,n1021_0,n520_1,n1372,n347,_w_6123,_w_13051,n427,N52_1,n1027_0,n110,n1272,n230,n170,_w_13811,n178,n487,n917_1,_w_13858,_w_5504,_w_7204,n1791_0,_w_9661,_w_9911,n1587_1,n214_1,n1552_0,N137_10,_w_9688,n1464_0,_w_7452,_w_13537,n1562,_w_5819,N528_3,_w_7928,n954_1,_w_9198,n1091_1,_w_12318,n165_1,n1330,_w_10308,_w_5527,_w_9350,n1189,n382,n171_0,n729,n604,n764,_w_6969,n1724_0,n68,_w_14954,n1247,_w_6884,n1800,n270,_w_5354,N460_6,_w_10680,N52_7,_w_13518,n41,n1035,_w_15476,n1554_0,_w_7996,n372_0,n1695,N171_4,N460_4,_w_13593,n1505,n45,n353_0,n1193_1,_w_7328,n556,n561_0,n308,n624,_w_12027,n1475_1,_w_6808,n74,n1497,_w_11015,n83,n1577,_w_10122,n1436_1,n483,_w_5860,n114_1,n596,n1372_1,n1074,n513_1,n948,_w_13344,_w_5613,n866_1,N307_13,_w_7676,n233_0,n449,n734,n1872_0,_w_5890,n868_0,n1509,n65,n84_0,n521,_w_13642,_w_12755,n1413_1,n904,n1339_1,n208_1,n205,_w_8728,n598,_w_11128,n774_1,n1174,_w_11174,n933,_w_13508,N494_19,_w_6266,n1716_1,n1752_0,n1185,n1547_1,n1540_1,n977,_w_15875,n1786_1,n1061,_w_8551,n560_1,n58,n75,_w_11802,_w_8635,n837_0,n637,_w_8439,n1758,_w_9971,n1680_1,_w_11294,N188_10,n551_1,_w_12277,n1327,n187,_w_13454,n43_1,n879,n443_1,n63_0,_w_7992,_w_8741,n1738_1,N477_3,N222_13,_w_14347,n1086,n1884_0,n786,n1485,_w_14628,n1466_1,_w_10052,n525_0,_w_13763,n1556,_w_7083,n745,n63_1,n1391,_w_6716,n288_0,n609_0,_w_16100,n280,n322,_w_13870,_w_8469,n699,_w_10384,_w_7523,n240,_w_11106,n176_1,_w_14615,n1003,N426_18,_w_5429,n1735_1,_w_11578,n1802,_w_13462,n1439,_w_6137,_w_10077,n235,_w_6074,n1820,_w_15229,_w_6686,n505,_w_7670,n155_0,n1424,_w_14402,n380,n843,n681_1,n477_1,_w_7794,_w_9825,n342,_w_9811,n243,n339_1,_w_8392,N443_2,n505_0,n321_0,_w_7438,n1491,_w_15503,_w_7710,n1062,n667_0,_w_7901,_w_8747,n378,n714,_w_15097,n1597_0,_w_13814,n759_1,n1274_0,n697,n889_1,n246,_w_7923,n1632_0,n249,n321,n1128_1,_w_10325,n948_1,n798,_w_10091,n418,n863,_w_6895,_w_13879,_w_8042,_w_9115,_w_12337,_w_6237,_w_13333,n250,_w_15487,N392_14,_w_11317,n826,_w_8587,_w_7002,n251,n1761_0,_w_9949,_w_7673,n1138,_w_15888,n1396,n1171_1,_w_9632,n1896_0,n539_0,n403,_w_12392,N222_15,_w_6167,n1155_0,n1296,n889_0,_w_10274,_w_8738,_w_13236,n1357,n558_0,n930,_w_9669,_w_6889,_w_13504,n994,_w_14943,n353_1,_w_8136,n563,n755,n967,_w_6347,_w_7786,n1115,_w_14334,n1238,n1761_1,n848_1,n313,_w_7547,n810,n1149,n274,_w_6970,n283_1,_w_10206,n1236_1,_w_13550,_w_12023,n1154,n609,_w_15227,_w_7558,_w_9642,n279,_w_12376,n976_0,n302,n331,N137_7,_w_12273,n1184,N511_13,n1051,n869,_w_15303,n508,_w_12970,n1551_1,n428,_w_11409,n412_1,n1291_0,n106_0,n307_0,n748_0,_w_11874,n182,n529_1,_w_7533,_w_8183,n1829_1,_w_7369,n432,n555,_w_8895,n1600_1,N273_11,n448,_w_13393,n269,_w_8278,_w_13067,n1039_1,n655_1,n1229_1,_w_12501,n167,n499,n277_0,n226,N460_15,n1575_1,n1874,N273_12,N494_7,_w_5393,n1699,n1518_1,_w_5821,_w_12717,n1901,_w_13821,_w_13186,_w_9336,n839_1,n709_0,_w_9014,_w_9670,_w_6840,n285,n1445_1,N120_0,n287,_w_7860,n1863_1,n1406_0,_w_13134,n1112_0,n271,n218,N324_7,n372,_w_12335,n241_0,_w_13218,_w_8310,n233,n301_0,n297,_w_15612,n1046_0,n977_1,n1136,_w_7686,n574,_w_14185,_w_13158,n1034,n523,N69_16,n572_1,n371,_w_6297,n1488_0,n633,n414,n508_0,n1665_1,_w_5569,n1767_1,n950,_w_13802,n671,_w_6145,N171_7,_w_10641,n296,_w_13239,n1597_1,_w_5722,n423,_w_9938,n1211_1,n129_0,n462_0,_w_8229,_w_8280,n1303_1,n1744,N409_6,n1844,n524_0,n759_0,n1381_1,_w_6020,n421_0,_w_15124,_w_12339,_w_11747,n1162,n199,n1455_0,_w_14232,_w_8454,n852_0,n156_0,n1819,_w_8907,_w_9433,N137_5,_w_5323,n814_0,n1870_1,_w_7725,_w_9744,n904_0,n239,_w_13536,n49_1,n310,n591,_w_15471,n1710,_w_10366,_w_6718,n1433_1,n1725_0,n358,_w_9711,_w_8135,_w_6457,n594,_w_14878,N460_19,n1101_1,n55_1,n685_1,n457,n319,_w_6218,n1668_1,n320,n1172,n661_1,n627_1,N307_19,n629_0,n362,n159_0,n1151_1,n690_0,_w_8125,_w_13434,N188_2,_w_12752,n729_0,_w_15729,n472_0,n402,n328,n186,n957_1,_w_5413,N222_4,n1760,n330,n703,_w_12643,n1141,n1524_0,N52_14,n338,n1456_0,n1811_1,_w_10358,n606,_w_14009,n420,_w_12617,n346,n581_0,n1741_0,n840,_w_7991,n348,_w_6698,n1242,_w_12990,_w_5993,N375_3,n92,n369_1,n1692,N290_6,n1582_1,n838,N86_8,n1511_0,_w_6572,N358_13,N137_3,N1_15,_w_5491,n1060_1,_w_11658,n937,n1280,n962,_w_12744,n1554,n1768_1,n1059,n424,n1284_0,n309_1,N69_5,_w_13192,_w_6641,N120_17,n1514_0,n626_1,_w_6995,_w_9311,n917,n928,n363,_w_8954,n986_0,_w_10478,n1895,n344,n973_1,n1784,n366,_w_15964,_w_15320,n1290_1,_w_5598,n1596,n958_1,_w_8919,n492_1,_w_9372,n1347,n339_0,_w_8724,_w_8413,n1022_1,n1780,_w_7413,_w_9607,n535_1,n1385_0,_w_14211,_w_7357,n266,n943,_w_12700,_w_7943,n407,_w_8344,n515,_w_16205,n455,n146,_w_15496,n351,N18_8,n1324_0,n167_1,n1252,N52_17,n1894_1,_w_15556,n1726,n1391_1,n1576_0,n35,n1454,n376,_w_8997,n264,_w_6435,_w_14341,_w_11140,N477_10,_w_12653,_w_11299,_w_8744,_w_12936,n593_0,n411,_w_15330,n1536_1,n1259_0,n70,n177,n44,n446,N188_7,N154_14,n1167,n935_1,n381_0,n1383_0,n195,_w_7354,_w_12515,n387,n865,n1254_0,_w_8489,N35_3,n1458_1,_w_6205,n351_1,_w_14599,_w_6960,_w_13169,_w_7011,n1136_0,n557,_w_9403,n395,_w_16277,n493_1,n98,_w_9973,n1343,n818,n1496,_w_6508,n1437,n894,_w_7044,_w_14915,n1876,n719,_w_7924,n1692_0,_w_8420,n406,n429,_w_10123,n409,_w_14431,_w_14104,n793_0,n514,n745_0,n1584_1,_w_8718,_w_8964,n220_0,n1418_0,_w_6654,_w_10257,n226_1,n314_1,_w_8543,_w_8743,n252_1,_w_11979,n425,n533_1,_w_9340,_w_11531,n1434,_w_10335,n1350_0,n474,n426,n981,n982_0,_w_7594,_w_9922,_w_9151,n1825_0,_w_9687,_w_7619,n452,_w_14942,_w_8416,_w_12188,_w_9237,n1260_0,n1467,n1800_0,n1614,_w_8279,_w_8736,n790_1,n1470_1,n486_0,_w_7222,n199_0,n1684,_w_13757,n433,n562,N290_10,_w_14127,N120_4,n1571,_w_7363,n1445_0,n1078,_w_10360,_w_5737,n847,n1181,_w_6726,_w_9786,_w_12586,n1626_0,_w_6865,n1617_0,_w_14614,n1603_1,_w_6098,_w_7268,_w_8891,n791,n234,n447_1,_w_9349,n1139_1,n439,_w_11242,_w_5741,_w_14811,_w_8778,n1439_0,n1369_0,_w_10511,_w_10269,_w_10350,n440,n1018,_w_14067,n224,_w_13257,n453,n1001_0,_w_14082,N460_18,_w_8432,N443_3,n1424_1,_w_8950,_w_9184,_w_13100,n922,n793,n93_1,n1169_0,_w_6593,_w_16015,_w_11634,n584,n405,n457_1,n1809,n739_1,n460,_w_12762,n872_1,_w_5688,n1747_0,_w_15478,_w_14606,n1620_0,_w_16200,_w_5601,n101_0,n1838,_w_7432,n1416_1,_w_5746,n463,n433_0,_w_7587,_w_8186,_w_9634,n1045_1,n1414,N188_6,_w_14224,n774,n376_1,N222_8,n243_0,n465,n93,N392_5,n784_0,_w_13053,_w_9562,N426_5,_w_10253,_w_14990,_w_6560,_w_13369,_w_10084,n1770_1,_w_11488,n573,n1455_1,_w_16071,_w_15205,n833_0,n118_1,_w_7977,_w_13900,n137_1,_w_8586,n1149_1,n33,_w_12246,n1777_0,n1066,_w_8822,n689,_w_10479,_w_6437,_w_8027,_w_8619,n678_0,n1746_1,_w_14463,n1520_1,_w_8649,_w_11092,n1878_1,n724,_w_13371,n1755,n1116_1,_w_10155,n253,_w_14525,n468,n469,n1728_0,_w_9639,_w_9707,n1102,_w_5316,n473,n816,n1043_1,n1075_1,_w_5782,n276_1,N18_12,_w_15560,_w_12328,n658,n1014,n1583,_w_7592,_w_6554,n311,_w_10789,n777,_w_5774,n1792,n1368_0,N528_17,n1528,_w_7555,n1721_0,n492,_w_5951,_w_8405,n798_0,_w_7758,_w_9950,_w_9746,n647,_w_15923,_w_15912,n1853,n538,n1848_1,_w_12609,n397_1,_w_10615,n564_1,_w_10792,n270_1,n1200_1,n1462,_w_11267,_w_10738,n577,_w_11744,_w_10791,n1073,n636_2,_w_7055,_w_15484,_w_15274,_w_5556,n205_1,N409_1,N477_4,_w_15853,n1206,n1478,_w_9334,_w_7983,N1_10,_w_5905,n169,_w_14642,n1823,_w_8235,_w_8809,_w_15173,n676_1,n63,_w_13308,n386,_w_7332,_w_14379,n1360,n973,n504,_w_12819,n512,n1367_0,n345_0,_w_13070,_w_10985,n1734_1,n600_0,n1701_1,n664,_w_9503,_w_9052,n1659_1,n518,n698,_w_15565,_w_7748,_w_9910,n602,n292,_w_12299,n1790,_w_6612,n202_0,n1430,_w_8236,n1648,n1703,n1099,_w_9768,n1100,_w_8002,n511_0,n1290,n1311,n1152_1,_w_12964,N477_13,n1105,_w_14202,_w_13329,n1743_0,n91,n72_1,_w_6039,n783,_w_7496,n180_1,n1276_0,_w_8442,n911,n531,n1634,n1247_0,_w_6656,n1743,_w_13801,n1117,n1301,_w_7936,_w_8107,n1118,_w_5314,n1121,n1306,_w_9286,n678_1,_w_6633,_w_8642,n1724,_w_12384,n1521_0,n1123,n1124,_w_12138,n1125,_w_9165,n1423,n1171_0,n615_0,_w_13231,n1771_1,_w_15334,n1127,_w_12524,n1469,n688_1,n1791,_w_8192,n873,n1623_0,_w_13610,n1128,n1146_1,n1607,_w_15737,_w_9790,_w_10154,n1129,n1856,_w_6760,n1130,_w_6010,N511_10,_w_7334,_w_8456,_w_8530,n1133,n1134,n1139,n1499_1,_w_6705,n1180_0,N392_7,_w_10513,n1672,n1612,_w_15365,_w_9455,N35_1,_w_5925,_w_5995,_w_12132,n1026,_w_7141,n1144,n592,N154_3,_w_13451,n1518,_w_10017,n881,_w_15318,n1811_0,n1148,n1456_1,n1882,_w_6648,n727,n437,n1667_0,n1016,n1651,n1153,n1155,_w_13793,n1027_1,_w_7338,n756,_w_12919,_w_12374,_w_5848,n1157,n862_1,_w_8049,n1163,_w_7728,n1854_1,_w_8780,n1861,n1165,n1170,_w_6990,_w_13512,n1173,n1842_1,n121_0,n1291_1,n1898,N35_5,_w_7128,_w_14445,_w_8127,_w_7576,_w_10048,_w_15929,n91_1,n1511_1,n1847_1,_w_10610,n1819_1,_w_7098,n1032,n529_0,_w_9708,_w_11582,_w_9387,_w_5978,_w_11114,n1100_1,n721_1,n1183,n785,_w_9447,n1480,_w_15865,_w_9721,n1608,n229_0,n1187,_w_12002,n1285_1,_w_8434,n1588_0,_w_10918,n573_1,_w_15537,n1045,N69_19,n1029,_w_8562,n1195,_w_11133,n1787,_w_12978,n1208,n387_1,_w_12904,_w_11167,n630_1,_w_8068,_w_8202,_w_7930,n1203,n1342,_w_12106,n1204,n822,n1664_0,_w_7835,_w_9110,n1205,n1210,n1535_1,_w_9147,_w_12599,_w_10134,n1000,_w_5970,n1211,_w_8773,n1212,_w_7519,_w_16017,n1218,n68_0,_w_6260,n1219,_w_15362,n597_0,_w_6414,_w_10748,n37,_w_11060,n1578,n157,n353,n1581,n823_0,n1241_0,_w_5593,_w_13734,n1728_1,n1235,_w_6120,n1236,n768,n1529_0,n450_0,_w_8459,n1685_1,_w_8145,n1487_1,n1845,_w_15139,N171_12,n837_1,n1707_0,n1245,n87_1,n555_0,_w_6617,_w_10690,n1688,n1253,n1233,n1055_0,n1254,_w_9595,_w_9841,n728,_w_9335,n1226_1,_w_13358,n1258,_w_14690,n1407_1,n1655_0,_w_15987,n1884_1,_w_5629,n1338_0,n76,n1260,n1398,n1723,_w_6863,_w_6200,n697_1,_w_9751,n1261,_w_5833,n1018_1,n1262,n1270,n1794_1,n684_1,n1478_0,n405_0,_w_5891,n441,_w_8665,_w_14736,n1278,n126,n1267,n1268,_w_7379,n1658_1,_w_7085,_w_10029,N188_4,_w_9390,n1271,n326_1,_w_14482,n1495,_w_8630,n1274,_w_15355,_w_7762,n126_1,n1279,n572_0,_w_9221,n1284,n1288,n908,_w_7785,n1713_1,_w_8048,_w_12798,n1737_0,n1408,_w_5509,n90_1,_w_6165,_w_11664,n609_1,_w_10743,n552_0,_w_15052,n181_1,_w_6348,n166,_w_5451,_w_15696,_w_8549,_w_13440,n1500,_w_12192,n1304,n1305,n1572_1,n745_1,n863_1,_w_13828,n1307,N137_12,_w_5370,n1758_1,n1886,n1309,_w_14553,n552,n825,n430_1,n558_1,_w_8846,n1313,_w_8067,_w_15166,n347_1,_w_10053,n554_1,N35_8,n1317,_w_5377,n480_1,n544,n1442,n667,n1320,n1321,n256_1,n1005,_w_9829,n1325,_w_13656,_w_6354,_w_12624,_w_8685,_w_14475,n945,n1326,n1376_1,n1328,n1425,n1744_0,_w_5752,N239_5,n117_0,_w_6345,n1333,_w_15501,_w_15451,n1334,_w_6496,n1335,N290_9,n292_0,_w_5624,_w_15183,_w_11916,n1364,_w_16245,n304,n1337,_w_8715,n1234,n396_0,_w_9030,n1368,n495_1,_w_10971,_w_6793,_w_10036,n1410_0,_w_13014,n1341,n1345,_w_11542,n1893_0,_w_7652,n1351,n1640,n527,n769,_w_10691,n1352,_w_14300,n1043_0,n1353,_w_13142,_w_5739,_w_8137,_w_7417,n1354,n853_1,_w_14182,_w_5470,_w_7712,_w_15904,_w_15704,_w_7651,n1673,n942_1,n1358,n1130_0,n970_0,_w_7703,n1361,n1263,_w_15404,n247_0,_w_7295,n497,_w_6402,_w_10104,n1366,n908_0,_w_5652,_w_6978,_w_6825,_w_7013,n1797,_w_10334,_w_6578,_w_14243,n139,_w_7472,n1788,n929_1,_w_8212,_w_10428,n1369,_w_8989,n1140,n1371,N18_3,_w_11024,n495,n1375,_w_5431,n1380,_w_14731,_w_5401,_w_6495,n926_1,_w_8947,n1382,n639,n154,_w_9055,n1383,_w_15014,n1386,n1880_1,n691_0,_w_5345,_w_9125,_w_5357,n1730_1,_w_13062,n1244_0,n416,_w_14805,n1759,n1308,_w_5404,n1833_1,_w_11984,n1393,n1394,n603_1,_w_7586,n1824_1,n1725_1,_w_14189,n1397,_w_12411,n164_0,_w_16168,n1019_1,n1263_1,_w_15813,n1400,_w_10386,n1418,n211_1,_w_12451,n1650_1,n525_1,n715,n1405,_w_15101,_w_7320,n257,_w_14790,_w_8450,_w_9738,n1620_1,N1_14,_w_7323,_w_8177,n69_0,_w_15644,_w_14252,n526,n1407,n1411,n496_0,n1412,_w_13078,n813_0,n1415,n1157_1,n1422,_w_12340,n597_1,n1416,_w_11877,_w_5923,n1436,n956_0,N392_18,n1563_1,_w_15995,n1417,n1618_1,n1419,_w_15354,_w_10435,n1421,n1857,_w_6019,_w_7927,n123_1,n826_0,n156,n1427,_w_15123,n630_0,_w_6358,_w_5813,_w_7075,n1429,n919,_w_9848,n1431,n1662_1,_w_12224,_w_10630,n210_0,n1435,_w_5324,n1440,_w_10082,n1444,n1445,n587_1,_w_6028,n1033,n1661_1,_w_12630,_w_6513,_w_12929,n1004_1,n1446,_w_11732,n1202_1,n1635,n1517,n1054,n1447,_w_14855,_w_11690,_w_6480,n1452,_w_16147,n307,_w_8180,_w_8411,n1674_0,n1363_1,_w_16266,_w_10834,n1803_0,n452_1,n168_1,N494_14,n321_1,n676,_w_5683,_w_13364,_w_10798,n1455,n1200_0,n1058_0,_w_5405,n1456,n246_2,n1457,_w_14705,_w_7848,n1458,N494_1,n517,_w_14704,n1852_1,_w_13706,n706_0,_w_13082,n1464,n303_1,n1465,_w_7383,_w_16106,N511_7,n979,n295,n343,n1753_1,_w_14921,_w_5747,_w_8106,_w_15293,_w_9188,n1289,n1474,_w_10304,_w_5516,_w_10614,_w_8791,_w_7263,_w_9784,_w_13540,n1896,_w_6535,n1785_1,_w_9260,n1616,_w_6665,n1022,n513,n1713,_w_15922,n1481,n1373,n1840,n1627,n1482,_w_12236,_w_6305,n1486,_w_8663,_w_11472,n939,_w_8745,n1487,_w_10914,_w_7048,n1350,n1488,_w_12402,n1490,_w_8529,n1492,n480_0,n1877_1,_w_9097,n1803_1,n1493,n1667,N528_14,n1676_1,n450_1,n1502,_w_14294,_w_8293,_w_8993,_w_10869,n1503,_w_13554,_w_10566,n924,_w_5582,_w_9023,n1704,_w_6988,n878,n472,n1504,n940,n811_0,_w_7642,n650,n323_1,n1508,_w_7053,n1326_1,n242_1,_w_7485,_w_6431,n1514,n546_0,n559,n1515,n892,n1516,_w_13726,_w_6744,n1597,N171_16,N290_2,_w_8401,n391_0,_w_11743,_w_5766,_w_14813,_w_14361,n1520,n439_0,n1522,_w_13429,_w_9270,n409_0,n1867_0,n928_1,n1524,_w_12678,n1525,_w_6443,_w_8051,n985,n76_1,_w_9162,_w_7852,_w_8820,_w_15428,n115_1,N426_1,_w_6981,n1530,n1667_1,N120_18,_w_6448,n1469_1,_w_8121,N86_1,n1696,_w_9502,_w_14175,n1575_0,n1535,n176_0,_w_8269,n1889,_w_12160,n1038,n534,_w_12458,_w_5674,_w_12768,n1538,n1054_0,n1539,_w_7921,n1534,_w_8987,_w_6957,n1461_1,n1544,_w_6542,n108_0,n1545,_w_14002,n1572_0,_w_10539,n1546,n1366_0,n1547,_w_13670,n349,N35_2,_w_15832,_w_9616,n502,n563_1,_w_15580,_w_5394,_w_10979,n1552,_w_6360,_w_9411,n1729_1,n1476,_w_7581,n1844_0,_w_13446,n584_0,n987,n1184_0,n1631_0,_w_15611,_w_9506,_w_10408,n1269_0,n854_0,n1557,n1559,n1403_1,_w_9347,_w_13903,_w_12747,_w_8403,n1640_0,_w_14666,N511_12,_w_12274,_w_9045,n1564,n1565,n1568,n615_1,n1569,_w_15846,n1248_0,N409_10,N171_11,_w_5984,_w_9212,_w_12578,n1585,n363_0,_w_9040,_w_14444,n744,_w_7929,n1574,_w_9457,n1558_1,_w_12692,n893,n1576,n1468,_w_9654,n367_1,n400,n474_0,n1580,_w_14640,N273_4,N239_8,_w_6596,n1582,n902_0,n404,n920_0,_w_10149,n672_1,n702_1,_w_7329,N494_5,_w_13115,n1586,_w_14025,n88_0,n1668,_w_12699,_w_7894,n628,_w_9022,n1589,N222_5,N239_1,n1590,_w_7429,_w_6910,n1282_1,_w_14719,_w_8437,n1591,n1329_0,n1587_0,_w_5805,_w_5935,_w_8767,n1592,n40,n1593,n1765,_w_9002,n1595,n1063,n1618,n350_0,_w_7236,_w_8526,n1607_0,_w_12571,n438_0,_w_10536,n1599,_w_9884,_w_10596,N324_14,n1600,_w_10299,_w_9753,n55,n739_0,n1604,_w_16014,n751_1,n1461_0,n1669,_w_15932,n1870,n1646_1,n1509_0,_w_14658,_w_7585,_w_5611,n84,n193_1,_w_5549,_w_14457,_w_7567,n133,_w_9830,n1552_1,_w_13156,n1285,n1302_0,_w_11076,n377_1,n1353_0,_w_12401,n600,n1404_0,n278,_w_12666,_w_9075,_w_10707,n1617,_w_11492,n1785_0,n601,n1691_1,n259_1,n1621,n1623,_w_10180,n1624,n1626,N358_19,n1493_0,_w_10092,n1677_1,n46_0,_w_15534,N307_0,n1629,N137_14,n1294_0,N494_0,_w_5781,_w_6230,n1893,n1512_0,_w_15059,_w_9921,n940_0,_w_14851,_w_14187,n393_0,n333,_w_6179,n1582_0,n65_1,n1632,n952_0,n139_1,_w_9145,n495_0,n1643_0,_w_7253,n619,_w_7511,_w_8579,n747,_w_15411,_w_5546,_w_13114,n1636,n1637,_w_16141,_w_9761,n1103_0,_w_5708,n1799_1,n657,_w_11215,_w_10994,n1771,N256_6,n637_0,n1877_0,n1643,_w_8363,n1644,_w_15154,n1645,_w_15138,n357,_w_7633,_w_15427,N35_15,n892_1,n1647,_w_8063,n1170_0,n1476_0,_w_7702,N273_3,_w_15122,_w_10374,_w_5840,_w_15555,_w_14720,_w_13302,_w_8566,n1649,_w_14493,_w_6735,n36_0,N494_6,_w_5681,n265,n1619,n456_0,_w_12704,n311_0,n1896_1,_w_10507,n1683_1,_w_11914,_w_7255,_w_7821,n1712_1,_w_14804,_w_10385,n1262_1,_w_8238,n1600_0,n1659,_w_7005,_w_14920,n537,n1660,n1786_0,n1663,n516_1,n537_1,n1665,_w_13313,n1149_0,_w_8800,_w_10300,n1425_0,n1677,_w_14562,_w_6932,_w_12010,n1680,n1079,_w_9316,n1681,n520,_w_6651,n1682,n610,n1380_1,n1685,_w_12839,_w_6781,n918,n1384_0,_w_7322,n1046_1,n1835_0,n1121_1,n443_0,n925_1,_w_6147,n1427_1,n1736,_w_15055,n1013_1,_w_7618,_w_9894,_w_6492,n1390,_w_14240,_w_12488,n1190_1,_w_13837,N154_5,n233_1,_w_11929,n1702,n1821_1,_w_8799,n1267_0,n1706,n1542,_w_9321,n1691_0,n760_0,_w_15045,_w_12596,n364,_w_9991,n1707,_w_11568,n288,_w_13081,n1860_1,_w_7782,_w_10827,n1714,_w_15876,n191,n1611_0,_w_7510,_w_11442,n950_1,n524_1,n1616_1,N171_0,n235_0,_w_9763,_w_12089,n1720,_w_5768,n1721,_w_12741,n1725,_w_15706,n1322,_w_14375,_w_7532,_w_14922,_w_8043,_w_12592,_w_11078,n1728,n832,_w_5983,n1805,n1729,n143,n651_0,n1830_1,_w_7994,n874,n1733,_w_6362,n155,_w_14126,n1450,_w_8028,n784,n1012,n1454_1,_w_14364,N222_17,N69_17,n106_1,n158,n511_1,n1742,n1497_0,_w_12342,_w_6087,_w_8628,_w_9787,_w_14585,_w_13121,n1745,n1536,_w_10735,N120_19,n1753,N273_10,n1754,_w_14917,n1757,N324_15,_w_8866,_w_9727,n1260_1,_w_10117,N171_6,_w_6791,n303,n1763,n886_1,n1175_0,n47,_w_13323,_w_11269,n1768,n1693,n1769,_w_11033,n1770,_w_7525,N1_17,_w_9709,_w_14088,n526_1,n725_0,n856,n1774,n1340,n1543_1,n1778,n158_1,_w_12670,_w_6341,n1786,n1410,N222_6,n1794,N426_15,_w_7778,n1223_0,n1192,n1796,N324_10,_w_9233,n391_1,_w_8808,n1798,n1799,_w_6732,_w_9917,n1349,n1801,n942,_w_5483,n393,_w_5592,n52,n100,n766_1,n1803,_w_12254,n796,_w_14264,n657_0,n1398_0,_w_10784,n619_0,n360_0,n350_1,n1807,_w_11474,n1788_0,_w_6689,_w_13937,_w_8548,n1810,_w_6983,_w_16127,n1813,n1709_1,n600_1,_w_6380,N18_2,n1814,n1460_0,_w_9926,N256_1,_w_15178,_w_7912,_w_9283,N494_3,n1821,_w_8504,n311_1,n314_0,_w_15653,_w_7661,_w_13638,_w_5562,n932,_w_8024,_w_8194,n613_0,_w_11590,_w_9370,N290_17,n1601,n504_1,_w_9782,_w_16157,n1825,_w_8546,_w_14937,_w_13789,_w_12569,n276,n1858,n1826,_w_13897,N341_14,N69_13,n381,n1828,_w_10761,N443_4,_w_7447,_w_8470,_w_9535,n1830,_w_15253,n1831,n861,_w_13335,_w_7239,_w_11508,_w_6854,n1523_0,_w_15455,n412_0,_w_7289,_w_14106,n973_0,_w_14500,_w_6930,n867,_w_11182,_w_6789,_w_8453,n1834,_w_8618,_w_8155,N239_6,n1465_1,n1179_1,N205_16,n1847,_w_10043,n1446_0,n355,n1897,_w_9155,n1849,n1731,_w_7097,n1851,n1739,n1631_1,n754,n1588,_w_6566,n1855,n1223_1,_w_7066,_w_9429,_w_9703,_w_10919,n1548,n1864,_w_7557,n1867,_w_16090,_w_8615,n1872,_w_15371,n1521,_w_7337,n696_1,n1877,n457_0,n1277_1,_w_6841,n1881,_w_8421,n1537_1,n1250,_w_13725,_w_13111,_w_8319,_w_9979,n56_1,n1279_0,n993,_w_8365,_w_10161,n315_0,_w_14194,n1890,n536_1,n635_1,_w_15854,_w_12684,n1666,_w_7101,_w_13788,n1891,_w_6142,n486_1,n1009_0,_w_14962,n152_1,n1868,_w_9197,_w_11097,n1895_0,_w_9247,n454_1,n510_1,N375_14,_w_9252,_w_7225,n1101,_w_7364,n1527_0,n1895_1,_w_6894,n1890_0,N103_4,n1890_1,_w_15280,n1397_0,_w_9892,n1887_0,n1887_1,n1806_1,_w_5477,n1082_1,_w_9630,n1881_0,_w_8506,_w_14306,n1833_0,n1872_1,_w_9148,_w_14727,n488,n114,_w_15458,n228,_w_6116,n436_0,n1863_0,n1858_1,n418_1,n1353_1,n1478_1,_w_15613,n737_1,_w_6601,_w_5668,_w_9591,n1851_0,_w_6844,_w_12294,n852,_w_9633,n1848_0,_w_8360,n390,N494_2,n481,n1422_1,_w_5312,N1_12,_w_6253,_w_13245,_w_8521,_w_15716,_w_13473,N154_4,_w_14426,_w_5918,N188_9,n1826_1,n249_0,_w_8441,_w_10362,n280_1,n1449,_w_13234,_w_10379,n1659_0,_w_9284,n1824_0,_w_7134,n1449_1,_w_8152,n145_1,n765_1,n744_1,n1091_0,_w_6192,n623_1,_w_14547,n434,n1814_0,n795_0,n245_0,_w_7220,n1448_1,n1812_0,n1594,N137_2,n1812_1,_w_6920,_w_12693,n1797_1,N18_15,_w_5901,N154_6,_w_9527,n1796_1,N324_17,n332_1,n1213,n1794_0,n962_1,N35_0,n1791_1,_w_6838,_w_13848,n1671_1,n1787_1,n991,N358_7,_w_7646,n38,_w_7969,n306,n1842,_w_13782,_w_7214,n1781_0,_w_6688,_w_9297,n264_0,n1521_1,n1656_1,n57_1,n1764_1,_w_14737,n1762_1,_w_15169,n1749_0,_w_9920,n1112_1,n1296_0,n190,_w_12625,_w_9413,_w_10353,_w_10010,n89,_w_8498,n1746,n1741_1,n1610_1,n1385,n1733_1,n370,n1729_0,_w_11225,_w_6349,n1199,n1719_1,N154_13,_w_14840,_w_10599,n1710_0,n830_1,_w_7100,n782,n254,_w_9925,N1_7,n1549,N222_9,_w_10174,n252,n1710_1,_w_5669,n123_0,n998_1,_w_8250,_w_12577,_w_12536,n1131_0,n1544_0,n827_1,_w_11513,_w_5452,n887_1,n1183_0,n1706_1,_w_12565,_w_9353,_w_5536,n362_0,_w_5776,n1208_0,_w_10185,_w_9699,_w_15439,n1176_0,n444_0,_w_12847,n1119,_w_16202,n447,n1689_1,n1688_0,_w_16241,_w_9619,_w_7680,_w_14893,n986,n1684_0,_w_11468,n100_1,_w_6941,_w_9389,_w_10051,_w_15714,n1683_0,n771,_w_9341,n1682_1,_w_15731,_w_5969,_w_12104,n622_0,n1644_0,n199_1,_w_14021,n1351_0,n1661_0,n1094_1,n1336_1,_w_5533,n1650_0,_w_12757,_w_10481,_w_6833,_w_8122,n1649_0,n1722_1,n390_0,_w_11324,N443_5,n1649_1,_w_9099,n1889_0,n1644_1,_w_5820,n643,_w_7636,n538_1,n1299,_w_5368,_w_7262,_w_14367,_w_11603,n323_0,_w_10090,n131,n1637_0,n1154_0,_w_13644,_w_11820,_w_9442,n1412_0,n1040_0,n658_0,_w_8994,n1609_1,_w_7705,_w_7109,N239_12,_w_9577,n693_0,n625_1,n1365_0,_w_8903,n1454_0,_w_10554,n1893_1,_w_11026,n923_0,n1626_1,_w_5563,_w_14117,n551_0,_w_9673,n1499,n1375_1,n1067,_w_6738,n1784_1,_w_6927,_w_8425,n198_0,_w_14677,_w_6033,n1617_1,n743,_w_7259,N426_4,_w_6044,n1870_0,n1464_1,_w_5333,_w_9774,n1618_0,_w_12208,_w_8688,n1120,n1407_0,_w_8643,n1593_1,_w_7034,n363_1,n1611_1,n1812,_w_10656,_w_6519,_w_13983,n1590_1,n1668_0,n1639,n1573_1,_w_11407,_w_11350,n1109_0,n1484_1,n1730_0,_w_14548,_w_5559,n1585_1,n1057_0,_w_9181,n1569_0,_w_7963,_w_9409,n1567_0,N307_6,n1110,_w_6979,_w_13910,n1037,n1557_0,_w_8315,_w_15645,n733_0,n1443_1,_w_12306,n1545_0,n670_0,n439_1,_w_10355,n1113_0,_w_10039,n40_1,_w_11996,N222_12,n564,n1110_1,n623_0,_w_7132,n584_1,n1275,n1524_1,n1053,n1749,_w_7283,_w_14319,_w_14228,n273,_w_9674,n1542_1,_w_12808,n1541_1,n649,_w_15131,_w_8316,n1538_0,n1889_1,n1827_0,n1530_1,n447_0,_w_15081,_w_11050,n1790_0,_w_5622,_w_16053,_w_11146,_w_8034,_w_14259,n895_0,n489_1,_w_9333,_w_6224,n1790_1,_w_6922,n936_0,_w_7953,n523_1,_w_9575,_w_13625,_w_5864,_w_9767,_w_15819,n1526_1,_w_7059,_w_15585,n1630,_w_7396,_w_15323,n46_1,n898_1,_w_6822,_w_10112,n375_0,n1523_1,n1827_1,n1520_0,_w_9516,_w_9833,_w_9219,n1514_1,_w_13717,n479,n1433_0,n1704_1,_w_9978,N358_18,_w_11740,_w_5684,n1419_0,_w_14867,n1503_1,_w_13010,n1502_0,N188_12,_w_6700,n1496_0,n505_1,N375_15,_w_7217,n1493_1,_w_7623,_w_7541,_w_12163,n699_1,n74_1,n1221_0,_w_9539,n649_0,n1491_0,n382_1,_w_9941,_w_10995,_w_5770,_w_9227,_w_9741,_w_13179,n1487_0,n1700,_w_12753,_w_12234,n1484_0,_w_16230,_w_8197,n1482_0,_w_15187,n1056_0,_w_14989,n843_0,_w_13104,_w_10559,n771_0,n1473_0,n1323,n1883_0,n1472_0,_w_13310,n245,n1823_0,n1823_1,n1007,_w_16158,N460_0,n1463_0,_w_15979,_w_12330,_w_5841,_w_7305,_w_7654,_w_14888,_w_14004,n1554_1,N18_11,n1133_1,n1463_1,_w_8431,n1161,n945_0,n1462_1,_w_11012,_w_9071,n1457_0,n1469_0,_w_11355,n961,n1453_0,_w_13853,n1496_1,_w_7345,n1453_1,n1448_0,_w_15332,_w_10312,n1446_1,_w_13163,_w_6049,N477_17,_w_14030,n378_2,_w_9435,_w_10150,n988,_w_16137,_w_9271,n1415_0,_w_7065,_w_11218,_w_7212,n1431_1,_w_10908,n1427_0,n1475,n1425_1,n632_1,n1857_0,_w_8507,n889,n1436_0,_w_14899,_w_5487,n1416_0,n957,_w_6094,_w_8752,n1415_1,n1406_1,_w_14757,n1359_1,n1400_1,n963_1,_w_8268,n1197_0,_w_12015,n1594_1,n142,n1197_1,n751,n962_0,_w_9282,n932_0,_w_7903,n1080_0,_w_13367,_w_13327,_w_9728,n1080_1,n1549_1,n1899_0,n1899_1,n937_0,n964_0,_w_8644,_w_14215,n1013_0,n42_1,n965_0,_w_8223,n357_1,_w_7859,n965_1,n1057_1,_w_5521,n1596_0,_w_7659,n968_0,n968_1,n1836,_w_9822,n1855_1,n464,n971_1,n318,n833_1,n736_0,n736_1,_w_9378,n1250_0,n1250_1,_w_11646,_w_9325,n979_0,_w_8275,n980_0,n980_1,_w_12124,n985_0,_w_11821,n988_0,_w_7875,_w_13569,n988_1,_w_8945,_w_8978,n989_0,n989_1,_w_15498,_w_13972,_w_13931,N341_17,n1188_1,N256_0,N256_4,N256_7,N256_8,n979_1,N256_9,_w_10618,_w_6386,n296_0,N256_10,N256_11,_w_8495,N256_12,N256_13,_w_8245,N256_15,n704,N256_17,N256_20,N256_21,n1748,n902_1,_w_8621,n991_0,n992_0,_w_14422,_w_13850,n1108,n992_1,_w_7956,_w_10496,n360_1,n210,n724_0,n724_1,_w_15512,_w_13994,_w_6826,n111_0,n1001_1,_w_6288,n1006_0,_w_14220,n1006_1,_w_10277,n1007_0,_w_13694,n1007_1,_w_7908,_w_14366,_w_13009,n317_0,n1510,_w_6225,n444_1,n1379_1,n1388_0,n900,n1388_1,_w_10648,n1506,n1033_1,n33_0,_w_5795,n33_1,_w_7074,n994_0,n545_1,_w_10108,n1034_0,n1034_1,_w_15572,n1036_0,_w_14350,_w_12803,n1036_1,_w_13779,_w_13468,n1563_0,N103_14,n1550_1,_w_6110,n783_0,n1434_1,n1050_0,_w_6264,_w_10242,n1050_1,n1738_0,n1051_1,n949_0,n949_1,n1546_1,n1052_0,_w_13173,N205_15,n570_0,n570_1,n1096,n1053_0,n1750_0,n1053_1,_w_5679,_w_10058,n441_1,_w_8219,_w_9118,n1286_1,_w_12826,n261,n187_0,n1058_1,_w_15937,_w_15002,_w_12439,_w_10529,n777_1,n1059_0,n1635_0,_w_14162,_w_8014,_w_10095,_w_11176,_w_10847,n1635_1,n1558_0,_w_6730,_w_8973,_w_14516,_w_6811,N137_19,n120_0,n1064_0,_w_5374,n1064_1,n1740_0,_w_5433,n1740_1,_w_12622,_w_6257,n1066_0,_w_12689,n883_0,n1066_1,_w_15698,_w_13042,_w_10731,_w_6992,n1071_1,N1_13,_w_7071,_w_9724,_w_12252,n1698_1,n203,n59_1,_w_11483,n1077_0,n1079_1,_w_7179,N52_0,N52_3,N52_4,n414_1,N52_9,n1021_1,_w_7427,N52_10,N52_11,N52_12,_w_5512,N52_13,N52_15,N52_16,_w_10603,_w_8486,_w_9346,_w_15219,n723_0,_w_9471,_w_14906,_w_10006,_w_10836,N52_19,_w_8496,_w_13208,n1083_0,n1220_0,_w_12834,_w_5408,_w_14624,n1220_1,_w_12375,n1196_1,_w_6169,_w_14776,n753_0,n753_1,_w_6743,n1098,n1088_0,_w_5784,n103_0,n1088_1,_w_15088,_w_12635,n1158,n1015_0,n1015_1,n1357_1,_w_8708,_w_9178,n1089_0,n192,_w_7387,n857_1,_w_7838,_w_5539,n1363_0,n1092_0,_w_15048,_w_5307,n1330_0,_w_5309,_w_6794,_w_5310,_w_13709,_w_5311,_w_5315,_w_13337,_w_5317,_w_7501,_w_14120,_w_7889,_w_5318,_w_5322,_w_11659,_w_5326,_w_6818,_w_12551,n151,_w_6636,_w_5335,_w_5336,_w_5337,_w_5338,_w_15094,n90,_w_5341,_w_7749,_w_5343,_w_12659,_w_8782,_w_5344,_w_5350,_w_15223,_w_12327,n205_0,_w_5351,_w_5352,_w_7561,_w_7602,_w_5355,_w_11236,_w_5358,n854_1,_w_7279,_w_5361,_w_8008,_w_6661,_w_5364,n1842_0,_w_5365,_w_13915,_w_5366,_w_5367,_w_8582,_w_5369,_w_5371,_w_5480,_w_5372,_w_5373,_w_5375,_w_6886,_w_5379,n884_0,_w_5381,n780_0,_w_5763,_w_5382,_w_5384,_w_5386,_w_14563,_w_11456,_w_11063,n761,_w_9839,_w_6551,_w_15927,_w_5387,_w_5388,_w_5389,_w_5390,_w_13939,_w_5391,_w_11404,n1830_0,_w_9836,_w_5392,_w_5395,_w_5396,_w_8500,_w_5397,_w_7208,_w_5398,_w_10067,_w_13565,_w_12107,_w_5399,_w_9386,_w_12827,_w_5402,_w_9573,_w_5403,_w_16129,_w_6580,_w_5406,_w_10280,_w_6472,_w_6208,_w_5407,_w_16210,n589,_w_5410,_w_7425,_w_5411,_w_6139,_w_11262,_w_7382,_w_5412,_w_8661,_w_5934,N392_13,_w_5415,_w_5416,_w_16078,_w_9936,_w_10158,_w_5417,_w_8477,_w_5418,_w_7898,n1332_0,_w_5419,_w_9620,_w_5420,_w_5423,_w_5424,_w_6856,_w_5425,n130_0,_w_5427,_w_9939,_w_13724,_w_5659,_w_8761,_w_5430,_w_5434,N358_5,_w_5436,_w_12321,_w_7266,n645_1,_w_5883,_w_5438,n1815_0,_w_5440,_w_15889,n551,_w_5441,_w_6004,_w_5443,_w_7139,_w_8646,_w_5444,_w_6151,_w_9053,_w_5445,_w_5446,_w_5448,_w_6459,_w_7516,_w_5453,_w_5454,_w_5456,_w_5457,_w_5824,_w_5591,_w_7870,_w_6892,_w_10137,_w_12427,_w_6365,_w_5458,_w_8321,_w_5459,_w_6949,_w_8545,_w_5461,_w_5462,_w_5463,_w_11281,_w_5325,_w_5464,_w_7209,_w_5465,_w_10506,_w_8837,_w_12155,_w_5466,_w_14959,_w_9100,_w_13060,_w_5467,_w_5468,_w_15163,_w_5975,n1157_0,_w_5472,_w_15222,_w_12848,n838_0,_w_6150,_w_8015,_w_12485,_w_8409,_w_12794,n1873_0,_w_5474,_w_15569,_w_7221,_w_5476,_w_15530,_w_5478,_w_5481,_w_5482,_w_5485,_w_5486,_w_6060,_w_8167,_w_9904,n669,_w_5488,_w_7988,_w_9578,_w_7742,_w_5489,_w_5492,n87_0,_w_5494,_w_5496,_w_5497,_w_12201,_w_9802,_w_7572,_w_5498,_w_5607,_w_6556,_w_10905,n522_0,_w_5499,_w_5500,_w_13617,_w_5849,_w_8481,_w_9380,N69_2,_w_5503,_w_11785,_w_7150,_w_13004,_w_7215,_w_16225,_w_13020,_w_7436,_w_5506,_w_7840,_w_5799,_w_12041,_w_9875,_w_5510,_w_13882,_w_8662,n153,_w_5400,_w_5511,n899_1,_w_9837,n560,_w_5514,_w_15818,_w_7242,_w_15782,N511_19,n837,_w_5515,n361_0,_w_7489,N460_8,n1077_1,_w_9840,n482,_w_5517,_w_13935,_w_10860,_w_5518,_w_7834,_w_5524,_w_14903,_w_13857,n839,_w_9418,_w_5526,_w_5528,_w_5529,_w_13303,_w_5531,_w_6537,_w_5537,_w_12070,n116,_w_5538,_w_6320,_w_5541,_w_5544,_w_13783,_w_5547,n765_0,_w_5772,_w_5548,_w_5551,_w_8407,_w_5690,N358_1,_w_6338,_w_7177,_w_5555,n925_0,_w_5558,n180,_w_5561,_w_10332,n317,_w_5564,_w_14717,_w_9234,_w_12250,_w_5565,_w_5567,_w_15652,_w_6954,_w_7143,_w_5571,_w_10240,_w_5572,_w_15086,_w_13902,_w_8568,_w_14291,_w_11959,_w_10022,_w_7579,_w_5576,_w_13021,_w_5577,_w_5578,_w_14114,_w_5579,_w_14237,_w_13929,_w_8285,_w_13824,_w_9081,_w_5580,_w_5581,_w_6040,_w_5583,_w_5847,_w_5586,_w_11296,n1406,_w_8047,_w_10376,n620_1,_w_5587,_w_5589,_w_5596,_w_10071,_w_13598,_w_11310,_w_5597,_w_7308,_w_5599,_w_13366,_w_6672,_w_5606,n1771_0,_w_5609,_w_8016,_w_5610,_w_6800,_w_5612,n1022_0,_w_6984,_w_5615,_w_9946,_w_5618,_w_5619,_w_13575,_w_5620,_w_5523,_w_8716,_w_8391,_w_8775,_w_11510,_w_5627,_w_15860,_w_5780,n590,n1560,_w_5630,_w_15373,_w_5634,_w_5636,n983_1,_w_9067,_w_5637,_w_11862,_w_6842,_w_9810,_w_5638,_w_13637,_w_5640,n820,_w_5642,n242,n120_1,_w_7706,_w_5644,_w_5646,_w_6558,n1442_0,_w_8949,_w_7818,_w_5647,_w_5648,_w_7426,n1822,_w_5650,_w_5651,_w_7615,_w_12125,_w_8915,_w_10239,_w_5653,n408_0,_w_5654,N443_19,_w_6893,_w_11933,_w_5656,_w_14352,_w_7608,_w_6162,_w_5658,_w_7553,_w_10238,_w_5660,_w_5661,_w_13977,n1364_0,_w_5662,_w_8603,_w_5664,_w_7938,_w_5666,_w_6908,_w_9547,n682_0,_w_5670,_w_14432,_w_5671,_w_12677,_w_6076,n992,_w_5675,_w_5677,_w_11035,n442,_w_5678,_w_5680,_w_15669,_w_7138,_w_5685,_w_10938,_w_10898,_w_10874,_w_5686,_w_16131,_w_5691,_w_16196,_w_14836,_w_9174,_w_15966,n717_1,_w_9585,_w_5692,_w_14089,_w_10070,_w_5695,_w_10837,_w_9622,_w_8565,_w_5697,_w_9689,n1557_1,_w_5698,_w_13781,_w_7508,_w_8574,_w_8674,_w_5699,_w_5701,_w_9610,n1845_1,_w_5702,_w_5703,_w_11440,_w_5705,_w_9327,_w_14388,_w_9624,_w_5709,_w_5605,_w_5711,_w_8666,_w_12721,_w_6853,n1517_0,_w_8750,N358_4,_w_5713,n1182,_w_5717,_w_16267,_w_5719,_w_8162,_w_8408,_w_5720,_w_5721,_w_8557,n579_1,_w_5723,n1461,n1500_0,_w_7439,_w_5724,_w_13467,n146_1,_w_5725,_w_5726,_w_5727,_w_10546,_w_7569,n1276_1,_w_7820,_w_5728,_w_6525,n1089,_w_9018,_w_13702,_w_5730,n552_1,_w_5731,_w_12561,_w_5733,_w_5734,_w_9244,n1356_1,n1472_1,_w_5735,_w_8213,_w_9816,_w_5736,n214_0,_w_6691,_w_5738,n985_1,n789_0,_w_9598,_w_5740,_w_12562,_w_5743,_w_5744,_w_5745,_w_12980,n842_1,_w_8217,_w_5748,_w_11030,_w_10281,_w_5755,_w_10247,_w_15855,_w_5756,n163,_w_5884,_w_5757,_w_7509,_w_5758,_w_5759,_w_11336,_w_5760,_w_5761,_w_5769,n193_0,_w_5771,n730,_w_9444,_w_5773,_w_13426,_w_12682,n267_1,_w_5775,_w_9280,_w_11379,_w_5777,n910,_w_5778,_w_5779,n375,_w_5788,_w_5793,_w_12575,_w_12011,n703_0,_w_8667,_w_14616,n1047,_w_7798,_w_5794,_w_14249,n1137_1,n232,_w_5796,_w_5938,_w_14241,n282,_w_9522,_w_5797,n1804,_w_5798,_w_6592,_w_14806,_w_11707,_w_9431,_w_13969,_w_5800,_w_16215,_w_5802,_w_5801,_w_11493,_w_10993,_w_5806,_w_10388,_w_5807,_w_16216,_w_5808,_w_5811,_w_5812,_w_5814,_w_9486,_w_5815,n963,_w_5816,_w_5818,_w_14156,N494_15,_w_8184,_w_7412,n1244,n1277,_w_5822,_w_10517,_w_5825,_w_8444,_w_9039,_w_5828,_w_11085,N69_7,_w_5829,_w_14051,_w_9752,_w_5831,_w_9764,_w_6324,N171_17,_w_10204,n1852,_w_5835,_w_8654,_w_5837,_w_12737,n43_0,_w_8026,_w_12261,n1400_0,_w_5839,_w_10131,_w_10033,_w_5843,_w_5850,_w_15864,_w_6236,n60_1,_w_7934,_w_5852,n1128_0,_w_5874,_w_5853,n1735,_w_5952,_w_7091,_w_6467,_w_5854,n1575,_w_5855,_w_5856,_w_5857,_w_13443,_w_5858,N239_14,_w_5861,_w_9406,_w_14263,_w_13686,_w_9446,_w_5863,_w_15347,_w_6336,_w_5865,_w_6199,_w_5866,_w_13746,_w_5867,_w_5869,_w_11529,_w_5871,_w_13046,_w_12368,_w_5872,_w_11169,n1488_1,_w_6902,_w_8696,_w_5876,_w_15745,n1443,_w_5877,_w_15827,_w_6799,_w_5879,_w_5880,_w_5882,_w_6539,_w_10962,_w_10850,N171_18,_w_5649,_w_10244,_w_12783,n1395,_w_7224,_w_5421,_w_5885,_w_13220,_w_12810,n1110_0,_w_5886,_w_11391,_w_5888,_w_11641,_w_5889,_w_5893,_w_5790,_w_6540,_w_5894,n1573_0,_w_9420,_w_5896,n105_1,_w_5898,n606_0,_w_9112,_w_5900,_w_5903,_w_14492,_w_5904,_w_9249,_w_7500,_w_5907,n523_0,_w_9123,_w_13513,n853_0,_w_7812,_w_5908,_w_14866,n1162_1,_w_5911,_w_6701,_w_5912,n162_0,_w_5913,_w_11611,_w_5916,_w_7707,_w_5917,_w_9866,_w_5919,_w_13851,N409_17,_w_6967,_w_5920,_w_6256,_w_12639,_w_5921,_w_5543,_w_5922,n925,_w_5924,_w_8157,_w_15574,_w_7708,_w_5926,n1634_0,_w_6762,_w_5929,_w_5930,_w_11543,_w_5931,_w_10825,n1608_0,_w_6516,_w_5933,_w_13555,_w_5936,_w_5937,_w_12203,_w_5939,_w_9869,_w_5941,_w_11745,_w_9399,_w_15266,_w_5943,_w_7191,_w_14627,_w_5944,_w_7914,_w_7644,_w_5947,_w_8930,_w_5948,_w_14316,_w_11040,N460_3,_w_5953,_w_5955,_w_5956,_w_5958,_w_7099,_w_5960,_w_10930,_w_7791,_w_5965,_w_5966,n775_1,_w_8645,_w_9469,n314,_w_5971,n613,_w_5972,_w_8040,_w_5363,_w_5973,n1166_0,_w_10167,_w_5974,_w_11593,_w_5976,_w_5977,_w_8251,_w_5979,_w_11062,_w_5980,n1613,_w_5981,_w_5982,_w_5985,n1753_0,_w_6734,n792_0,_w_8187,_w_15019,_w_9684,_w_5986,_w_5987,_w_14648,_w_9795,n1661,_w_5991,_w_8977,n1620,_w_5992,_w_9049,_w_7949,n1894_0,_w_10079,_w_5999,_w_6000,N120_11,_w_6001,_w_6002,_w_11370,_w_6003,n762_1,_w_6005,_w_14521,n1357_0,_w_6006,_w_6007,n645,_w_5626,_w_6550,n298,_w_6008,_w_11752,_w_6009,_w_8992,_w_6013,_w_6860,_w_13201,_w_6014,_w_15499,_w_6016,N239_15,_w_6017,_w_12193,_w_6022,_w_6025,_w_8170,n494,_w_6026,_w_15718,_w_13244,_w_6985,_w_13488,_w_6027,_w_9778,_w_6029,_w_5475,_w_6030,_w_6031,_w_6034,n1676,_w_6035,_w_6037,N392_1,_w_6038,_w_12688,_w_6042,_w_8301,_w_6043,_w_11640,_w_6046,_w_6047,N52_18,_w_6050,_w_9515,_w_6561,_w_5360,_w_7353,_w_8656,_w_5997,_w_8979,_w_6639,_w_6056,_w_15643,_w_5906,N511_4,n408,_w_6057,_w_6058,_w_6059,_w_7783,_w_6063,_w_8352,_w_6064,n721_0,_w_8169,_w_13297,_w_5994,_w_6070,n262,_w_6371,_w_6071,n1705,_w_6075,_w_6077,_w_11227,n913_0,n1303,n496_1,_w_7922,_w_6078,_w_9473,n268,_w_6079,_w_15426,N477_6,_w_6083,_w_15744,_w_6084,_w_6086,_w_6088,_w_14262,n1286,n248,_w_6091,_w_6092,_w_6152,_w_6093,_w_6095,_w_6101,_w_6102,_w_14601,N392_6,_w_6103,_w_10606,_w_6104,_w_6105,_w_8368,_w_12481,_w_6109,_w_6112,_w_15345,_w_6114,_w_6117,_w_10021,_w_6121,n124_1,_w_9854,_w_6124,_w_15148,n1437_1,_w_6125,_w_6126,_w_6219,_w_6127,_w_6812,_w_9031,_w_6128,_w_6129,_w_6130,n1016_1,_w_6378,_w_6131,_w_8894,_w_6132,_w_7430,_w_6134,n186_1,_w_7522,_w_6136,_w_6138,_w_6140,_w_6155,_w_14320,_w_8255,_w_9524,_w_13031,n536_0,_w_6158,_w_10172,_w_6160,_w_6279,_w_8938,_w_6161,_w_6163,n478,_w_8215,_w_10111,_w_6164,n1561_1,_w_7700,_w_6168,_w_6170,n890_1,_w_6255,n1537,_w_6172,_w_11748,_w_6173,_w_11649,n265_1,_w_6174,_w_8798,_w_6177,_w_8044,_w_15089,_w_13407,_w_6178,_w_6183,_w_9132,_w_11737,_w_6184,_w_9102,_w_11196,_w_6185,_w_6187,_w_6189,_w_6190,_w_6191,_w_6196,n1211_0,_w_6202,n1529_1,_w_7634,_w_16120,n382_0,_w_6203,n336,_w_8472,_w_6206,_w_6207,_w_14417,_w_13109,_w_6210,_w_7435,_w_13697,n880_0,_w_6211,_w_6213,_w_6217,_w_6222,_w_10576,_w_9756,n532,_w_6223,_w_10929,_w_7745,_w_5473,_w_6226,_w_9158,_w_14605,_w_13312,_w_6228,_w_6238,n379,_w_7662,_w_6231,_w_6497,_w_7873,_w_6233,_w_7069,_w_6234,_w_6235,_w_6240,_w_7876,_w_6242,_w_13966,_w_6243,_w_14590,_w_5957,_w_8046,_w_6244,_w_11943,_w_6245,_w_7679,n1788_1,_w_6246,n1585_0,_w_10248,_w_13006,_w_6247,_w_6249,_w_6251,_w_6252,_w_7713,_w_8465,_w_6258,_w_6261,_w_6262,_w_11170,n117,_w_6268,_w_9740,n687_1,n308_2,_w_5878,_w_6269,_w_6271,_w_6273,_w_10521,_w_6275,N205_0,_w_5870,_w_7352,_w_9735,_w_6276,_w_6559,_w_8071,_w_13255,_w_8467,_w_8290,_w_12405,_w_9974,_w_13825,_w_7453,_w_6282,_w_6285,n370_0,_w_6286,_w_8166,_w_15883,_w_6287,_w_6289,_w_9788,_w_15963,_w_6291,_w_7577,_w_8230,n1239_0,_w_6333,_w_7068,_w_8317,_w_5750,_w_6294,N120_6,_w_6299,_w_13647,_w_6303,n1226_0,_w_6304,_w_6307,_w_6309,n595,_w_6310,_w_10602,_w_6311,_w_7105,n1370,_w_6312,_w_6313,_w_6314,_w_6315,_w_7640,_w_7604,_w_6317,_w_6533,_w_7094,_w_6318,_w_12801,_w_6319,_w_10125,n1632_1,_w_6321,_w_15454,_w_8867,_w_8899,_w_8734,_w_6323,_w_15845,_w_10868,n633_1,_w_5932,_w_6325,_w_8608,_w_9662,_w_6326,_w_9497,_w_6330,n77_0,n1121_0,_w_6332,_w_14932,_w_13334,_w_6334,_w_6337,_w_7146,_w_14092,n327_0,_w_6340,_w_9201,_w_7514,_w_6342,_w_13546,_w_5767,_w_6350,_w_12126,_w_6351,_w_6352,_w_6353,_w_12977,_w_6250,_w_6355,_w_6359,_w_14401,_w_6364,_w_16031,_w_8585,n477_0,_w_6367,_w_9947,_w_14297,_w_6368,_w_6373,_w_6369,n1072_0,_w_6370,n605,_w_9065,_w_6372,_w_6375,_w_6379,_w_7251,_w_6381,_w_8195,_w_6387,_w_16181,_w_6390,_w_13357,_w_8735,_w_6391,_w_14589,_w_6394,_w_11564,_w_6395,_w_6397,_w_15951,_w_14747,_w_6401,_w_14966,_w_12354,_w_6403,_w_10706,_w_6405,_w_7856,_w_6407,_w_9352,_w_12206,N103_13,_w_6408,_w_6409,_w_6410,_w_6220,_w_6411,_w_12916,_w_6412,_w_7216,_w_6413,_w_6415,_w_15119,_w_6418,_w_6419,_w_6420,_w_15712,_w_7433,_w_8227,_w_13438,_w_9010,_w_6423,_w_6647,_w_6427,_w_6429,_w_6430,_w_8940,_w_6432,n1824,_w_6434,n1638,_w_6436,_w_6439,_w_6680,_w_5834,_w_6440,_w_6441,_w_6442,_w_7892,_w_6444,_w_14329,_w_8976,_w_14423,n845_1,_w_6089,_w_6446,n1103,_w_6447,_w_6449,_w_14595,_w_12530,n558,_w_9163,_w_6675,_w_6451,_w_11175,_w_6452,_w_8558,_w_6455,_w_6383,_w_7517,_w_6456,_w_6461,N375_11,_w_8818,_w_14992,_w_10484,_w_6463,n614,_w_6464,_w_6465,_w_6466,_w_6469,n824_1,_w_5712,_w_6474,_w_10072,N239_13,_w_7410,_w_6478,_w_15125,_w_6481,_w_14685,_w_6483,_w_11712,_w_6484,_w_6486,_w_6488,n1191_0,_w_6489,_w_6493,n1853_1,_w_8304,_w_6494,_w_15245,_w_12253,_w_6499,_w_6500,n1237,_w_6503,_w_6504,_w_8544,_w_15893,n369,_w_6506,_w_6509,_w_6510,_w_6514,_w_6490,_w_6515,_w_15928,_w_9243,_w_6517,n953_0,_w_6518,_w_10088,_w_15100,_w_6520,_w_14062,_w_6521,n726,_w_6522,n1490_0,_w_6527,N69_12,_w_7721,_w_6529,_w_14186,_w_6530,_w_13427,_w_7341,_w_6532,_w_9094,_w_9190,_w_6536,_w_6684,_w_6543,_w_9891,_w_6546,_w_6548,_w_6553,n1732_0,n244,_w_6562,_w_8095,_w_6567,_w_6568,_w_6569,_w_9923,n695,_w_6570,_w_5810,_w_6571,_w_13868,n1590_0,_w_6624,_w_6575,_w_10915,_w_6576,_w_6577,n369_0,_w_6579,_w_7825,_w_10568,_w_6583,_w_6584,_w_6585,_w_6587,_w_15405,_w_6590,_w_10454,n1255,_w_6591,_w_10391,_w_9454,_w_6594,_w_13603,_w_6595,_w_6602,_w_6603,_w_6604,_w_6605,_w_7469,_w_9393,_w_6607,_w_13216,_w_6608,_w_6609,_w_6610,_w_13807,_w_6611,n1360_0,_w_6613,_w_6614,_w_7234,n1171,_w_6615,n1114,_w_6616,_w_11693,_w_6477,_w_6888,_w_6618,_w_11711,n188,n1174_0,_w_6619,_w_5600,_w_10085,_w_6620,N222_2,n215,_w_10205,n721,_w_6622,_w_6780,_w_6625,_w_14395,_w_6626,n1386_0,_w_6627,_w_6628,n582,_w_6629,_w_6631,_w_9743,n216_0,_w_6632,n1288_1,_w_7494,_w_7982,_w_14345,_w_10212,_w_6634,_w_6635,_w_6637,_w_14673,_w_6638,_w_6640,_w_7348,_w_5594,_w_6642,_w_6643,_w_6644,n557_0,_w_6649,_w_6652,n1439_1,_w_6655,_w_13948,n649_1,n1622_0,_w_7944,_w_6657,_w_9256,_w_6658,_w_15597,_w_6660,_w_15470,_w_14506,_w_13228,_w_8807,_w_6662,n1180,_w_6663,n967_1,n628_0,_w_6667,_w_6668,_w_13659,_w_6673,_w_8221,_w_6676,_w_7932,_w_6679,_w_11301,_w_6681,_w_11120,_w_8207,_w_11607,_w_6682,_w_7801,_w_6847,_w_6685,_w_7483,_w_6692,_w_12836,_w_6693,n1221,_w_6694,_w_6695,_w_6699,n1142_1,_w_6702,N409_2,_w_6704,n318_1,_w_6706,_w_6707,_w_15429,n1719,_w_6708,_w_7677,_w_8086,_w_10805,_w_6712,_w_8854,_w_6713,n90_0,_w_6714,N460_14,n50,_w_10230,_w_9330,_w_6715,_w_6717,_w_6719,_w_7685,_w_11263,n1509_1,_w_6720,N52_5,_w_7333,_w_6721,_w_14864,_w_6724,_w_6725,_w_9298,n1251,_w_6727,n476,_w_6729,_w_6731,_w_13881,_w_6733,_w_8889,_w_12058,_w_9489,n653,_w_6736,_w_6388,_w_6739,n666_1,_w_6740,n1282,_w_6742,_w_6747,N290_18,_w_6748,n112_0,n440_0,_w_6396,_w_6749,_w_13090,_w_5568,_w_7317,_w_6750,_w_14844,_w_9025,_w_6015,_w_6751,_w_14251,_w_6752,_w_6753,_w_6755,n971_0,_w_6758,_w_7888,_w_6453,_w_6759,_w_6761,_w_9103,_w_5328,_w_6763,_w_9478,_w_10109,_w_14502,_w_6765,_w_14674,_w_7041,_w_9048,_w_6767,_w_6768,_w_8350,_w_15167,_w_6772,_w_15032,_w_14438,_w_6774,_w_5950,_w_6645,_w_6775,n865_0,_w_6776,_w_6425,_w_8902,_w_14304,_w_9967,_w_11082,n1350_1,n684_0,_w_6777,_w_6778,_w_11278,_w_6023,_w_6779,_w_10846,_w_5432,_w_6782,N528_18,_w_6784,n554_0,_w_6785,n1744_1,n1109,_w_10047,_w_10951,_w_9499,N511_9,_w_6786,n576,n1647_1,_w_6788,_w_6792,_w_10186,_w_8588,_w_6796,_w_6646,_w_6797,_w_11144,_w_9959,_w_6802,_w_15184,_w_6272,_w_5552,_w_6803,_w_7476,n217,_w_6804,_w_12830,_w_12749,_w_6805,_w_15607,_w_6815,_w_6265,_w_7881,n1482_1,_w_6670,_w_6816,_w_6817,_w_9538,_w_6819,_w_8932,_w_6820,n1864_1,_w_6823,_w_11418,_w_6824,_w_13894,_w_8958,_w_6828,n1674,_w_6829,_w_6830,_w_6831,_w_15711,_w_6834,_w_6835,_w_6836,n756_1,_w_6837,_w_11504,n541,_w_6067,_w_6839,_w_6843,_w_11366,_w_6845,_w_9364,_w_6849,_w_6851,_w_6855,N477_9,n1656_0,n524,_w_6857,_w_6858,_w_6876,n105,_w_6859,_w_6861,_w_6959,_w_9267,_w_6862,_w_6864,_w_14136,_w_6866,_w_6867,n1527_1,_w_6868,_w_12939,_w_6869,n149_0,_w_6875,_w_8885,_w_10992,_w_6877,_w_10245,_w_6878,_w_5575,_w_9459,_w_6879,_w_8199,_w_6882,_w_11724,_w_6883,_w_8946,_w_6887,_w_6890,_w_15418,_w_6891,_w_6897,_w_14046,_w_6898,_w_8839,_w_10227,_w_6899,_w_12671,_w_6900,_w_6061,_w_6901,_w_9056,_w_6903,_w_10236,_w_7971,_w_6904,_w_6905,_w_6906,_w_8860,_w_6907,_w_6909,n1271_0,_w_6913,n871_1,_w_6914,_w_9179,_w_6919,_w_6924,_w_9205,_w_6926,_w_6929,_w_9723,_w_6931,_w_9077,_w_8277,_w_10526,n789_1,_w_6933,_w_13072,_w_6934,_w_5710,_w_6937,_w_6938,_w_6939,_w_11193,_w_6940,_w_6942,_w_6944,_w_14841,_w_6945,_w_8189,_w_15133,_w_8599,n1839,_w_6947,_w_7858,n1764_0,_w_9206,_w_6948,_w_11307,_w_6952,_w_13246,_w_6953,n989,_w_6955,_w_7624,n1546_0,_w_6956,_w_7584,_w_6961,_w_6962,_w_6963,n82,_w_6574,_w_9533,_w_9074,_w_6964,_w_8982,N494_10,_w_6965,_w_6872,_w_6968,_w_6971,_w_6974,_w_6975,_w_6976,_w_6980,_w_7170,n207_0,_w_6982,_w_6986,_w_13976,_w_7765,_w_6987,_w_6989,_w_6991,_w_6993,_w_14503,_w_6994,_w_6996,_w_6997,_w_13693,_w_7663,_w_14443,n1044,n1395_1,_w_6998,n468_1,_w_6999,_w_15817,_w_7003,_w_7006,_w_7008,_w_13288,_w_7009,n521_1,n329_1,_w_7012,_w_7014,_w_7016,_w_9542,_w_7017,_w_7018,_w_7019,_w_9660,_w_6221,_w_7021,_w_7546,_w_11777,N341_9,_w_7022,_w_14845,_w_7023,_w_7025,_w_16058,_w_7026,_w_12510,_w_8927,_w_10946,n1501,_w_7027,_w_7031,_w_7032,_w_6166,n947,_w_7033,_w_7035,_w_7458,_w_7038,_w_9140,_w_7039,_w_9248,_w_15289,_w_7596,_w_7040,_w_11596,_w_9319,n716,_w_7042,_w_7043,_w_15406,_w_6923,_w_9569,_w_14081,_w_7045,_w_10774,_w_6589,_w_10143,_w_10724,_w_10466,_w_8591,N511_11,_w_7050,_w_7052,_w_5998,_w_7054,_w_8237,_w_7771,_w_9111,_w_9980,_w_7056,_w_15144,_w_7057,_w_7060,n40_0,_w_7062,_w_7063,_w_14520,_w_7067,_w_7070,n868,_w_8602,_w_16172,_w_11767,n496,n1867_1,_w_7015,_w_7073,_w_7079,n982_1,_w_7080,n1756_0,_w_7822,n561_1,_w_6757,_w_7958,_w_6874,_w_7084,_w_7086,_w_7087,_w_7088,_w_6421,_w_9037,_w_6534,_w_7089,_w_8624,_w_10037,_w_14957,N460_11,_w_7092,_w_15374,_w_7096,_w_7372,_w_7102,n1264,_w_7106,_w_13522,_w_7108,n61,_w_7110,_w_7111,_w_14933,_w_8144,_w_9611,_w_7112,n1689_0,_w_7113,_w_13798,n75_1,_w_7114,_w_10258,_w_7115,_w_15953,_w_7118,n134,_w_7119,_w_12185,n241,_w_7123,_w_7125,_w_7127,_w_7129,_w_13817,_w_7809,_w_7136,_w_13341,_w_7142,_w_7144,_w_7145,_w_16257,_w_10193,_w_7151,_w_7498,_w_9540,_w_15171,_w_6741,_w_7154,_w_9120,_w_7156,_w_5729,_w_7157,_w_7158,_w_8703,_w_7159,_w_7160,_w_13684,_w_7162,_w_7163,_w_10770,_w_7165,n1477,_w_8897,n603,_w_7166,N290_16,_w_8463,_w_7169,n929_0,_w_7171,_w_11067,_w_9888,_w_5614,_w_7172,_w_7174,_w_7175,_w_7176,_w_13164,_w_7178,_w_10220,_w_7180,n239_0,_w_7184,_w_7187,_w_7188,_w_7195,_w_9546,_w_15128,_w_7196,_w_7198,_w_7199,_w_13003,_w_12979,_w_9789,n802_1,_w_7200,_w_13133,_w_7625,_w_5845,_w_8900,_w_7201,_w_8520,_w_7203,_w_13797,_w_7205,N273_19,_w_7206,_w_15771,_w_7207,_w_12508,_w_7210,_w_7211,_w_16002,_w_9823,_w_13191,_w_7219,_w_14946,_w_7223,_w_14462,_w_5895,_w_7226,_w_7711,_w_9518,_w_7227,_w_16206,_w_7228,_w_7229,_w_14083,_w_7230,_w_15931,_w_8298,_w_7232,n672,_w_7233,_w_14856,n1677_0,_w_7235,N222_16,_w_7237,_w_10018,n719_0,n1291,n1835,_w_7238,_w_7626,_w_6810,_w_7240,_w_7241,_w_15504,_w_7244,n854,n1146,_w_7482,_w_7246,_w_12386,_w_8372,_w_10156,_w_7248,_w_11857,_w_8433,_w_7257,_w_13913,n1858_0,_w_7258,_w_16094,_w_8680,_w_9003,_w_7260,_w_8914,_w_6051,_w_9258,_w_7264,_w_8871,n340,_w_7267,n1019,_w_7269,_w_13268,_w_7271,n964,_w_7272,_w_7276,_w_7277,n1146_0,_w_7280,_w_7281,_w_16238,_w_6298,_w_7282,_w_7285,_w_7287,_w_7288,_w_7290,_w_7293,_w_7294,_w_8287,N460_13,_w_7296,_w_7297,_w_8815,_w_7298,_w_16250,n891,_w_8523,_w_12074,_w_7299,_w_7300,_w_7306,_w_11738,_w_10175,_w_7313,_w_11165,_w_7314,_w_7315,_w_7319,_w_7324,_w_13264,_w_7449,_w_10124,_w_7325,_w_7326,_w_9210,_w_7330,_w_7335,n463_1,_w_7339,_w_13166,_w_9934,n1228,_w_7829,_w_7340,n772_1,_w_8908,n1227,_w_7342,_w_12461,_w_8556,_w_7343,_w_7344,_w_7346,_w_14419,_w_7349,_w_7351,_w_7359,_w_7360,_w_7362,_w_13012,_w_7365,_w_7366,_w_14823,_w_7368,_w_7370,_w_7371,_w_8120,_w_12958,_w_6770,_w_7374,N86_11,_w_7367,_w_7376,_w_8011,_w_14022,_w_7377,n528_0,n654,_w_7380,_w_7381,_w_7384,_w_7385,_w_7386,_w_7388,_w_7390,_w_7391,_w_14174,_w_8759,_w_8779,n341,_w_7392,_w_15677,_w_7393,_w_7394,_w_14926,_w_13396,_w_8139,n143_1,_w_8967,_w_14034,_w_7397,_w_15351,_w_7398,_w_11764,_w_7399,_w_10967,_w_7402,_w_7403,_w_9491,N358_2,_w_7404,_w_7406,n887,_w_7407,_w_7408,n646,_w_6300,_w_7612,_w_7414,n1080,_w_9054,_w_16076,_w_15735,_w_5753,_w_7415,_w_10064,_w_11733,_w_7418,_w_13534,_w_7421,_w_8297,_w_5832,_w_7422,_w_7423,_w_13956,_w_7424,_w_7899,n109,_w_7428,_w_9231,_w_7434,_w_7437,_w_13891,_w_7440,_w_7395,_w_9057,_w_7442,_w_15784,_w_12487,_w_8534,_w_7443,_w_11343,_w_7448,_w_12395,_w_7450,_w_7451,_w_7456,_w_16214,_w_16029,_w_9304,_w_7457,_w_7459,_w_8009,_w_9576,_w_7461,_w_16153,_w_14511,_w_9481,_w_13980,_w_7462,_w_7463,n55_0,n1629_1,_w_7464,_w_9308,_w_7465,_w_14963,n227,_w_7468,n542_2,_w_7470,n1688_1,_w_7478,_w_7484,_w_9965,_w_7487,_w_9781,_w_7488,_w_11801,N18_4,_w_9804,_w_6470,_w_7490,n1240,_w_7491,_w_7497,_w_14892,_w_6581,_w_7499,_w_7502,_w_12727,_w_7503,_w_7504,_w_13690,_w_7505,_w_16211,_w_8968,_w_7507,n813,_w_9425,n242_0,_w_7513,_w_7518,_w_12895,_w_10422,_w_7521,n1463,_w_7524,_w_8299,_w_16162,_w_5450,_w_7526,_w_13614,n480,_w_7527,_w_5439,_w_7528,_w_15812,_w_7529,_w_11316,_w_11288,_w_6417,_w_7530,_w_7531,_w_14947,_w_7535,_w_12049,_w_7537,_w_8452,_w_12353,_w_9315,_w_7540,_w_7542,_w_15834,_w_6424,_w_7543,_w_7549,_w_12640,_w_10767,_w_7552,_w_10407,_w_7556,_w_12231,n115_0,_w_7559,_w_7560,_w_7562,_w_8118,_w_16069,_w_7563,_w_7564,n56,_w_8699,n1653_0,_w_7565,_w_9428,_w_7566,_w_7568,_w_7570,_w_13940,_w_7573,_w_7575,_w_6538,_w_7779,_w_5964,_w_7578,_w_8853,n829_0,n927,n286_1,N103_0,_w_7582,_w_12520,_w_9692,_w_7583,_w_7588,_w_10472,_w_10233,_w_7590,_w_7591,_w_7593,_w_6722,_w_7599,_w_13941,_w_7600,_w_7601,N222_20,_w_7606,n1169_1,_w_9438,_w_7607,_w_5362,_w_7609,n1012_1,_w_7611,n509,n411_1,_w_7613,_w_11152,n320_0,n910_1,_w_7616,_w_7617,_w_8516,_w_7620,_w_7621,_w_7622,_w_16041,_w_12060,_w_7627,n238_1,n1885,_w_7628,_w_7629,_w_15938,_w_10393,n486,n449_0,_w_7630,_w_7631,_w_7632,_w_7638,_w_7639,_w_12117,_w_8313,_w_7641,_w_7643,_w_14787,_w_6012,_w_7645,_w_12365,_w_7647,_w_7648,_w_7650,_w_15180,_w_7653,_w_12890,_w_7655,_w_9013,_w_7656,_w_7657,_w_7658,_w_7665,_w_10676,_w_10485,_w_7666,_w_7667,_w_8801,_w_7668,_w_14652,n1202,_w_7669,_w_7674,_w_7304,_w_7153,_w_7675,_w_7678,_w_7093,_w_7683,_w_6541,_w_7688,_w_7689,_w_13189,_w_7690,_w_7691,_w_9228,_w_7692,n555_1,_w_7693,n415_1,_w_7694,N511_0,_w_7695,_w_7696,_w_8335,_w_7699,_w_7704,n1344_0,_w_7714,n875_1,n1293,_w_7715,n1145_0,_w_9036,n324,_w_7716,_w_7718,_w_13961,_w_8045,_w_12176,_w_7719,_w_7723,_w_10012,_w_14583,_w_7727,_w_7729,n1424_0,n184,_w_7730,_w_5707,_w_7731,_w_7411,_w_7732,_w_16154,_w_7733,_w_7751,_w_12962,_w_7735,_w_7737,_w_11686,N69_11,_w_7738,_w_13723,n162,_w_8337,_w_7739,_w_7740,_w_7746,_w_16155,_w_5786,_w_7747,n299_0,_w_7752,_w_9019,_w_15333,_w_11624,n672_0,_w_7979,_w_12776,n702,_w_9171,n1179,n1168,_w_7755,_w_7756,_w_14713,n700_1,_w_9417,_w_12338,_w_7759,_w_13923,_w_8840,_w_7760,_w_13855,_w_7181,_w_7761,_w_7764,_w_9421,_w_7766,_w_7767,_w_13993,_w_7768,_w_7770,n1431_0,_w_10210,_w_7772,N426_0,n808,_w_9101,_w_14775,n1363,_w_7774,_w_7775,n877,_w_7776,_w_8484,_w_9658,_w_7777,_w_15705,_w_8188,_w_7780,_w_7473,_w_7781,_w_7493,_w_7784,_w_15570,_w_10902,_w_7787,_w_7550,_w_7788,_w_7789,_w_7790,_w_7795,_w_7800,_w_13248,N443_12,_w_7802,_w_5910,_w_7803,_w_7806,_w_7807,_w_8390,_w_7808,n335_0,_w_7810,_w_7813,_w_15400,_w_7815,_w_9004,n1095_1,_w_7816,_w_5574,_w_7817,_w_7823,_w_9776,_w_7824,_w_5689,_w_6366,_w_7827,_w_11882,n1074_0,_w_7769,_w_7830,_w_7831,n644,_w_9202,n708,_w_7082,_w_7832,_w_15686,n1367_1,_w_7833,_w_7839,_w_14602,n1866_0,n175,_w_8742,_w_7844,n66_1,_w_7847,_w_10153,_w_7850,_w_7851,_w_7853,_w_14427,_w_7854,_w_7970,n596_0,_w_7120,_w_7701,_w_7855,_w_7861,n786_1,_w_7863,_w_15065,_w_8203,_w_7864,n1679,_w_7961,_w_7865,_w_7869,n1302,_w_7871,_w_5505,_w_7872,_w_9009,_w_8448,_w_6278,_w_7709,_w_7878,_w_8537,_w_7880,_w_7883,_w_11220,_w_10166,_w_7885,_w_7886,_w_7887,_w_5428,_w_7893,_w_7895,_w_7896,n1747_1,_w_7897,_w_9651,_w_8105,_w_10009,_w_11482,_w_7902,_w_12397,_w_10197,_w_16252,_w_14936,_w_7909,_w_14074,_w_13810,_w_13085,n502_1,_w_9720,_w_5508,_w_8072,N511_8,_w_7915,_w_16212,_w_9394,_w_7916,_w_15507,_w_9555,_w_5633,_w_7918,_w_7919,_w_8328,_w_10697,_w_7925,_w_7926,_w_7931,n289_0,_w_5553,_w_7935,_w_8636,n1059_1,_w_10001,_w_7940,n263,_w_9129,_w_7941,_w_9196,_w_7942,_w_14772,n654_0,_w_7471,_w_7076,_w_7945,_w_7946,n1076,n511,_w_7947,_w_12493,n46,_w_7948,_w_7950,_w_7951,n1844_1,_w_7952,_w_7954,_w_7955,_w_6925,_w_9153,_w_10425,_w_7959,_w_7962,n1564_0,_w_8862,_w_7964,_w_15397,_w_10711,n1561,_w_9016,_w_7966,_w_8345,n1566_0,n939_1,_w_9157,_w_7968,n451_0,_w_7972,_w_16128,_w_8091,_w_7973,n1573,_w_7974,_w_11320,_w_7976,_w_7877,_w_9952,N222_10,n1749_1,_w_7980,_w_7984,_w_8774,_w_7985,_w_9177,_w_7986,n188_0,_w_7987,_w_7989,_w_7990,_w_7993,_w_7997,_w_7998,n1148_1,_w_7999,_w_8625,_w_12858,_w_9338,_w_8000,_w_8001,_w_12966,n836_1,_w_8005,n1888,_w_8012,_w_13118,N341_1,_w_8013,_w_8017,_w_8018,_w_13079,_w_8019,_w_8020,_w_8021,_w_5342,_w_8023,_w_9873,N188_0,_w_8029,_w_9073,_w_8031,_w_8032,_w_8033,_w_10231,_w_9066,_w_9970,_w_7867,_w_8037,_w_9680,_w_8038,n450,_w_8041,n1308_0,_w_8050,_w_8053,_w_8054,_w_8676,_w_9747,_w_8059,_w_15203,_w_6871,_w_8060,_w_6599,_w_8062,_w_10921,n1401,_w_8064,_w_12140,_w_8065,N222_21,_w_5319,_w_9799,_w_8070,_w_8074,_w_8906,_w_8075,n1470,_w_7681,_w_5535,_w_8077,_w_8078,n168,_w_8270,_w_5353,_w_8079,_w_8080,_w_8081,_w_12934,_w_7077,_w_8083,n64,_w_8084,_w_6108,_w_9852,_w_10135,_w_8085,_w_6392,_w_8087,_w_14994,_w_8089,_w_15026,_w_6552,_w_8090,_w_8094,n279_0,_w_8096,_w_8099,N103_19,_w_8101,_w_8102,_w_8104,_w_15268,_w_9361,_w_9992,_w_8109,_w_6677,_w_9465,_w_8110,n1368_1,_w_8111,_w_12722,_w_8113,_w_8115,n389,_w_7506,_w_8294,n516,_w_8116,n336_0,_w_8117,N307_14,_w_8119,_w_8124,n660_0,n630,_w_9232,_w_12843,n665,_w_8129,_w_13343,_w_8130,_w_8131,_w_8133,_w_8138,_w_11041,_w_9020,_w_8140,_w_8196,_w_8142,n1365,_w_8143,n1336,_w_8146,_w_8147,_w_10141,_w_8149,n1162_0,_w_8382,_w_14325,_w_6406,_w_8151,_w_15939,_w_8153,n1216,_w_9262,_w_8156,_w_14651,_w_10338,n1505_1,_w_5954,_w_8158,_w_8159,_w_12442,_w_8491,_w_11533,_w_8160,_w_5332,_w_8161,_w_8163,_w_5522,_w_8165,_w_13846,_w_11238,_w_8171,_w_11459,n465_0,_w_8905,_w_5530,_w_8172,_w_10065,n229_1,_w_8174,_w_8175,_w_8178,_w_8181,_w_8660,_w_10107,_w_6771,_w_9827,_w_8182,_w_8185,_w_7193,_w_8190,_w_9617,_w_9666,_w_8191,_w_10665,_w_10008,_w_8198,_w_7302,n961_1,_w_8200,n1471_0,_w_8204,_w_15241,n1655,_w_8205,n1092_1,_w_8206,_w_8209,_w_9717,n1212_1,_w_10000,_w_8218,_w_8550,_w_8222,_w_8224,_w_8225,_w_8226,_w_10830,n1602_1,_w_8231,_w_8233,_w_8234,_w_8239,N324_4,n582_1,_w_8241,_w_8980,_w_7336,_w_8242,_w_8243,_w_15236,_w_15057,_w_14449,n128,_w_6281,_w_8247,_w_8248,_w_9850,_w_8249,_w_8252,_w_7036,_w_8253,_w_9695,_w_9448,_w_8254,_w_6156,_w_8737,_w_8256,_w_8257,_w_8258,_w_15543,n1716,_w_8259,_w_6194,_w_8260,_w_6678,_w_8684,_w_8263,_w_10025,_w_8264,_w_8265,_w_13080,n282_0,_w_8266,_w_7534,_w_9091,_w_7164,_w_8267,_w_8309,_w_8300,_w_5573,_w_8271,_w_8272,_w_14728,_w_8578,_w_8273,_w_8274,_w_8276,_w_14970,_w_14016,_w_8282,n1327_1,_w_8283,_w_14336,n1579_1,n1377_0,_w_8286,_w_15523,_w_13150,_w_8572,_w_13214,n1354_0,_w_7754,_w_9001,_w_9603,_w_8289,_w_9912,_w_13363,_w_13167,_w_8291,_w_8295,_w_8610,_w_8296,_w_8302,n902,_w_8303,_w_8306,_w_14796,_w_8308,_w_8314,_w_12869,_w_8318,_w_8148,_w_8418,_w_9731,_w_14984,_w_11997,_w_8320,_w_8324,_w_9453,_w_13472,_w_11746,n49,_w_9495,_w_6062,_w_8325,_w_8327,_w_8334,_w_8765,_w_8336,_w_12108,n1681_1,_w_8338,_w_15285,_w_8339,_w_12724,n1061_0,_w_6055,_w_8340,n174_0,_w_9739,n963_0,_w_8341,_w_8910,_w_15098,_w_5331,_w_8342,_w_11184,_w_5645,_w_8343,_w_10934,_w_7072,_w_8346,_w_14246,n244_0,_w_8423,_w_15116,_w_7061,_w_8347,_w_15046,_w_8981,_w_6209,_w_8348,n268_1,_w_8353,_w_9192,_w_11445,N477_11,_w_9299,n578_0,_w_8354,_w_8357,_w_9681,_w_7192,_w_8358,_w_15349,N290_7,_w_8359,N154_2,_w_8362,_w_8364,_w_10613,_w_8366,_w_7149,_w_8367,n1312_1,_w_9878,_w_8369,_w_11606,_w_9382,_w_8371,_w_8374,_w_15420,_w_9033,_w_8375,_w_8376,_w_8953,_w_8377,_w_7773,_w_10214,n1318,_w_8380,_w_9130,_w_8381,_w_10660,_w_8383,_w_6054,n1143_1,_w_8386,_w_10191,_w_8387,_w_9770,_w_8388,n725,_w_8389,_w_9734,n1373_1,N409_7,_w_10115,_w_8393,_w_9209,_w_7726,_w_8397,_w_15402,_w_8398,_w_8399,_w_9076,_w_8400,n804_1,_w_8406,n545_0,_w_8410,_w_12343,_w_11880,_w_9682,n298_0,n1230_1,_w_8414,_w_13415,_w_8419,_w_9170,_w_15460,n219_1,_w_8539,_w_8422,_w_8424,N273_14,_w_8426,n219_0,_w_8427,_w_6216,_w_8428,_w_8429,n142_1,_w_8436,_w_8440,_w_8445,n1811,_w_8446,_w_8455,_w_8457,_w_8458,n371_1,_w_8461,_w_15747,_w_5422,_w_8462,_w_8464,_w_8466,_w_8468,_w_8471,_w_8473,_w_11108,_w_8474,_w_13771,_w_8476,_w_13460,_w_8478,_w_8036,_w_8480,_w_8869,_w_9089,_w_8483,_w_8485,_w_8487,N375_5,_w_8490,_w_16270,_w_8493,_w_8494,_w_8502,n974,_w_8503,n1774_0,_w_8505,_w_15623,_w_8569,_w_15435,_w_8508,_w_8510,_w_9356,_w_10520,_w_8511,_w_12418,_w_6697,_w_8512,_w_8607,_w_8513,_w_8514,_w_13481,_w_6606,n445_1,n797,_w_8211,_w_8515,_w_8517,_w_8518,n202_1,_w_8522,_w_14577,_w_8524,_w_7254,_w_8525,_w_8528,n775_0,_w_8969,_w_8533,n548_1,_w_9173,_w_14007,_w_8536,_w_8538,_w_15364,_w_8541,_w_8542,_w_6565,_w_8547,_w_8552,n1434_0,_w_8553,_w_8554,_w_8563,_w_10076,_w_8571,n1738,_w_9514,_w_8573,_w_8576,_w_7837,_w_8577,_w_6696,n1698_0,_w_10040,_w_7431,_w_8580,_w_8581,_w_7965,_w_9697,_w_8584,_w_8589,_w_15842,_w_8351,_w_8592,n1164,_w_8594,_w_8595,_w_14581,_w_10199,_w_8596,_w_11420,_w_8597,_w_8598,N409_16,_w_8600,_w_8601,_w_8604,_w_12777,_w_8605,_w_10855,_w_8606,N290_12,_w_9501,_w_8609,_w_14905,_w_8611,_w_8612,n123,_w_8620,_w_12807,_w_8623,_w_5716,_w_8627,_w_15197,_w_6201,_w_8629,_w_8633,_w_8726,_w_8634,_w_8637,n1869_0,_w_8639,_w_8641,_w_14041,_w_8647,_w_8648,_w_9461,_w_9812,_w_14950,_w_8650,_w_8651,_w_8929,n1737,_w_8652,_w_15690,_w_13800,_w_6361,_w_8653,_w_8655,_w_6327,_w_10130,_w_8657,_w_8664,_w_8670,_w_12733,_w_9613,_w_9638,_w_8672,_w_8677,_w_8795,_w_14223,_w_8679,_w_8681,_w_8683,_w_6754,_w_7250,_w_9230,_w_12676,N239_3,_w_8686,_w_8687,_w_8689,_w_8560,_w_8690,n1570_1,_w_8692,_w_8693,_w_8694,_w_13548,_w_10709,n216_1,_w_8697,_w_13490,_w_8698,_w_9694,_w_8700,_w_14956,_w_8704,_w_9241,_w_8705,_w_8706,_w_8707,_w_16193,_w_10365,_w_6573,_w_8789,_w_9930,n1722,_w_8709,_w_8711,_w_14818,_w_9898,_w_11794,_w_8712,_w_14073,_w_7920,_w_8713,_w_9998,_w_15338,_w_8719,_w_12087,_w_8721,_w_15824,_w_13433,n149_1,_w_10264,_w_11118,_w_8723,_w_14307,n1613_0,_w_8640,_w_8725,_w_11205,n1241,_w_8727,_w_14976,_w_13206,_w_10329,n1539_0,_w_8730,_w_8731,_w_8732,n1498,_w_8740,_w_8746,_w_9927,_w_8748,n907_0,_w_6531,_w_5320,_w_8751,_w_15793,_w_8753,_w_8754,_w_8755,_w_8757,_w_8762,_w_8763,_w_8764,n1166_1,_w_8766,_w_14415,_w_8768,n1277_0,n1616_0,_w_8769,_w_13380,n72_0,_w_8771,_w_8772,_w_11043,_w_8776,_w_9046,_w_10346,_w_8777,n1625_0,_w_8890,_w_8783,_w_13315,_w_8784,_w_5437,_w_8787,n78_0,_w_8788,_w_14097,_w_8792,_w_15316,_w_8793,_w_8797,_w_8802,_w_8803,_w_8804,_w_12146,n618_1,n1404_1,_w_8810,_w_9732,_w_8811,_w_8035,_w_8812,_w_13141,_w_12413,_w_8813,_w_7321,_w_6683,_w_8501,_w_8816,n779,_w_9200,_w_8819,n821_1,n400_0,_w_8821,_w_8823,_w_8824,_w_8825,_w_8826,_w_8827,_w_10783,_w_8831,_w_8834,N52_2,_w_8835,_w_8836,_w_8838,_w_8843,_w_8844,_w_7910,_w_8845,_w_8849,_w_8850,_w_8851,_w_10229,_w_8852,_w_8856,_w_8858,_w_10633,_w_8859,_w_14362,_w_8861,n856_0,_w_9796,_w_8863,_w_10237,_w_8864,_w_8865,_w_16208,n1073_1,_w_8868,_w_6426,_w_8870,_w_6277,_w_8872,n996,_w_10100,n1832_1,_w_9530,_w_8873,_w_6917,_w_5534,_w_8874,_w_9011,n412,_w_8875,_w_8882,_w_9114,_w_8883,_w_8884,_w_10404,N409_0,n1664,_w_8886,_w_11830,n1042_1,n1766,_w_8887,_w_10370,_w_8888,_w_8893,_w_8896,_w_8901,_w_8904,_w_15749,_w_14672,_w_11099,_w_8913,n1283,_w_8100,_w_8916,_w_14999,_w_8920,_w_8921,_w_8924,N69_18,_w_8925,n569_1,_w_8928,_w_11245,_w_9384,_w_8933,_w_8935,n860,_w_8936,_w_11203,_w_8965,_w_8939,_w_14029,_w_8941,_w_8943,n73_1,_w_8948,_w_8951,_w_14254,_w_7049,_w_8955,_w_15608,_w_8956,_w_8957,_w_8963,_w_15746,_w_8970,_w_13576,n636,n1298,_w_6097,_w_8971,n1238_0,_w_8972,_w_8974,_w_14059,_w_8975,_w_11491,_w_8983,_w_8984,N494_4,_w_8985,_w_15925,N188_11,_w_8986,_w_8988,_w_14967,n271_1,N137_4,_w_8991,_w_8995,n1172_0,_w_8996,n1030_0,n408_1,_w_8998,_w_8999,_w_9005,_w_12333,_w_10891,n106,_w_9006,_w_13154,n1861_0,_w_9160,_w_9007,_w_5785,n633_0,n1266,_w_9017,_w_15917,_w_9024,_w_15959,_w_9026,_w_15692,_w_9240,_w_9027,_w_16249,_w_9028,_w_9029,_w_10444,_w_9554,_w_6157,_w_9032,_w_6328,_w_9034,_w_9337,_w_15258,_w_9035,_w_11952,_w_9041,_w_9042,_w_16110,_w_9043,_w_9047,n756_0,_w_9051,n1767,_w_9058,_w_9059,_w_9060,_w_12748,_w_11910,_w_9063,_w_5603,_w_9064,_w_7047,_w_9068,_w_9070,n1473,_w_9072,_w_16248,_w_5560,_w_9078,_w_15064,_w_9079,_w_14535,_w_13499,_w_9082,_w_14751,_w_9085,_w_9090,_w_9092,_w_9093,_w_9517,_w_9095,_w_9589,_w_9098,_w_9104,n1137_0,_w_7270,_w_7133,_w_9105,_w_9107,N86_2,_w_9108,n631_0,_w_5455,_w_9109,_w_13184,n1233_1,_w_6398,_w_9671,_w_9113,_w_9116,_w_14914,_w_7197,_w_9117,_w_7486,_w_7939,_w_9119,_w_9121,_w_15214,_w_9124,_w_6737,_w_9127,_w_15090,N426_6,_w_9131,_w_7189,_w_9133,_w_9135,_w_9357,_w_7202,_w_9136,_w_9139,_w_9141,_w_9144,_w_8176,_w_9154,_w_9156,n1242_1,_w_9159,_w_9166,_w_13055,_w_9167,n1773_0,_w_9168,_w_9792,_w_7637,_w_9169,_w_9172,n1551,_w_9175,N307_4,_w_9180,_w_9182,_w_14784,_w_13342,_w_9183,_w_5715,_w_9186,_w_9187,_w_9189,_w_12475,_w_9191,_w_9193,_w_12022,_w_9195,_w_9199,_w_14631,_w_14394,_w_7687,_w_9203,_w_13751,_w_10872,_w_6146,_w_9204,_w_9213,_w_9214,_w_9215,_w_7717,_w_7131,_w_9218,_w_12369,N460_10,N18_19,_w_9224,_w_16118,_w_11000,_w_7539,_w_9225,_w_16232,_w_9226,_w_9229,_w_9235,_w_9238,_w_9239,n1567,_w_9242,n391,_w_9245,_w_8415,_w_9246,_w_9250,_w_9253,_w_9257,_w_9263,_w_7261,_w_9264,_w_9265,_w_15085,_w_9872,n1119_0,_w_9268,N528_16,_w_9269,_w_9272,_w_11340,_w_9273,_w_9274,n375_1,_w_6880,_w_9275,_w_12887,_w_9276,_w_9277,_w_6274,_w_10226,_w_9281,_w_9285,_w_9287,_w_10099,_w_9289,_w_9526,_w_13040,n445_0,_w_9290,_w_9292,_w_14611,_w_9293,_w_8952,_w_9294,_w_10575,n1539_1,_w_9295,n1027,_w_9296,N103_10,_w_9301,n1346,_w_9302,_w_14706,_w_9303,_w_6756,_w_9305,_w_9309,_w_9310,_w_9320,_w_9322,_w_9323,_w_8262,_w_9138,_w_9326,_w_9329,_w_12655,_w_9332,_w_9339,_w_9343,_w_15708,_w_9344,_w_15031,_w_12943,n1214_0,_w_9345,_w_12952,_w_11375,n849,_w_9351,_w_13914,_w_9354,_w_9355,_w_10290,_w_9360,_w_12999,_w_9362,_w_10083,_w_9363,n124,n1567_1,_w_9365,_w_11935,_w_9366,n1161_1,_w_9367,_w_13044,_w_7024,_w_9368,_w_13584,_w_9371,_w_12618,_w_10344,_w_9373,_w_9374,_w_9434,_w_9375,_w_12611,N341_11,_w_9376,_w_10249,_w_9381,_w_11804,n1701_0,_w_9383,_w_6798,_w_9385,_w_12258,N443_1,_w_9592,_w_8876,_w_9388,_w_9391,_w_9392,_w_10073,n937_1,_w_9395,_w_9396,_w_15270,_w_9398,_w_9400,_w_9401,_w_9404,_w_9405,n691,_w_9410,_w_9412,_w_9414,_w_9416,_w_15921,_w_9422,_w_9359,_w_9423,_w_10285,_w_9426,_w_9427,_w_12371,_w_7905,_w_9437,_w_16222,_w_9439,_w_5846,_w_8361,_w_9443,_w_6389,n1752,_w_9445,_w_12932,_w_9080,_w_9493,_w_9449,_w_9452,_w_10471,_w_9456,_w_9458,_w_9460,_w_7004,_w_9462,_w_13271,_w_9466,_w_14028,_w_9467,_w_9606,_w_8479,_w_9468,_w_11955,n1671_0,_w_10062,_w_6072,_w_9470,_w_9594,_w_15728,_w_6107,_w_9474,_w_9475,_w_9476,_w_14276,_w_9477,n1694,_w_10268,_w_9480,n130,_w_6450,_w_9483,N273_5,_w_9868,n173_0,_w_9862,_w_9484,_w_9485,_w_14327,_w_9488,N154_0,_w_10219,_w_11058,_w_10627,n694_0,_w_9496,_w_7310,_w_9498,_w_14076,_w_9508,n413,_w_9510,n1200,_w_9511,n1042_0,_w_9513,n834,_w_9519,_w_5959,_w_9521,_w_9525,_w_9528,_w_9529,_w_12069,_w_9531,_w_9532,_w_9541,_w_9543,_w_13346,_w_9890,_w_9548,_w_9012,_w_9550,_w_5830,_w_9757,_w_15681,_w_9551,n1623_1,_w_6445,_w_9328,_w_9556,_w_9558,_w_9559,_w_9561,_w_11154,_w_6316,_w_9565,_w_9567,_w_12241,_w_5676,_w_5479,_w_9568,_w_15035,n1122_1,_w_9570,_w_9574,n1805_1,_w_6664,_w_9579,_w_9581,_w_14958,_w_9582,_w_11972,_w_8714,_w_9583,_w_9586,_w_9588,_w_9590,_w_9597,_w_6711,_w_9599,_w_5826,_w_9602,_w_7544,_w_9604,_w_9608,_w_9612,_w_9614,_w_10509,N171_10,n1294_1,_w_9618,_w_15535,_w_13298,_w_5380,_w_9621,_w_9623,_w_9625,_w_7347,_w_9626,_w_9844,_w_9629,_w_8385,_w_6135,_w_9631,n876,_w_9636,_w_9637,_w_9640,_w_12975,_w_9780,_w_9641,_w_6215,_w_9643,_w_9793,n947_0,n841_0,_w_8396,_w_9646,_w_9648,_w_9652,_w_9655,_w_15254,_w_12579,_w_7303,_w_9657,_w_9659,_w_10429,n323,_w_9667,_w_9668,_w_5330,n1642,_w_9672,n1887,_w_9675,_w_9509,_w_9677,_w_16167,_w_9678,_w_6669,_w_9685,_w_9686,_w_9690,_w_9693,_w_9696,_w_9698,_w_12003,N443_8,_w_9701,_w_9702,_w_9704,_w_9705,_w_9706,_w_13912,_w_9710,_w_14207,_w_11274,_w_9713,_w_9615,_w_9715,_w_9716,_w_9722,_w_9725,_w_13886,n1235_0,_w_9726,_w_9729,_w_16119,n1056_1,_w_9733,_w_9736,_w_15493,_w_9737,_w_9742,_w_9745,_w_8402,_w_9750,_w_6296,_w_9754,n1443_0,_w_9755,_w_9758,_w_5765,_w_9759,_w_9760,_w_9765,_w_9766,_w_9772,_w_9773,N409_15,_w_6885,_w_10093,_w_9779,_w_12257,_w_9785,_w_11514,_w_8039,_w_9794,_w_12358,_w_9798,n1857_1,_w_9803,_w_10588,n1508_0,_w_9805,_w_11162,_w_9806,_w_9807,_w_9808,_w_9809,n1576_1,_w_9814,_w_8841,_w_9817,_w_9818,_w_9819,_w_9820,_w_13718,_w_9824,_w_9826,_w_9828,_w_6564,_w_9834,_w_9842,_w_9843,_w_15344,n722,n568,_w_9845,_w_5875,_w_9846,_w_9847,n1384_1,_w_9849,_w_9851,_w_9534,_w_9855,N341_15,_w_9857,_w_15410,_w_9859,_w_9863,_w_14885,_w_9865,_w_16156,_w_14687,n53,_w_9867,_w_6204,_w_9870,N205_18,_w_8942,_w_9871,_w_15551,n1106_0,n220,_w_9876,n780_1,n1003_1,_w_9877,_w_9879,_w_9649,_w_9883,_w_9885,_w_9889,_w_8240,_w_6766,_w_9893,_w_9897,_w_9899,_w_9901,_w_13988,_w_5718,_w_9902,_w_9903,_w_9905,_w_7882,_w_9907,_w_9908,_w_10677,n432_0,_w_9909,_w_5349,_w_9913,_w_12095,_w_9914,_w_9915,_w_9916,_w_9450,_w_9918,_w_9924,_w_11742,_w_9928,_w_12004,_w_9929,_w_15480,n648_0,n1610_0,_w_9931,n1740,_w_9935,n1333_0,n342_1,_w_9937,n167_0,_w_9942,n1266_1,_w_9944,n1718_0,_w_9945,n1292,_w_9948,_w_14829,_w_9955,_w_9956,_w_9957,_w_9958,_w_5700,_w_9961,_w_9962,_w_12685,n1177_0,n956,_w_7000,_w_9963,n701,_w_9966,_w_5823,_w_9972,_w_10585,n1681_0,_w_9975,_w_14686,_w_9977,_w_9987,_w_9982,_w_9985,_w_9986,n1348,_w_9164,_w_9988,_w_15416,_w_11081,n1538_1,_w_9989,_w_9990,_w_9993,_w_7126,_w_9994,_w_9152,_w_9995,_w_9996,_w_9999,_w_10003,_w_10004,_w_14814,_w_6181,_w_10007,n1072,_w_10011,n1224,_w_10013,_w_15113,_w_10014,_w_14593,_w_10015,_w_11976,_w_9964,n336_1,_w_10016,_w_10019,_w_10023,_w_10026,_w_10030,_w_10031,_w_13416,_w_13278,_w_10032,_w_10035,_w_10041,_w_10042,_w_10494,_w_10044,_w_10046,_w_10049,_w_10050,_w_7671,_w_10054,_w_14298,_w_10055,_w_10057,_w_10059,_w_10060,n591_1,N256_5,_w_10063,_w_10066,_w_13589,_w_10717,n1678_0,_w_10068,_w_10069,_w_13437,_w_10075,_w_7538,_w_10086,_w_10087,_w_10094,_w_13277,_w_9861,n261_0,_w_10096,_w_9777,n1441,_w_10097,n659,_w_10098,_w_10102,_w_14782,_w_7311,_w_10105,_w_10106,_w_15563,_w_7400,_w_10110,_w_10113,_w_10114,_w_10116,_w_10118,_w_9719,_w_10120,n952,_w_10121,n627_0,_w_10126,n1718,n173_1,_w_10127,N256_16,_w_9523,_w_9050,_w_10128,_w_10129,N103_3,_w_10133,_w_10136,n1152,_w_8499,_w_10139,_w_10140,_w_15269,_w_10144,_w_10145,_w_10146,_w_13041,_w_10148,_w_14045,_w_10151,_w_10152,_w_10159,_w_10160,_w_11171,_w_10162,_w_6384,_w_10165,n699_0,n156_1,_w_10168,_w_10169,n1829,_w_6053,_w_10170,_w_10171,N443_11,_w_9557,_w_10176,_w_10178,_w_15121,N307_15,_w_10179,_w_10181,_w_10184,_w_10187,_w_14170,_w_10189,_w_10190,_w_10194,_w_14514,_w_10195,_w_15848,_w_11715,_w_10196,_w_10200,_w_10201,_w_10202,_w_14487,_w_13382,_w_9512,_w_6113,_w_5590,_w_10208,_w_10209,_w_10211,_w_11655,_w_10213,_w_10215,_w_7046,_w_10216,_w_10217,_w_10218,_w_10223,_w_10225,_w_7904,_w_10228,n726_0,_w_10241,_w_10246,_w_14065,_w_8210,_w_10250,_w_14879,N120_9,_w_10251,_w_10255,n255,_w_10259,_w_10261,_w_10270,_w_5340,_w_5764,_w_10272;

  bfr _b_14386(.a(N86),.q(_w_16288));
  bfr _b_14385(.a(N69),.q(_w_16287));
  bfr _b_14384(.a(_w_16286),.q(_w_16198));
  bfr _b_14380(.a(_w_16282),.q(_w_16283));
  bfr _b_14379(.a(_w_16281),.q(_w_16282));
  bfr _b_14377(.a(_w_16279),.q(_w_16280));
  bfr _b_14374(.a(_w_16276),.q(_w_16277));
  bfr _b_14372(.a(_w_16274),.q(_w_16275));
  bfr _b_14367(.a(_w_16269),.q(_w_16270));
  bfr _b_14364(.a(_w_16266),.q(_w_16267));
  bfr _b_14363(.a(_w_16265),.q(_w_16266));
  bfr _b_14362(.a(_w_16264),.q(_w_16265));
  bfr _b_14360(.a(_w_16262),.q(_w_16263));
  bfr _b_14359(.a(_w_16261),.q(_w_16262));
  bfr _b_14358(.a(_w_16260),.q(_w_16261));
  bfr _b_14355(.a(_w_16257),.q(_w_16258));
  bfr _b_14354(.a(_w_16256),.q(_w_16257));
  bfr _b_14350(.a(_w_16252),.q(_w_16253));
  bfr _b_14345(.a(_w_16247),.q(_w_16248));
  bfr _b_14344(.a(_w_16246),.q(_w_16247));
  bfr _b_14337(.a(_w_16239),.q(_w_16240));
  bfr _b_14336(.a(_w_16238),.q(_w_16239));
  bfr _b_14335(.a(_w_16237),.q(_w_16238));
  bfr _b_14334(.a(_w_16236),.q(_w_16237));
  bfr _b_14332(.a(_w_16234),.q(_w_16235));
  bfr _b_14331(.a(_w_16233),.q(_w_16234));
  bfr _b_14330(.a(_w_16232),.q(_w_16233));
  bfr _b_14329(.a(_w_16231),.q(_w_16232));
  bfr _b_14327(.a(_w_16229),.q(_w_16230));
  bfr _b_14325(.a(_w_16227),.q(_w_16228));
  bfr _b_14324(.a(_w_16226),.q(_w_16227));
  bfr _b_14320(.a(_w_16222),.q(_w_16223));
  bfr _b_14319(.a(_w_16221),.q(_w_16222));
  bfr _b_14318(.a(_w_16220),.q(_w_16221));
  bfr _b_14317(.a(_w_16219),.q(_w_16220));
  bfr _b_14316(.a(_w_16218),.q(_w_16219));
  bfr _b_14313(.a(_w_16215),.q(_w_16216));
  bfr _b_14310(.a(_w_16212),.q(_w_16213));
  bfr _b_14308(.a(_w_16210),.q(_w_16211));
  bfr _b_14307(.a(_w_16209),.q(_w_16210));
  bfr _b_14306(.a(_w_16208),.q(_w_16209));
  bfr _b_14303(.a(_w_16205),.q(_w_16206));
  bfr _b_14301(.a(_w_16203),.q(_w_16204));
  bfr _b_14298(.a(_w_16200),.q(_w_16201));
  bfr _b_14297(.a(_w_16199),.q(_w_16200));
  bfr _b_14296(.a(N528),.q(_w_16199));
  bfr _b_14293(.a(_w_16195),.q(_w_16196));
  bfr _b_14291(.a(_w_16193),.q(_w_16194));
  bfr _b_14290(.a(_w_16192),.q(_w_16193));
  bfr _b_14287(.a(_w_16189),.q(_w_16190));
  bfr _b_14285(.a(_w_16187),.q(_w_16188));
  bfr _b_14283(.a(_w_16185),.q(_w_16186));
  bfr _b_14280(.a(_w_16182),.q(_w_16183));
  bfr _b_14277(.a(_w_16179),.q(_w_16180));
  bfr _b_14276(.a(_w_16178),.q(_w_16179));
  bfr _b_14274(.a(_w_16176),.q(_w_16177));
  bfr _b_14273(.a(_w_16175),.q(_w_16176));
  bfr _b_14269(.a(_w_16171),.q(_w_16172));
  bfr _b_14265(.a(_w_16167),.q(_w_16168));
  bfr _b_14264(.a(_w_16166),.q(_w_16167));
  bfr _b_14262(.a(_w_16164),.q(_w_16165));
  bfr _b_14261(.a(_w_16163),.q(_w_16164));
  bfr _b_14257(.a(_w_16159),.q(_w_16160));
  bfr _b_14256(.a(_w_16158),.q(_w_16159));
  bfr _b_14255(.a(_w_16157),.q(_w_16158));
  bfr _b_14254(.a(_w_16156),.q(_w_16157));
  bfr _b_14250(.a(_w_16152),.q(_w_16153));
  bfr _b_14247(.a(_w_16149),.q(_w_16150));
  bfr _b_14246(.a(_w_16148),.q(_w_16149));
  bfr _b_14244(.a(_w_16146),.q(_w_16147));
  bfr _b_14243(.a(_w_16145),.q(_w_16146));
  bfr _b_14242(.a(_w_16144),.q(_w_16145));
  bfr _b_14240(.a(_w_16142),.q(_w_16143));
  bfr _b_14239(.a(_w_16141),.q(_w_16142));
  bfr _b_14237(.a(_w_16139),.q(_w_16140));
  bfr _b_14236(.a(_w_16138),.q(_w_16139));
  bfr _b_14233(.a(_w_16135),.q(_w_16136));
  bfr _b_14231(.a(_w_16133),.q(_w_16134));
  bfr _b_14226(.a(_w_16128),.q(_w_16129));
  bfr _b_14221(.a(_w_16123),.q(_w_16124));
  bfr _b_14217(.a(_w_16119),.q(_w_16120));
  bfr _b_14214(.a(_w_16116),.q(_w_16117));
  bfr _b_14213(.a(_w_16115),.q(_w_16116));
  bfr _b_14212(.a(_w_16114),.q(_w_16115));
  bfr _b_14208(.a(_w_16110),.q(_w_16111));
  bfr _b_14328(.a(_w_16230),.q(_w_16231));
  bfr _b_14207(.a(_w_16109),.q(_w_16110));
  bfr _b_14201(.a(_w_16103),.q(_w_16104));
  bfr _b_14200(.a(_w_16102),.q(_w_16103));
  bfr _b_14198(.a(_w_16100),.q(_w_16101));
  bfr _b_14196(.a(_w_16098),.q(_w_16099));
  bfr _b_14195(.a(_w_16097),.q(_w_16098));
  bfr _b_14192(.a(_w_16094),.q(_w_16095));
  bfr _b_14188(.a(_w_16090),.q(_w_16091));
  bfr _b_14184(.a(_w_16086),.q(_w_16087));
  bfr _b_14182(.a(_w_16084),.q(_w_16085));
  bfr _b_14181(.a(_w_16083),.q(_w_16084));
  bfr _b_14180(.a(_w_16082),.q(_w_16083));
  bfr _b_14179(.a(_w_16081),.q(_w_16082));
  bfr _b_14176(.a(_w_16078),.q(_w_16079));
  bfr _b_14175(.a(_w_16077),.q(_w_16078));
  bfr _b_14174(.a(_w_16076),.q(_w_16077));
  bfr _b_14171(.a(_w_16073),.q(_w_16074));
  bfr _b_14168(.a(_w_16070),.q(_w_16071));
  bfr _b_14166(.a(_w_16068),.q(_w_16069));
  bfr _b_14165(.a(_w_16067),.q(_w_16068));
  bfr _b_14260(.a(_w_16162),.q(_w_16163));
  bfr _b_14162(.a(_w_16064),.q(_w_16065));
  bfr _b_14160(.a(_w_16062),.q(_w_16063));
  bfr _b_14158(.a(_w_16060),.q(_w_16061));
  bfr _b_14156(.a(_w_16058),.q(_w_16059));
  bfr _b_14155(.a(_w_16057),.q(_w_16058));
  bfr _b_14154(.a(_w_16056),.q(_w_16057));
  bfr _b_14153(.a(_w_16055),.q(_w_16056));
  bfr _b_14150(.a(_w_16052),.q(_w_16053));
  bfr _b_14147(.a(_w_16049),.q(_w_16050));
  bfr _b_14146(.a(_w_16048),.q(_w_16049));
  bfr _b_14143(.a(_w_16045),.q(_w_16046));
  bfr _b_14142(.a(_w_16044),.q(_w_16045));
  bfr _b_14141(.a(_w_16043),.q(_w_16044));
  bfr _b_14140(.a(_w_16042),.q(_w_16043));
  bfr _b_14137(.a(_w_16039),.q(_w_16040));
  bfr _b_14136(.a(_w_16038),.q(_w_16039));
  bfr _b_14135(.a(_w_16037),.q(_w_16038));
  bfr _b_14133(.a(_w_16035),.q(_w_16036));
  bfr _b_14131(.a(_w_16033),.q(_w_16034));
  bfr _b_14130(.a(_w_16032),.q(_w_16033));
  bfr _b_14128(.a(_w_16030),.q(_w_16031));
  bfr _b_14125(.a(_w_16027),.q(_w_16028));
  bfr _b_14122(.a(_w_16024),.q(_w_16025));
  bfr _b_14121(.a(_w_16023),.q(_w_16024));
  bfr _b_14120(.a(_w_16022),.q(_w_16023));
  bfr _b_14119(.a(_w_16021),.q(_w_16022));
  bfr _b_14117(.a(N494),.q(_w_16020));
  bfr _b_14116(.a(_w_16018),.q(_w_15930));
  bfr _b_14114(.a(_w_16016),.q(_w_16017));
  bfr _b_14113(.a(_w_16015),.q(_w_16016));
  bfr _b_14112(.a(_w_16014),.q(_w_16015));
  bfr _b_14111(.a(_w_16013),.q(_w_16014));
  bfr _b_14110(.a(_w_16012),.q(_w_16013));
  bfr _b_14109(.a(_w_16011),.q(_w_16012));
  bfr _b_14108(.a(_w_16010),.q(_w_16011));
  bfr _b_14103(.a(_w_16005),.q(_w_16006));
  bfr _b_14102(.a(_w_16004),.q(_w_16005));
  bfr _b_14101(.a(_w_16003),.q(_w_16004));
  bfr _b_14099(.a(_w_16001),.q(_w_16002));
  bfr _b_14098(.a(_w_16000),.q(_w_16001));
  bfr _b_14097(.a(_w_15999),.q(_w_16000));
  bfr _b_14096(.a(_w_15998),.q(_w_15999));
  bfr _b_14093(.a(_w_15995),.q(_w_15996));
  bfr _b_14092(.a(_w_15994),.q(_w_15995));
  bfr _b_14090(.a(_w_15992),.q(_w_15993));
  bfr _b_14089(.a(_w_15991),.q(_w_15992));
  bfr _b_14086(.a(_w_15988),.q(_w_15989));
  bfr _b_14082(.a(_w_15984),.q(_w_15985));
  bfr _b_14080(.a(_w_15982),.q(_w_15983));
  bfr _b_14079(.a(_w_15981),.q(_w_15982));
  bfr _b_14078(.a(_w_15980),.q(_w_15981));
  bfr _b_14076(.a(_w_15978),.q(_w_15979));
  bfr _b_14073(.a(_w_15975),.q(_w_15976));
  bfr _b_14071(.a(_w_15973),.q(_w_15974));
  bfr _b_14067(.a(_w_15969),.q(_w_15970));
  bfr _b_14064(.a(_w_15966),.q(_w_15967));
  bfr _b_14063(.a(_w_15965),.q(_w_15966));
  bfr _b_14062(.a(_w_15964),.q(_w_15965));
  bfr _b_14060(.a(_w_15962),.q(_w_15963));
  bfr _b_14059(.a(_w_15961),.q(_w_15962));
  bfr _b_14057(.a(_w_15959),.q(_w_15960));
  bfr _b_14048(.a(_w_15950),.q(_w_15951));
  bfr _b_14046(.a(_w_15948),.q(_w_15949));
  bfr _b_14044(.a(_w_15946),.q(_w_15947));
  bfr _b_14043(.a(_w_15945),.q(_w_15946));
  bfr _b_14042(.a(_w_15944),.q(_w_15945));
  bfr _b_14041(.a(_w_15943),.q(_w_15944));
  bfr _b_14040(.a(_w_15942),.q(_w_15943));
  bfr _b_14038(.a(_w_15940),.q(_w_15941));
  bfr _b_14036(.a(_w_15938),.q(_w_15939));
  bfr _b_14030(.a(_w_15932),.q(_w_15933));
  bfr _b_14029(.a(_w_15931),.q(_w_15932));
  bfr _b_14027(.a(_w_15929),.q(_w_15861));
  bfr _b_14025(.a(_w_15927),.q(_w_15928));
  bfr _b_14023(.a(_w_15925),.q(_w_15926));
  bfr _b_14022(.a(_w_15924),.q(_w_15925));
  bfr _b_14020(.a(_w_15922),.q(_w_15923));
  bfr _b_14015(.a(_w_15917),.q(_w_15918));
  bfr _b_14013(.a(_w_15915),.q(_w_15916));
  bfr _b_14010(.a(_w_15912),.q(_w_15913));
  bfr _b_14008(.a(_w_15910),.q(_w_15911));
  bfr _b_14007(.a(_w_15909),.q(_w_15910));
  bfr _b_14006(.a(_w_15908),.q(_w_15909));
  bfr _b_14004(.a(_w_15906),.q(_w_15907));
  bfr _b_14002(.a(_w_15904),.q(_w_15905));
  bfr _b_13996(.a(_w_15898),.q(_w_15899));
  bfr _b_13995(.a(_w_15897),.q(_w_15898));
  bfr _b_13993(.a(_w_15895),.q(_w_15896));
  bfr _b_13991(.a(_w_15893),.q(_w_15894));
  bfr _b_13989(.a(_w_15891),.q(_w_15892));
  bfr _b_13984(.a(_w_15886),.q(_w_15887));
  bfr _b_13983(.a(_w_15885),.q(_w_15886));
  bfr _b_13982(.a(_w_15884),.q(_w_15885));
  bfr _b_13977(.a(_w_15879),.q(_w_15880));
  bfr _b_13975(.a(_w_15877),.q(_w_15878));
  bfr _b_13973(.a(_w_15875),.q(_w_15876));
  bfr _b_13972(.a(_w_15874),.q(_w_15875));
  bfr _b_13970(.a(_w_15872),.q(_w_15873));
  bfr _b_13968(.a(_w_15870),.q(_w_15871));
  bfr _b_13967(.a(_w_15869),.q(_w_15870));
  bfr _b_13966(.a(_w_15868),.q(_w_15869));
  bfr _b_13964(.a(_w_15866),.q(_w_15867));
  bfr _b_13963(.a(_w_15865),.q(_w_15866));
  bfr _b_13962(.a(_w_15864),.q(_w_15865));
  bfr _b_13961(.a(_w_15863),.q(_w_15864));
  bfr _b_13959(.a(N460),.q(_w_15862));
  bfr _b_13957(.a(_w_15859),.q(_w_15860));
  bfr _b_13956(.a(_w_15858),.q(_w_15859));
  bfr _b_13953(.a(_w_15855),.q(_w_15856));
  bfr _b_13952(.a(_w_15854),.q(_w_15855));
  bfr _b_13951(.a(_w_15853),.q(_w_15854));
  bfr _b_13950(.a(_w_15852),.q(_w_15853));
  bfr _b_13948(.a(_w_15850),.q(_w_15851));
  bfr _b_13947(.a(_w_15849),.q(_w_15850));
  bfr _b_13945(.a(_w_15847),.q(_w_15848));
  bfr _b_13944(.a(_w_15846),.q(_w_15847));
  bfr _b_13942(.a(_w_15844),.q(_w_15845));
  bfr _b_13941(.a(_w_15843),.q(_w_15844));
  bfr _b_13940(.a(_w_15842),.q(_w_15843));
  bfr _b_13939(.a(_w_15841),.q(_w_15842));
  bfr _b_13938(.a(_w_15840),.q(_w_15841));
  bfr _b_13936(.a(_w_15838),.q(_w_15839));
  bfr _b_13934(.a(_w_15836),.q(_w_15837));
  bfr _b_13933(.a(_w_15835),.q(_w_15836));
  bfr _b_13932(.a(_w_15834),.q(_w_15835));
  bfr _b_13930(.a(_w_15832),.q(_w_15833));
  bfr _b_13929(.a(_w_15831),.q(_w_15832));
  bfr _b_13926(.a(_w_15828),.q(_w_15829));
  bfr _b_13924(.a(_w_15826),.q(_w_15827));
  bfr _b_13921(.a(_w_15823),.q(_w_15824));
  bfr _b_14129(.a(_w_16031),.q(_w_16032));
  bfr _b_14069(.a(_w_15971),.q(_w_15972));
  bfr _b_13920(.a(_w_15822),.q(_w_15823));
  bfr _b_13917(.a(_w_15819),.q(_w_15820));
  bfr _b_13916(.a(_w_15818),.q(_w_15819));
  bfr _b_13915(.a(_w_15817),.q(_w_15818));
  bfr _b_13911(.a(_w_15813),.q(_w_15814));
  bfr _b_13909(.a(_w_15811),.q(_w_15812));
  bfr _b_13904(.a(_w_15806),.q(_w_15807));
  bfr _b_13902(.a(_w_15804),.q(_w_15805));
  bfr _b_13899(.a(_w_15801),.q(_w_15802));
  bfr _b_13897(.a(_w_15799),.q(_w_15800));
  bfr _b_13895(.a(_w_15797),.q(_w_15798));
  bfr _b_13891(.a(_w_15793),.q(_w_15794));
  bfr _b_13890(.a(N443),.q(_w_15793));
  bfr _b_13887(.a(_w_15789),.q(_w_15790));
  bfr _b_13886(.a(_w_15788),.q(_w_15789));
  bfr _b_13885(.a(_w_15787),.q(_w_15788));
  bfr _b_13884(.a(_w_15786),.q(_w_15787));
  bfr _b_13883(.a(_w_15785),.q(_w_15786));
  bfr _b_13882(.a(_w_15784),.q(_w_15785));
  bfr _b_13881(.a(_w_15783),.q(_w_15784));
  bfr _b_13880(.a(_w_15782),.q(_w_15783));
  bfr _b_13879(.a(_w_15781),.q(_w_15782));
  bfr _b_13878(.a(_w_15780),.q(_w_15781));
  bfr _b_13877(.a(_w_15779),.q(_w_15780));
  bfr _b_13876(.a(_w_15778),.q(_w_15779));
  bfr _b_13874(.a(_w_15776),.q(_w_15777));
  bfr _b_13873(.a(_w_15775),.q(_w_15776));
  bfr _b_13871(.a(_w_15773),.q(_w_15774));
  bfr _b_13869(.a(_w_15771),.q(_w_15772));
  bfr _b_13865(.a(_w_15767),.q(_w_15768));
  bfr _b_13862(.a(_w_15764),.q(_w_15765));
  bfr _b_13861(.a(_w_15763),.q(_w_15764));
  bfr _b_13859(.a(_w_15761),.q(_w_15762));
  bfr _b_13858(.a(_w_15760),.q(_w_15761));
  bfr _b_13857(.a(_w_15759),.q(_w_15760));
  bfr _b_13855(.a(_w_15757),.q(_w_15758));
  bfr _b_13854(.a(_w_15756),.q(_w_15757));
  bfr _b_13853(.a(_w_15755),.q(_w_15756));
  bfr _b_13851(.a(_w_15753),.q(_w_15754));
  bfr _b_13849(.a(_w_15751),.q(_w_15752));
  bfr _b_13848(.a(_w_15750),.q(_w_15751));
  bfr _b_13847(.a(_w_15749),.q(_w_15750));
  bfr _b_13843(.a(_w_15745),.q(_w_15746));
  bfr _b_13842(.a(_w_15744),.q(_w_15745));
  bfr _b_13840(.a(_w_15742),.q(_w_15743));
  bfr _b_13838(.a(_w_15740),.q(_w_15741));
  bfr _b_13837(.a(_w_15739),.q(_w_15740));
  bfr _b_13835(.a(_w_15737),.q(_w_15738));
  bfr _b_14163(.a(_w_16065),.q(_w_16066));
  bfr _b_13833(.a(_w_15735),.q(_w_15736));
  bfr _b_13830(.a(_w_15732),.q(_w_15733));
  bfr _b_13829(.a(_w_15731),.q(_w_15732));
  bfr _b_13825(.a(N426),.q(_w_15728));
  bfr _b_13823(.a(_w_15725),.q(_w_15726));
  bfr _b_13822(.a(_w_15724),.q(_w_15725));
  bfr _b_13819(.a(_w_15721),.q(_w_15722));
  bfr _b_13813(.a(_w_15715),.q(_w_15716));
  bfr _b_13811(.a(_w_15713),.q(_w_15714));
  bfr _b_13810(.a(_w_15712),.q(_w_15713));
  bfr _b_13807(.a(_w_15709),.q(_w_15710));
  bfr _b_13806(.a(_w_15708),.q(_w_15709));
  bfr _b_13804(.a(_w_15706),.q(_w_15707));
  bfr _b_13803(.a(_w_15705),.q(_w_15706));
  bfr _b_13802(.a(_w_15704),.q(_w_15705));
  bfr _b_13801(.a(_w_15703),.q(_w_15704));
  bfr _b_13800(.a(_w_15702),.q(_w_15703));
  bfr _b_13796(.a(_w_15698),.q(_w_15699));
  bfr _b_13794(.a(_w_15696),.q(_w_15697));
  bfr _b_13793(.a(_w_15695),.q(_w_15696));
  bfr _b_13792(.a(_w_15694),.q(_w_15695));
  bfr _b_13787(.a(_w_15689),.q(_w_15690));
  bfr _b_13786(.a(_w_15688),.q(_w_15689));
  bfr _b_13785(.a(_w_15687),.q(_w_15688));
  bfr _b_13784(.a(_w_15686),.q(_w_15687));
  bfr _b_13782(.a(_w_15684),.q(_w_15685));
  bfr _b_13781(.a(_w_15683),.q(_w_15684));
  bfr _b_13780(.a(_w_15682),.q(_w_15683));
  bfr _b_13777(.a(_w_15679),.q(_w_15680));
  bfr _b_13776(.a(_w_15678),.q(_w_15679));
  bfr _b_13772(.a(_w_15674),.q(_w_15675));
  bfr _b_13771(.a(_w_15673),.q(_w_15674));
  bfr _b_13770(.a(_w_15672),.q(_w_15673));
  bfr _b_13769(.a(_w_15671),.q(_w_15672));
  bfr _b_13765(.a(_w_15667),.q(_w_15668));
  bfr _b_13762(.a(_w_15664),.q(_w_15665));
  bfr _b_13760(.a(_w_15662),.q(_w_15663));
  bfr _b_13757(.a(_w_15659),.q(_w_15660));
  bfr _b_13753(.a(_w_15655),.q(_w_15656));
  bfr _b_13751(.a(_w_15653),.q(_w_15654));
  bfr _b_13748(.a(_w_15650),.q(_w_15651));
  bfr _b_13747(.a(_w_15649),.q(_w_15650));
  bfr _b_13746(.a(_w_15648),.q(_w_15649));
  bfr _b_13745(.a(_w_15647),.q(_w_15648));
  bfr _b_13744(.a(_w_15646),.q(_w_15647));
  bfr _b_13743(.a(_w_15645),.q(_w_15646));
  bfr _b_13739(.a(_w_15641),.q(_w_15642));
  bfr _b_13738(.a(_w_15640),.q(_w_15641));
  bfr _b_13737(.a(_w_15639),.q(_w_15640));
  bfr _b_13736(.a(_w_15638),.q(_w_15639));
  bfr _b_14203(.a(_w_16105),.q(_w_16106));
  bfr _b_13731(.a(_w_15633),.q(_w_15634));
  bfr _b_13730(.a(_w_15632),.q(_w_15633));
  bfr _b_13729(.a(_w_15631),.q(_w_15632));
  bfr _b_13728(.a(_w_15630),.q(_w_15631));
  bfr _b_13727(.a(_w_15629),.q(_w_15630));
  bfr _b_13726(.a(_w_15628),.q(_w_15629));
  bfr _b_13724(.a(_w_15626),.q(_w_15627));
  bfr _b_13723(.a(_w_15625),.q(_w_15626));
  bfr _b_13722(.a(_w_15624),.q(_w_15625));
  bfr _b_13721(.a(_w_15623),.q(_w_15624));
  bfr _b_13719(.a(N392),.q(_w_15622));
  bfr _b_13717(.a(_w_15619),.q(_w_15620));
  bfr _b_13716(.a(_w_15618),.q(_w_15619));
  bfr _b_13715(.a(_w_15617),.q(_w_15618));
  bfr _b_13714(.a(_w_15616),.q(_w_15617));
  bfr _b_13711(.a(_w_15613),.q(_w_15614));
  bfr _b_13709(.a(_w_15611),.q(_w_15612));
  bfr _b_13708(.a(_w_15610),.q(_w_15611));
  bfr _b_13707(.a(_w_15609),.q(_w_15610));
  bfr _b_13705(.a(_w_15607),.q(_w_15608));
  bfr _b_13702(.a(_w_15604),.q(_w_15605));
  bfr _b_13701(.a(_w_15603),.q(_w_15604));
  bfr _b_13697(.a(_w_15599),.q(_w_15600));
  bfr _b_13696(.a(_w_15598),.q(_w_15599));
  bfr _b_13695(.a(_w_15597),.q(_w_15598));
  bfr _b_13694(.a(N375),.q(_w_15597));
  bfr _b_13692(.a(_w_15594),.q(_w_15595));
  bfr _b_13691(.a(_w_15593),.q(_w_15594));
  bfr _b_13689(.a(_w_15591),.q(_w_15592));
  bfr _b_13688(.a(_w_15590),.q(_w_15591));
  bfr _b_13686(.a(_w_15588),.q(_w_15589));
  bfr _b_13683(.a(_w_15585),.q(_w_15586));
  bfr _b_13682(.a(_w_15584),.q(_w_15585));
  bfr _b_13681(.a(_w_15583),.q(_w_15584));
  bfr _b_13680(.a(_w_15582),.q(_w_15583));
  bfr _b_14031(.a(_w_15933),.q(_w_15934));
  bfr _b_13679(.a(_w_15581),.q(_w_15582));
  bfr _b_13677(.a(_w_15579),.q(_w_15580));
  bfr _b_13676(.a(_w_15578),.q(_w_15579));
  bfr _b_13673(.a(_w_15575),.q(_w_15576));
  bfr _b_13668(.a(N35),.q(_w_15570));
  bfr _b_13664(.a(_w_15566),.q(_w_15567));
  bfr _b_13663(.a(_w_15565),.q(_w_15566));
  bfr _b_13662(.a(_w_15564),.q(_w_15565));
  bfr _b_13658(.a(_w_15560),.q(_w_15561));
  bfr _b_13657(.a(_w_15559),.q(_w_15560));
  bfr _b_13655(.a(_w_15557),.q(_w_15558));
  bfr _b_13647(.a(_w_15549),.q(_w_15550));
  bfr _b_13645(.a(_w_15547),.q(_w_15548));
  bfr _b_13642(.a(_w_15544),.q(_w_15542));
  bfr _b_13638(.a(_w_15540),.q(_w_15541));
  bfr _b_13637(.a(N307),.q(_w_15540));
  bfr _b_13635(.a(N273),.q(_w_15537));
  bfr _b_13634(.a(_w_15536),.q(_w_15534));
  bfr _b_13633(.a(_w_15535),.q(_w_15536));
  bfr _b_13631(.a(N239),.q(_w_15533));
  bfr _b_13630(.a(N205),.q(_w_15532));
  bfr _b_13628(.a(N18),.q(_w_15530));
  bfr _b_13625(.a(N137),.q(_w_15527));
  bfr _b_13623(.a(N103),.q(_w_15525));
  bfr _b_13905(.a(_w_15807),.q(_w_15808));
  bfr _b_13621(.a(_w_15523),.q(_w_15524));
  bfr _b_13620(.a(N1),.q(_w_15523));
  bfr _b_13619(.a(_w_15521),.q(n779));
  bfr _b_13618(.a(_w_15520),.q(N18_15));
  bfr _b_13617(.a(_w_15519),.q(_w_15520));
  bfr _b_13616(.a(_w_15518),.q(_w_15519));
  bfr _b_13615(.a(_w_15517),.q(_w_15518));
  bfr _b_13613(.a(_w_15515),.q(_w_15516));
  bfr _b_13611(.a(_w_15513),.q(_w_15514));
  bfr _b_13605(.a(_w_15507),.q(_w_15508));
  bfr _b_13604(.a(_w_15506),.q(_w_15507));
  bfr _b_14210(.a(_w_16112),.q(_w_16113));
  bfr _b_13602(.a(_w_15504),.q(_w_15505));
  bfr _b_13600(.a(_w_15502),.q(_w_15503));
  bfr _b_13599(.a(_w_15501),.q(_w_15502));
  bfr _b_13597(.a(_w_15499),.q(_w_15500));
  bfr _b_13596(.a(_w_15498),.q(_w_15499));
  bfr _b_13594(.a(_w_15496),.q(N18_13));
  bfr _b_13593(.a(_w_15495),.q(_w_15496));
  bfr _b_13592(.a(_w_15494),.q(_w_15495));
  bfr _b_13591(.a(_w_15493),.q(_w_15494));
  bfr _b_13587(.a(_w_15489),.q(_w_15490));
  bfr _b_13585(.a(_w_15487),.q(_w_15488));
  bfr _b_13584(.a(_w_15486),.q(N18_6));
  bfr _b_13582(.a(_w_15484),.q(N18_3));
  bfr _b_13579(.a(_w_15481),.q(_w_15482));
  bfr _b_13577(.a(_w_15479),.q(_w_15480));
  bfr _b_13574(.a(_w_15476),.q(_w_15477));
  bfr _b_13573(.a(_w_15475),.q(_w_15476));
  bfr _b_13571(.a(_w_15473),.q(_w_15474));
  bfr _b_13566(.a(_w_15468),.q(_w_15469));
  bfr _b_13564(.a(_w_15466),.q(_w_15467));
  bfr _b_13563(.a(_w_15465),.q(_w_15466));
  bfr _b_13562(.a(_w_15464),.q(_w_15465));
  bfr _b_13561(.a(_w_15463),.q(_w_15464));
  bfr _b_13560(.a(_w_15462),.q(_w_15463));
  bfr _b_13559(.a(_w_15461),.q(_w_15462));
  bfr _b_13558(.a(_w_15460),.q(_w_15461));
  bfr _b_13556(.a(_w_15458),.q(_w_15459));
  bfr _b_13553(.a(_w_15455),.q(_w_15456));
  bfr _b_13551(.a(_w_15453),.q(_w_15454));
  bfr _b_13546(.a(_w_15448),.q(_w_15449));
  bfr _b_13544(.a(_w_15446),.q(_w_15447));
  bfr _b_13542(.a(_w_15444),.q(_w_15445));
  bfr _b_13541(.a(_w_15443),.q(_w_15444));
  bfr _b_13539(.a(_w_15441),.q(_w_15442));
  bfr _b_13538(.a(_w_15440),.q(_w_15441));
  bfr _b_13537(.a(_w_15439),.q(_w_15440));
  bfr _b_13536(.a(_w_15438),.q(_w_15439));
  bfr _b_13535(.a(_w_15437),.q(_w_15438));
  bfr _b_13534(.a(_w_15436),.q(_w_15437));
  bfr _b_13532(.a(_w_15434),.q(_w_15435));
  bfr _b_13529(.a(_w_15431),.q(_w_15432));
  bfr _b_13528(.a(_w_15430),.q(_w_15431));
  bfr _b_13527(.a(_w_15429),.q(_w_15430));
  bfr _b_13526(.a(_w_15428),.q(_w_15429));
  bfr _b_13524(.a(_w_15426),.q(_w_15427));
  bfr _b_13523(.a(_w_15425),.q(_w_15426));
  bfr _b_13522(.a(_w_15424),.q(_w_15425));
  bfr _b_13521(.a(_w_15423),.q(_w_15424));
  bfr _b_13519(.a(_w_15421),.q(_w_15422));
  bfr _b_13518(.a(_w_15420),.q(_w_15421));
  bfr _b_13517(.a(_w_15419),.q(_w_15420));
  bfr _b_13513(.a(_w_15415),.q(_w_15416));
  bfr _b_13508(.a(_w_15410),.q(_w_15411));
  bfr _b_13507(.a(_w_15409),.q(_w_15410));
  bfr _b_13504(.a(_w_15406),.q(_w_15407));
  bfr _b_13500(.a(_w_15402),.q(_w_15403));
  bfr _b_13497(.a(_w_15399),.q(_w_15400));
  bfr _b_13496(.a(_w_15398),.q(_w_15399));
  bfr _b_13494(.a(_w_15396),.q(N18_2));
  bfr _b_13492(.a(_w_15394),.q(_w_15395));
  bfr _b_13491(.a(_w_15393),.q(_w_15394));
  bfr _b_13712(.a(_w_15614),.q(_w_15615));
  bfr _b_13489(.a(_w_15391),.q(_w_15392));
  bfr _b_13486(.a(_w_15388),.q(_w_15389));
  bfr _b_13485(.a(_w_15387),.q(_w_15388));
  bfr _b_13788(.a(_w_15690),.q(_w_15691));
  bfr _b_13483(.a(_w_15385),.q(_w_15386));
  bfr _b_13480(.a(_w_15382),.q(_w_15383));
  bfr _b_13479(.a(_w_15381),.q(_w_15382));
  bfr _b_13478(.a(_w_15380),.q(_w_15381));
  bfr _b_13476(.a(_w_15378),.q(_w_15379));
  bfr _b_13471(.a(_w_15373),.q(_w_15374));
  bfr _b_13470(.a(_w_15372),.q(_w_15373));
  bfr _b_13468(.a(_w_15370),.q(_w_15371));
  bfr _b_13467(.a(_w_15369),.q(_w_15370));
  bfr _b_13699(.a(_w_15601),.q(_w_15602));
  bfr _b_13466(.a(_w_15368),.q(_w_15369));
  bfr _b_13465(.a(_w_15367),.q(_w_15368));
  bfr _b_13464(.a(_w_15366),.q(_w_15367));
  bfr _b_13463(.a(_w_15365),.q(_w_15366));
  bfr _b_13461(.a(_w_15363),.q(_w_15364));
  bfr _b_13456(.a(_w_15358),.q(_w_15359));
  bfr _b_13455(.a(_w_15357),.q(_w_15358));
  bfr _b_13453(.a(_w_15355),.q(_w_15356));
  bfr _b_13872(.a(_w_15774),.q(_w_15775));
  bfr _b_13448(.a(_w_15350),.q(_w_15351));
  bfr _b_13447(.a(_w_15349),.q(_w_15350));
  bfr _b_13445(.a(_w_15347),.q(_w_15348));
  bfr _b_13444(.a(_w_15346),.q(_w_15347));
  bfr _b_13443(.a(_w_15345),.q(_w_15346));
  bfr _b_13441(.a(_w_15343),.q(_w_15344));
  bfr _b_13440(.a(_w_15342),.q(_w_15343));
  bfr _b_13439(.a(_w_15341),.q(_w_15342));
  bfr _b_13438(.a(_w_15340),.q(N18_1));
  bfr _b_13437(.a(_w_15339),.q(_w_15340));
  bfr _b_13815(.a(_w_15717),.q(_w_15718));
  bfr _b_13434(.a(_w_15336),.q(_w_15337));
  bfr _b_13433(.a(_w_15335),.q(_w_15336));
  bfr _b_13432(.a(_w_15334),.q(_w_15335));
  bfr _b_13429(.a(_w_15331),.q(_w_15332));
  bfr _b_13426(.a(_w_15328),.q(_w_15329));
  bfr _b_13422(.a(_w_15324),.q(_w_15325));
  bfr _b_13421(.a(_w_15323),.q(_w_15324));
  bfr _b_13419(.a(_w_15321),.q(_w_15322));
  bfr _b_13416(.a(_w_15318),.q(_w_15319));
  bfr _b_13415(.a(_w_15317),.q(_w_15318));
  bfr _b_13412(.a(_w_15314),.q(_w_15315));
  bfr _b_13404(.a(_w_15306),.q(_w_15307));
  bfr _b_13402(.a(_w_15304),.q(n422));
  bfr _b_13398(.a(_w_15300),.q(_w_15301));
  bfr _b_13395(.a(_w_15297),.q(n56_1));
  bfr _b_13394(.a(_w_15296),.q(_w_15297));
  bfr _b_13925(.a(_w_15827),.q(_w_15828));
  bfr _b_13392(.a(_w_15294),.q(n1143_1));
  bfr _b_13391(.a(_w_15293),.q(_w_15294));
  bfr _b_13390(.a(_w_15292),.q(_w_15293));
  bfr _b_13389(.a(_w_15291),.q(_w_15292));
  bfr _b_13388(.a(_w_15290),.q(N69_3));
  bfr _b_13386(.a(_w_15288),.q(_w_15289));
  bfr _b_13385(.a(_w_15287),.q(_w_15288));
  bfr _b_13383(.a(_w_15285),.q(_w_15286));
  bfr _b_13382(.a(_w_15284),.q(_w_15285));
  bfr _b_13380(.a(_w_15282),.q(_w_15283));
  bfr _b_13379(.a(_w_15281),.q(_w_15282));
  bfr _b_13378(.a(_w_15280),.q(_w_15281));
  bfr _b_13377(.a(_w_15279),.q(_w_15280));
  bfr _b_13376(.a(_w_15278),.q(_w_15279));
  bfr _b_13373(.a(_w_15275),.q(_w_15276));
  bfr _b_13372(.a(_w_15274),.q(_w_15275));
  bfr _b_13371(.a(_w_15273),.q(_w_15274));
  bfr _b_13370(.a(_w_15272),.q(_w_15273));
  bfr _b_13369(.a(_w_15271),.q(_w_15272));
  bfr _b_13368(.a(_w_15270),.q(_w_15271));
  bfr _b_13366(.a(_w_15268),.q(_w_15269));
  bfr _b_13361(.a(_w_15263),.q(_w_15264));
  bfr _b_13360(.a(_w_15262),.q(_w_15263));
  bfr _b_13358(.a(_w_15260),.q(_w_15261));
  bfr _b_13354(.a(_w_15256),.q(_w_15257));
  bfr _b_13351(.a(_w_15253),.q(_w_15254));
  bfr _b_13350(.a(_w_15252),.q(_w_15253));
  bfr _b_13346(.a(_w_15248),.q(_w_15249));
  bfr _b_13343(.a(_w_15245),.q(_w_15246));
  bfr _b_13342(.a(_w_15244),.q(_w_15245));
  bfr _b_13341(.a(_w_15243),.q(_w_15244));
  bfr _b_13340(.a(_w_15242),.q(_w_15243));
  bfr _b_13335(.a(_w_15237),.q(_w_15238));
  bfr _b_13332(.a(_w_15234),.q(_w_15235));
  bfr _b_13330(.a(_w_15232),.q(_w_15233));
  bfr _b_13327(.a(_w_15229),.q(_w_15230));
  bfr _b_13326(.a(_w_15228),.q(_w_15229));
  bfr _b_13325(.a(_w_15227),.q(_w_15228));
  bfr _b_13324(.a(_w_15226),.q(_w_15227));
  bfr _b_13323(.a(_w_15225),.q(_w_15226));
  bfr _b_13319(.a(_w_15221),.q(_w_15222));
  bfr _b_13318(.a(_w_15220),.q(_w_15221));
  bfr _b_13316(.a(_w_15218),.q(_w_15219));
  bfr _b_13312(.a(_w_15214),.q(_w_15215));
  bfr _b_13311(.a(_w_15213),.q(_w_15214));
  bfr _b_13308(.a(_w_15210),.q(_w_15211));
  bfr _b_13303(.a(_w_15205),.q(_w_15206));
  bfr _b_13302(.a(_w_15204),.q(_w_15205));
  bfr _b_13300(.a(_w_15202),.q(N69_2));
  bfr _b_13299(.a(_w_15201),.q(_w_15202));
  bfr _b_13292(.a(_w_15194),.q(_w_15195));
  bfr _b_13288(.a(_w_15190),.q(_w_15191));
  bfr _b_13287(.a(_w_15189),.q(_w_15190));
  bfr _b_13282(.a(_w_15184),.q(_w_15185));
  bfr _b_13281(.a(_w_15183),.q(_w_15184));
  bfr _b_13279(.a(_w_15181),.q(_w_15182));
  bfr _b_13277(.a(_w_15179),.q(_w_15180));
  bfr _b_14191(.a(_w_16093),.q(_w_16094));
  bfr _b_13276(.a(_w_15178),.q(_w_15179));
  bfr _b_13275(.a(_w_15177),.q(_w_15178));
  bfr _b_13274(.a(_w_15176),.q(_w_15177));
  bfr _b_13271(.a(_w_15173),.q(_w_15174));
  bfr _b_13270(.a(_w_15172),.q(_w_15173));
  bfr _b_13267(.a(_w_15169),.q(_w_15170));
  bfr _b_13265(.a(_w_15167),.q(_w_15168));
  bfr _b_13263(.a(_w_15165),.q(_w_15166));
  bfr _b_13261(.a(_w_15163),.q(_w_15164));
  bfr _b_13260(.a(_w_15162),.q(_w_15163));
  bfr _b_13259(.a(_w_15161),.q(_w_15162));
  bfr _b_13257(.a(_w_15159),.q(_w_15160));
  bfr _b_13253(.a(_w_15155),.q(_w_15156));
  bfr _b_13252(.a(_w_15154),.q(_w_15155));
  bfr _b_13251(.a(_w_15153),.q(_w_15154));
  bfr _b_13248(.a(_w_15150),.q(_w_15151));
  bfr _b_13247(.a(_w_15149),.q(_w_15150));
  bfr _b_13246(.a(_w_15148),.q(_w_15149));
  bfr _b_13985(.a(_w_15887),.q(_w_15888));
  bfr _b_13245(.a(_w_15147),.q(_w_15148));
  bfr _b_13244(.a(_w_15146),.q(N69_1));
  bfr _b_13242(.a(_w_15144),.q(_w_15145));
  bfr _b_13240(.a(_w_15142),.q(_w_15143));
  bfr _b_13239(.a(_w_15141),.q(_w_15142));
  bfr _b_13238(.a(_w_15140),.q(_w_15141));
  bfr _b_13236(.a(_w_15138),.q(_w_15139));
  bfr _b_13234(.a(_w_15136),.q(_w_15137));
  bfr _b_13233(.a(_w_15135),.q(_w_15136));
  bfr _b_13232(.a(_w_15134),.q(_w_15135));
  bfr _b_13230(.a(_w_15132),.q(_w_15133));
  bfr _b_13229(.a(_w_15131),.q(_w_15132));
  bfr _b_13228(.a(_w_15130),.q(_w_15131));
  bfr _b_13227(.a(_w_15129),.q(_w_15130));
  bfr _b_13225(.a(_w_15127),.q(_w_15128));
  bfr _b_13224(.a(_w_15126),.q(_w_15127));
  bfr _b_13442(.a(_w_15344),.q(_w_15345));
  bfr _b_13222(.a(_w_15124),.q(_w_15125));
  bfr _b_13221(.a(_w_15123),.q(_w_15124));
  bfr _b_13220(.a(_w_15122),.q(n652_1));
  bfr _b_13219(.a(_w_15121),.q(_w_15122));
  bfr _b_13217(.a(_w_15119),.q(_w_15120));
  bfr _b_13216(.a(_w_15118),.q(n808_1));
  bfr _b_13215(.a(_w_15117),.q(_w_15118));
  bfr _b_13214(.a(_w_15116),.q(_w_15117));
  bfr _b_13213(.a(_w_15115),.q(_w_15116));
  bfr _b_13211(.a(_w_15113),.q(n1212_1));
  bfr _b_13799(.a(_w_15701),.q(_w_15702));
  bfr _b_13210(.a(_w_15112),.q(_w_15113));
  bfr _b_13209(.a(_w_15111),.q(_w_15112));
  bfr _b_13208(.a(_w_15110),.q(_w_15111));
  bfr _b_13207(.a(_w_15109),.q(n410));
  bfr _b_13206(.a(_w_15108),.q(n1248_1));
  bfr _b_13205(.a(_w_15107),.q(_w_15108));
  bfr _b_13204(.a(_w_15106),.q(_w_15107));
  bfr _b_13202(.a(_w_15104),.q(n1260_1));
  bfr _b_13200(.a(_w_15102),.q(_w_15103));
  bfr _b_13199(.a(_w_15101),.q(_w_15102));
  bfr _b_13197(.a(_w_15099),.q(_w_15100));
  bfr _b_13196(.a(_w_15098),.q(_w_15099));
  bfr _b_13193(.a(_w_15095),.q(_w_15096));
  bfr _b_13192(.a(_w_15094),.q(_w_15095));
  bfr _b_13191(.a(_w_15093),.q(_w_15094));
  bfr _b_13187(.a(_w_15089),.q(_w_15090));
  bfr _b_13185(.a(_w_15087),.q(_w_15088));
  bfr _b_13184(.a(_w_15086),.q(_w_15087));
  bfr _b_13183(.a(_w_15085),.q(_w_15086));
  bfr _b_13182(.a(_w_15084),.q(n1345_1));
  bfr _b_13181(.a(_w_15083),.q(_w_15084));
  bfr _b_13180(.a(_w_15082),.q(_w_15083));
  bfr _b_13178(.a(_w_15080),.q(n92));
  bfr _b_13177(.a(_w_15079),.q(n1788_1));
  bfr _b_13176(.a(_w_15078),.q(_w_15079));
  bfr _b_13173(.a(_w_15075),.q(n1155_1));
  bfr _b_13171(.a(_w_15073),.q(_w_15074));
  bfr _b_13170(.a(_w_15072),.q(_w_15073));
  bfr _b_13168(.a(_w_15070),.q(n1386_1));
  bfr _b_13167(.a(_w_15069),.q(_w_15070));
  bfr _b_13166(.a(_w_15068),.q(_w_15069));
  bfr _b_13165(.a(_w_15067),.q(_w_15068));
  bfr _b_13164(.a(_w_15066),.q(n476));
  bfr _b_13163(.a(_w_15065),.q(n1416_1));
  bfr _b_13162(.a(_w_15064),.q(_w_15065));
  bfr _b_13161(.a(_w_15063),.q(_w_15064));
  bfr _b_13160(.a(_w_15062),.q(_w_15063));
  bfr _b_13159(.a(_w_15061),.q(n1422_1));
  bfr _b_13157(.a(_w_15059),.q(_w_15060));
  bfr _b_13155(.a(_w_15057),.q(n1198));
  bfr _b_13153(.a(_w_15055),.q(_w_15056));
  bfr _b_13626(.a(N154),.q(_w_15528));
  bfr _b_13151(.a(_w_15053),.q(_w_15054));
  bfr _b_13678(.a(_w_15580),.q(_w_15581));
  bfr _b_13149(.a(_w_15051),.q(n1491_1));
  bfr _b_13148(.a(_w_15050),.q(_w_15051));
  bfr _b_13146(.a(_w_15048),.q(_w_15049));
  bfr _b_13144(.a(_w_15046),.q(_w_15047));
  bfr _b_13137(.a(_w_15039),.q(n236));
  bfr _b_13136(.a(_w_15038),.q(_w_15039));
  bfr _b_13133(.a(_w_15035),.q(_w_15036));
  bfr _b_13128(.a(_w_15030),.q(_w_15031));
  bfr _b_13127(.a(_w_15029),.q(_w_15030));
  bfr _b_13124(.a(_w_15026),.q(_w_15027));
  bfr _b_13121(.a(_w_15023),.q(n1503_1));
  bfr _b_13116(.a(_w_15018),.q(n1722_1));
  bfr _b_13113(.a(_w_15015),.q(_w_15016));
  bfr _b_13111(.a(_w_15013),.q(_w_15014));
  bfr _b_13108(.a(_w_15010),.q(n1107_1));
  bfr _b_13107(.a(_w_15009),.q(_w_15010));
  bfr _b_13106(.a(_w_15008),.q(_w_15009));
  bfr _b_13104(.a(_w_15006),.q(n485));
  bfr _b_13103(.a(_w_15005),.q(n1665_1));
  bfr _b_13102(.a(_w_15004),.q(_w_15005));
  bfr _b_13100(.a(_w_15002),.q(_w_15003));
  bfr _b_13099(.a(_w_15001),.q(n1444));
  bfr _b_13098(.a(_w_15000),.q(n436));
  bfr _b_14321(.a(_w_16223),.q(_w_16224));
  bfr _b_13097(.a(_w_14999),.q(_w_15000));
  bfr _b_13096(.a(_w_14998),.q(_w_14999));
  bfr _b_13095(.a(_w_14997),.q(_w_14998));
  bfr _b_13094(.a(_w_14996),.q(_w_14997));
  bfr _b_13758(.a(_w_15660),.q(_w_15661));
  bfr _b_13091(.a(_w_14993),.q(_w_14994));
  bfr _b_13090(.a(_w_14992),.q(_w_14993));
  bfr _b_13088(.a(_w_14990),.q(_w_14991));
  bfr _b_13086(.a(_w_14988),.q(n1539));
  bfr _b_13085(.a(_w_14987),.q(_w_14988));
  bfr _b_13083(.a(_w_14985),.q(_w_14986));
  bfr _b_13082(.a(_w_14984),.q(_w_14985));
  bfr _b_13081(.a(_w_14983),.q(_w_14984));
  bfr _b_13074(.a(_w_14976),.q(n1753_1));
  bfr _b_13073(.a(_w_14975),.q(_w_14976));
  bfr _b_13072(.a(_w_14974),.q(_w_14975));
  bfr _b_13071(.a(_w_14973),.q(_w_14974));
  bfr _b_13070(.a(_w_14972),.q(n1765_1));
  bfr _b_13068(.a(_w_14970),.q(_w_14971));
  bfr _b_13067(.a(_w_14969),.q(_w_14970));
  bfr _b_13064(.a(_w_14966),.q(_w_14967));
  bfr _b_13061(.a(_w_14963),.q(_w_14964));
  bfr _b_13060(.a(_w_14962),.q(_w_14963));
  bfr _b_13059(.a(_w_14961),.q(_w_14962));
  bfr _b_13056(.a(_w_14958),.q(_w_14959));
  bfr _b_13065(.a(_w_14967),.q(n1357));
  bfr _b_13055(.a(_w_14957),.q(_w_14958));
  bfr _b_13053(.a(_w_14955),.q(n1794_1));
  bfr _b_13052(.a(_w_14954),.q(_w_14955));
  bfr _b_13051(.a(_w_14953),.q(_w_14954));
  bfr _b_13050(.a(_w_14952),.q(_w_14953));
  bfr _b_13049(.a(_w_14951),.q(n1589));
  bfr _b_13047(.a(_w_14949),.q(_w_14950));
  bfr _b_13045(.a(_w_14947),.q(_w_14948));
  bfr _b_13040(.a(_w_14942),.q(n1895_1));
  bfr _b_13037(.a(_w_14939),.q(_w_14940));
  bfr _b_13036(.a(_w_14938),.q(n1901));
  bfr _b_13035(.a(_w_14937),.q(n1897));
  bfr _b_13034(.a(_w_14936),.q(_w_14937));
  bfr _b_13032(.a(_w_14934),.q(_w_14935));
  bfr _b_13031(.a(_w_14933),.q(_w_14934));
  bfr _b_13029(.a(_w_14931),.q(_w_14932));
  bfr _b_13028(.a(_w_14930),.q(_w_14931));
  bfr _b_13026(.a(_w_14928),.q(_w_14929));
  bfr _b_13024(.a(_w_14926),.q(_w_14927));
  bfr _b_13022(.a(_w_14924),.q(_w_14925));
  bfr _b_13021(.a(_w_14923),.q(_w_14924));
  bfr _b_13020(.a(_w_14922),.q(_w_14923));
  bfr _b_13019(.a(_w_14921),.q(_w_14922));
  bfr _b_13018(.a(_w_14920),.q(_w_14921));
  bfr _b_13016(.a(_w_14918),.q(_w_14919));
  bfr _b_13014(.a(_w_14916),.q(_w_14917));
  bfr _b_13010(.a(_w_14912),.q(_w_14913));
  bfr _b_13009(.a(_w_14911),.q(_w_14912));
  bfr _b_13007(.a(_w_14909),.q(_w_14910));
  bfr _b_13005(.a(_w_14907),.q(_w_14908));
  bfr _b_13003(.a(_w_14905),.q(_w_14906));
  bfr _b_13000(.a(_w_14902),.q(_w_14903));
  bfr _b_12997(.a(_w_14899),.q(_w_14900));
  bfr _b_12996(.a(_w_14898),.q(_w_14899));
  bfr _b_12995(.a(_w_14897),.q(_w_14898));
  bfr _b_12992(.a(_w_14894),.q(_w_14895));
  bfr _b_14342(.a(_w_16244),.q(_w_16245));
  bfr _b_12990(.a(_w_14892),.q(_w_14893));
  bfr _b_12988(.a(_w_14890),.q(_w_14891));
  bfr _b_12987(.a(_w_14889),.q(_w_14890));
  bfr _b_13805(.a(_w_15707),.q(_w_15708));
  bfr _b_12986(.a(_w_14888),.q(_w_14889));
  bfr _b_12984(.a(_w_14886),.q(_w_14887));
  bfr _b_12983(.a(_w_14885),.q(_w_14886));
  bfr _b_12982(.a(_w_14884),.q(n1895));
  bfr _b_12978(.a(_w_14880),.q(_w_14881));
  bfr _b_12977(.a(_w_14879),.q(_w_14880));
  bfr _b_12975(.a(_w_14877),.q(_w_14878));
  bfr _b_12974(.a(_w_14876),.q(_w_14877));
  bfr _b_12973(.a(_w_14875),.q(_w_14876));
  bfr _b_12972(.a(_w_14874),.q(_w_14875));
  bfr _b_12970(.a(_w_14872),.q(_w_14873));
  bfr _b_12968(.a(_w_14870),.q(_w_14871));
  bfr _b_12967(.a(_w_14869),.q(_w_14870));
  bfr _b_12965(.a(_w_14867),.q(_w_14868));
  bfr _b_12963(.a(_w_14865),.q(_w_14866));
  bfr _b_12962(.a(_w_14864),.q(_w_14865));
  bfr _b_12961(.a(_w_14863),.q(_w_14864));
  bfr _b_12960(.a(_w_14862),.q(_w_14863));
  bfr _b_12957(.a(_w_14859),.q(_w_14860));
  bfr _b_12956(.a(_w_14858),.q(_w_14859));
  bfr _b_12955(.a(_w_14857),.q(_w_14858));
  bfr _b_12954(.a(_w_14856),.q(_w_14857));
  bfr _b_12953(.a(_w_14855),.q(_w_14856));
  bfr _b_12951(.a(_w_14853),.q(_w_14854));
  bfr _b_12950(.a(_w_14852),.q(_w_14853));
  bfr _b_12945(.a(_w_14847),.q(_w_14848));
  bfr _b_12939(.a(_w_14841),.q(_w_14842));
  bfr _b_12937(.a(_w_14839),.q(_w_14840));
  bfr _b_12936(.a(_w_14838),.q(_w_14839));
  bfr _b_12935(.a(_w_14837),.q(_w_14838));
  bfr _b_12934(.a(_w_14836),.q(_w_14837));
  bfr _b_12933(.a(_w_14835),.q(_w_14836));
  bfr _b_12931(.a(_w_14833),.q(_w_14834));
  bfr _b_13610(.a(_w_15512),.q(_w_15513));
  bfr _b_12930(.a(_w_14832),.q(n542_2));
  bfr _b_13867(.a(_w_15769),.q(_w_15770));
  bfr _b_12929(.a(_w_14831),.q(_w_14832));
  bfr _b_14185(.a(_w_16087),.q(_w_16088));
  bfr _b_12926(.a(_w_14828),.q(N6280));
  bfr _b_12924(.a(_w_14826),.q(_w_14827));
  bfr _b_12922(.a(_w_14824),.q(n1411));
  bfr _b_12921(.a(_w_14823),.q(n1888));
  bfr _b_12920(.a(_w_14822),.q(n438));
  bfr _b_12917(.a(_w_14819),.q(_w_14820));
  bfr _b_12916(.a(_w_14818),.q(n1886));
  bfr _b_12915(.a(_w_14817),.q(_w_14818));
  bfr _b_12914(.a(_w_14816),.q(_w_14817));
  bfr _b_12913(.a(_w_14815),.q(_w_14816));
  bfr _b_12912(.a(_w_14814),.q(_w_14815));
  bfr _b_12911(.a(_w_14813),.q(_w_14814));
  bfr _b_12909(.a(_w_14811),.q(_w_14812));
  bfr _b_12907(.a(_w_14809),.q(_w_14810));
  bfr _b_12906(.a(_w_14808),.q(_w_14809));
  bfr _b_12905(.a(_w_14807),.q(_w_14808));
  bfr _b_12904(.a(_w_14806),.q(_w_14807));
  bfr _b_12903(.a(_w_14805),.q(_w_14806));
  bfr _b_12901(.a(_w_14803),.q(_w_14804));
  bfr _b_12900(.a(_w_14802),.q(_w_14803));
  bfr _b_12899(.a(_w_14801),.q(_w_14802));
  bfr _b_12898(.a(_w_14800),.q(_w_14801));
  bfr _b_12892(.a(_w_14794),.q(_w_14795));
  bfr _b_12891(.a(_w_14793),.q(_w_14794));
  bfr _b_12890(.a(_w_14792),.q(_w_14793));
  bfr _b_12888(.a(_w_14790),.q(_w_14791));
  bfr _b_12887(.a(_w_14789),.q(_w_14790));
  bfr _b_12884(.a(_w_14786),.q(_w_14787));
  bfr _b_12883(.a(_w_14785),.q(_w_14786));
  bfr _b_12940(.a(_w_14842),.q(_w_14843));
  bfr _b_12881(.a(_w_14783),.q(_w_14784));
  bfr _b_12880(.a(_w_14782),.q(_w_14783));
  bfr _b_12874(.a(_w_14776),.q(_w_14777));
  bfr _b_12873(.a(_w_14775),.q(_w_14776));
  bfr _b_12870(.a(_w_14772),.q(_w_14773));
  bfr _b_12869(.a(_w_14771),.q(_w_14772));
  bfr _b_12867(.a(_w_14769),.q(n1882));
  bfr _b_12866(.a(_w_14768),.q(n1576_1));
  bfr _b_12865(.a(_w_14767),.q(_w_14768));
  bfr _b_12864(.a(_w_14766),.q(_w_14767));
  bfr _b_12863(.a(_w_14765),.q(_w_14766));
  bfr _b_12861(.a(_w_14763),.q(_w_14764));
  bfr _b_12860(.a(_w_14762),.q(_w_14763));
  bfr _b_12859(.a(_w_14761),.q(_w_14762));
  bfr _b_12858(.a(_w_14760),.q(n1878));
  bfr _b_12857(.a(_w_14759),.q(_w_14760));
  bfr _b_12856(.a(_w_14758),.q(_w_14759));
  bfr _b_12855(.a(_w_14757),.q(_w_14758));
  bfr _b_12854(.a(_w_14756),.q(_w_14757));
  bfr _b_12853(.a(_w_14755),.q(_w_14756));
  bfr _b_12850(.a(_w_14752),.q(_w_14753));
  bfr _b_12849(.a(_w_14751),.q(_w_14752));
  bfr _b_12848(.a(_w_14750),.q(_w_14751));
  bfr _b_12845(.a(_w_14747),.q(_w_14748));
  bfr _b_12844(.a(_w_14746),.q(_w_14747));
  bfr _b_12843(.a(_w_14745),.q(_w_14746));
  bfr _b_12842(.a(_w_14744),.q(_w_14745));
  bfr _b_12840(.a(_w_14742),.q(_w_14743));
  bfr _b_12839(.a(_w_14741),.q(_w_14742));
  bfr _b_12836(.a(_w_14738),.q(_w_14739));
  bfr _b_12834(.a(_w_14736),.q(n1877));
  bfr _b_12831(.a(_w_14733),.q(_w_14734));
  bfr _b_12830(.a(_w_14732),.q(_w_14733));
  bfr _b_13549(.a(_w_15451),.q(_w_15452));
  bfr _b_12829(.a(_w_14731),.q(_w_14732));
  bfr _b_12827(.a(_w_14729),.q(_w_14730));
  bfr _b_12826(.a(_w_14728),.q(_w_14729));
  bfr _b_12825(.a(_w_14727),.q(_w_14728));
  bfr _b_12824(.a(_w_14726),.q(_w_14727));
  bfr _b_12823(.a(_w_14725),.q(_w_14726));
  bfr _b_12822(.a(_w_14724),.q(_w_14725));
  bfr _b_12821(.a(_w_14723),.q(_w_14724));
  bfr _b_13817(.a(_w_15719),.q(_w_15720));
  bfr _b_12817(.a(_w_14719),.q(_w_14720));
  bfr _b_12816(.a(_w_14718),.q(_w_14719));
  bfr _b_12814(.a(_w_14716),.q(_w_14717));
  bfr _b_12813(.a(_w_14715),.q(_w_14716));
  bfr _b_12812(.a(_w_14714),.q(_w_14715));
  bfr _b_12811(.a(_w_14713),.q(_w_14714));
  bfr _b_12808(.a(_w_14710),.q(_w_14711));
  bfr _b_12806(.a(_w_14708),.q(_w_14709));
  bfr _b_12804(.a(_w_14706),.q(_w_14707));
  bfr _b_12803(.a(_w_14705),.q(_w_14706));
  bfr _b_12802(.a(_w_14704),.q(_w_14705));
  bfr _b_12799(.a(_w_14701),.q(_w_14702));
  bfr _b_12837(.a(_w_14739),.q(_w_14740));
  bfr _b_12797(.a(_w_14699),.q(_w_14700));
  bfr _b_12792(.a(_w_14694),.q(_w_14695));
  bfr _b_12790(.a(_w_14692),.q(_w_14693));
  bfr _b_12789(.a(_w_14691),.q(_w_14692));
  bfr _b_12787(.a(_w_14689),.q(_w_14690));
  bfr _b_12785(.a(_w_14687),.q(n1868));
  bfr _b_12784(.a(_w_14686),.q(n1859));
  bfr _b_12782(.a(_w_14684),.q(_w_14685));
  bfr _b_12780(.a(_w_14682),.q(_w_14683));
  bfr _b_12779(.a(_w_14681),.q(_w_14682));
  bfr _b_12778(.a(_w_14680),.q(_w_14681));
  bfr _b_12776(.a(_w_14678),.q(_w_14679));
  bfr _b_12775(.a(_w_14677),.q(_w_14678));
  bfr _b_12774(.a(_w_14676),.q(_w_14677));
  bfr _b_12773(.a(_w_14675),.q(_w_14676));
  bfr _b_12771(.a(_w_14673),.q(n1855));
  bfr _b_12770(.a(_w_14672),.q(_w_14673));
  bfr _b_12769(.a(_w_14671),.q(_w_14672));
  bfr _b_12768(.a(_w_14670),.q(_w_14671));
  bfr _b_12767(.a(_w_14669),.q(_w_14670));
  bfr _b_12766(.a(_w_14668),.q(_w_14669));
  bfr _b_12762(.a(_w_14664),.q(_w_14665));
  bfr _b_12760(.a(_w_14662),.q(_w_14663));
  bfr _b_12759(.a(_w_14661),.q(_w_14662));
  bfr _b_12758(.a(_w_14660),.q(_w_14661));
  bfr _b_12754(.a(_w_14656),.q(_w_14657));
  bfr _b_12753(.a(_w_14655),.q(_w_14656));
  bfr _b_12752(.a(_w_14654),.q(_w_14655));
  bfr _b_12751(.a(_w_14653),.q(_w_14654));
  bfr _b_12748(.a(_w_14650),.q(_w_14651));
  bfr _b_12746(.a(_w_14648),.q(_w_14649));
  bfr _b_12745(.a(_w_14647),.q(_w_14648));
  bfr _b_12744(.a(_w_14646),.q(_w_14647));
  bfr _b_12743(.a(_w_14645),.q(_w_14646));
  bfr _b_12742(.a(_w_14644),.q(_w_14645));
  bfr _b_12741(.a(_w_14643),.q(_w_14644));
  bfr _b_12740(.a(_w_14642),.q(_w_14643));
  bfr _b_12738(.a(_w_14640),.q(_w_14641));
  bfr _b_12737(.a(_w_14639),.q(_w_14640));
  bfr _b_12735(.a(_w_14637),.q(_w_14638));
  bfr _b_12732(.a(_w_14634),.q(_w_14635));
  bfr _b_12729(.a(_w_14631),.q(_w_14632));
  bfr _b_12728(.a(_w_14630),.q(_w_14631));
  bfr _b_12725(.a(_w_14627),.q(_w_14628));
  bfr _b_12724(.a(_w_14626),.q(_w_14627));
  bfr _b_12723(.a(_w_14625),.q(_w_14626));
  bfr _b_12721(.a(_w_14623),.q(_w_14624));
  bfr _b_12720(.a(_w_14622),.q(_w_14623));
  bfr _b_12719(.a(_w_14621),.q(_w_14622));
  bfr _b_12718(.a(_w_14620),.q(_w_14621));
  bfr _b_12717(.a(_w_14619),.q(_w_14620));
  bfr _b_12713(.a(_w_14615),.q(_w_14616));
  bfr _b_12711(.a(_w_14613),.q(n1432));
  bfr _b_12710(.a(_w_14612),.q(n1845));
  bfr _b_12709(.a(_w_14611),.q(_w_14612));
  bfr _b_12708(.a(_w_14610),.q(_w_14611));
  bfr _b_12707(.a(_w_14609),.q(_w_14610));
  bfr _b_12699(.a(_w_14601),.q(_w_14602));
  bfr _b_12697(.a(_w_14599),.q(_w_14600));
  bfr _b_12695(.a(_w_14597),.q(_w_14598));
  bfr _b_12694(.a(_w_14596),.q(_w_14597));
  bfr _b_12693(.a(_w_14595),.q(_w_14596));
  bfr _b_12691(.a(_w_14593),.q(_w_14594));
  bfr _b_12689(.a(_w_14591),.q(_w_14592));
  bfr _b_12686(.a(_w_14588),.q(_w_14589));
  bfr _b_12685(.a(_w_14587),.q(_w_14588));
  bfr _b_12684(.a(_w_14586),.q(_w_14587));
  bfr _b_12938(.a(_w_14840),.q(_w_14841));
  bfr _b_12682(.a(_w_14584),.q(_w_14585));
  bfr _b_12680(.a(_w_14582),.q(_w_14583));
  bfr _b_12678(.a(_w_14580),.q(_w_14581));
  bfr _b_12677(.a(_w_14579),.q(_w_14580));
  bfr _b_12676(.a(_w_14578),.q(_w_14579));
  bfr _b_12675(.a(_w_14577),.q(_w_14578));
  bfr _b_12673(.a(_w_14575),.q(_w_14576));
  bfr _b_12670(.a(_w_14572),.q(n1837));
  bfr _b_12669(.a(_w_14571),.q(n1831));
  bfr _b_12666(.a(_w_14568),.q(n1825));
  bfr _b_12665(.a(_w_14567),.q(_w_14568));
  bfr _b_12993(.a(_w_14895),.q(_w_14896));
  bfr _b_12664(.a(_w_14566),.q(_w_14567));
  bfr _b_12663(.a(_w_14565),.q(_w_14566));
  bfr _b_12661(.a(_w_14563),.q(_w_14564));
  bfr _b_12660(.a(_w_14562),.q(_w_14563));
  bfr _b_12659(.a(_w_14561),.q(_w_14562));
  bfr _b_13420(.a(_w_15322),.q(_w_15323));
  bfr _b_12658(.a(_w_14560),.q(_w_14561));
  bfr _b_12656(.a(_w_14558),.q(_w_14559));
  bfr _b_12654(.a(_w_14556),.q(N6250));
  bfr _b_12653(.a(_w_14555),.q(_w_14556));
  bfr _b_12652(.a(_w_14554),.q(_w_14555));
  bfr _b_12647(.a(_w_14549),.q(_w_14550));
  bfr _b_12645(.a(_w_14547),.q(_w_14548));
  bfr _b_12643(.a(_w_14545),.q(_w_14546));
  bfr _b_12636(.a(_w_14538),.q(_w_14539));
  bfr _b_12634(.a(_w_14536),.q(_w_14537));
  bfr _b_12631(.a(_w_14533),.q(_w_14534));
  bfr _b_12629(.a(_w_14531),.q(_w_14532));
  bfr _b_12628(.a(_w_14530),.q(_w_14531));
  bfr _b_14383(.a(_w_16285),.q(_w_16286));
  bfr _b_12872(.a(_w_14774),.q(_w_14775));
  bfr _b_12626(.a(_w_14528),.q(_w_14529));
  bfr _b_12624(.a(_w_14526),.q(_w_14527));
  bfr _b_12621(.a(_w_14523),.q(n1801));
  bfr _b_12619(.a(_w_14521),.q(N2548));
  bfr _b_12618(.a(_w_14520),.q(_w_14521));
  bfr _b_13870(.a(_w_15772),.q(_w_15773));
  bfr _b_12617(.a(_w_14519),.q(_w_14520));
  bfr _b_13142(.a(_w_15044),.q(_w_15045));
  bfr _b_12615(.a(_w_14517),.q(_w_14518));
  bfr _b_12614(.a(_w_14516),.q(_w_14517));
  bfr _b_12610(.a(_w_14512),.q(_w_14513));
  bfr _b_12609(.a(_w_14511),.q(_w_14512));
  bfr _b_12608(.a(_w_14510),.q(_w_14511));
  bfr _b_12606(.a(_w_14508),.q(_w_14509));
  bfr _b_13141(.a(_w_15043),.q(n1839_1));
  bfr _b_12605(.a(_w_14507),.q(_w_14508));
  bfr _b_12604(.a(_w_14506),.q(_w_14507));
  bfr _b_12603(.a(_w_14505),.q(_w_14506));
  bfr _b_12601(.a(_w_14503),.q(_w_14504));
  bfr _b_12600(.a(_w_14502),.q(_w_14503));
  bfr _b_12596(.a(_w_14498),.q(_w_14499));
  bfr _b_12595(.a(_w_14497),.q(_w_14498));
  bfr _b_12594(.a(_w_14496),.q(_w_14497));
  bfr _b_12593(.a(_w_14495),.q(_w_14496));
  bfr _b_12592(.a(_w_14494),.q(_w_14495));
  bfr _b_12590(.a(_w_14492),.q(_w_14493));
  bfr _b_12589(.a(_w_14491),.q(_w_14492));
  bfr _b_12588(.a(_w_14490),.q(_w_14491));
  bfr _b_13125(.a(_w_15027),.q(_w_15028));
  bfr _b_12587(.a(_w_14489),.q(_w_14490));
  bfr _b_12584(.a(_w_14486),.q(_w_14487));
  bfr _b_12583(.a(_w_14485),.q(_w_14486));
  bfr _b_12582(.a(_w_14484),.q(_w_14485));
  bfr _b_12581(.a(_w_14483),.q(_w_14484));
  bfr _b_12579(.a(_w_14481),.q(_w_14482));
  bfr _b_12576(.a(_w_14478),.q(_w_14479));
  bfr _b_12575(.a(_w_14477),.q(_w_14478));
  bfr _b_12570(.a(_w_14472),.q(_w_14473));
  bfr _b_12569(.a(_w_14471),.q(_w_14472));
  bfr _b_12568(.a(_w_14470),.q(_w_14471));
  bfr _b_12567(.a(_w_14469),.q(_w_14470));
  bfr _b_12565(.a(_w_14467),.q(_w_14468));
  bfr _b_12563(.a(_w_14465),.q(_w_14466));
  bfr _b_12561(.a(_w_14463),.q(_w_14464));
  bfr _b_13698(.a(_w_15600),.q(_w_15601));
  bfr _b_12560(.a(_w_14462),.q(_w_14463));
  bfr _b_12559(.a(_w_14461),.q(_w_14462));
  bfr _b_12558(.a(_w_14460),.q(_w_14461));
  bfr _b_12630(.a(_w_14532),.q(_w_14533));
  bfr _b_12557(.a(_w_14459),.q(_w_14460));
  bfr _b_12554(.a(_w_14456),.q(_w_14457));
  bfr _b_12550(.a(_w_14452),.q(_w_14453));
  bfr _b_12546(.a(_w_14448),.q(_w_14449));
  bfr _b_12545(.a(_w_14447),.q(_w_14448));
  bfr _b_12544(.a(_w_14446),.q(_w_14447));
  bfr _b_12543(.a(_w_14445),.q(_w_14446));
  bfr _b_12539(.a(_w_14441),.q(_w_14442));
  bfr _b_12538(.a(_w_14440),.q(_w_14441));
  bfr _b_12537(.a(_w_14439),.q(_w_14440));
  bfr _b_12535(.a(_w_14437),.q(_w_14438));
  bfr _b_12534(.a(_w_14436),.q(_w_14437));
  bfr _b_12533(.a(_w_14435),.q(_w_14436));
  bfr _b_14070(.a(_w_15972),.q(_w_15973));
  bfr _b_12531(.a(_w_14433),.q(_w_14434));
  bfr _b_12528(.a(_w_14430),.q(_w_14431));
  bfr _b_13718(.a(_w_15620),.q(_w_15596));
  bfr _b_12525(.a(_w_14427),.q(_w_14428));
  bfr _b_12522(.a(_w_14424),.q(_w_14425));
  bfr _b_12521(.a(_w_14423),.q(_w_14424));
  bfr _b_12519(.a(_w_14421),.q(_w_14422));
  bfr _b_14347(.a(_w_16249),.q(_w_16250));
  bfr _b_12518(.a(_w_14420),.q(_w_14421));
  bfr _b_13169(.a(_w_15071),.q(n218));
  bfr _b_12517(.a(_w_14419),.q(_w_14420));
  bfr _b_12516(.a(_w_14418),.q(_w_14419));
  bfr _b_12515(.a(_w_14417),.q(_w_14418));
  bfr _b_14066(.a(_w_15968),.q(_w_15969));
  bfr _b_12513(.a(_w_14415),.q(_w_14416));
  bfr _b_12510(.a(_w_14412),.q(_w_14413));
  bfr _b_12509(.a(_w_14411),.q(_w_14412));
  bfr _b_12508(.a(_w_14410),.q(_w_14411));
  bfr _b_12507(.a(_w_14409),.q(_w_14410));
  bfr _b_12504(.a(_w_14406),.q(_w_14407));
  bfr _b_12503(.a(_w_14405),.q(_w_14406));
  bfr _b_12502(.a(_w_14404),.q(_w_14405));
  bfr _b_12501(.a(_w_14403),.q(_w_14404));
  bfr _b_12497(.a(_w_14399),.q(_w_14400));
  bfr _b_12492(.a(_w_14394),.q(_w_14395));
  bfr _b_13997(.a(_w_15899),.q(_w_15900));
  bfr _b_12491(.a(_w_14393),.q(_w_14394));
  bfr _b_13912(.a(_w_15814),.q(_w_15815));
  bfr _b_12488(.a(_w_14390),.q(_w_14391));
  bfr _b_12487(.a(_w_14389),.q(_w_14390));
  bfr _b_12486(.a(_w_14388),.q(_w_14389));
  bfr _b_12485(.a(_w_14387),.q(_w_14388));
  bfr _b_12483(.a(_w_14385),.q(_w_14386));
  bfr _b_12481(.a(_w_14383),.q(_w_14384));
  bfr _b_12480(.a(_w_14382),.q(_w_14383));
  bfr _b_12476(.a(_w_14378),.q(_w_14379));
  bfr _b_12472(.a(_w_14374),.q(_w_14375));
  bfr _b_12471(.a(_w_14373),.q(N69_7));
  bfr _b_12702(.a(_w_14604),.q(_w_14605));
  bfr _b_12469(.a(_w_14371),.q(N69_6));
  bfr _b_12467(.a(_w_14369),.q(n1792));
  bfr _b_12465(.a(_w_14367),.q(_w_14368));
  bfr _b_12464(.a(_w_14366),.q(_w_14367));
  bfr _b_12461(.a(_w_14363),.q(_w_14364));
  bfr _b_12456(.a(_w_14358),.q(_w_14359));
  bfr _b_12455(.a(_w_14357),.q(_w_14358));
  bfr _b_12454(.a(_w_14356),.q(_w_14357));
  bfr _b_12450(.a(_w_14352),.q(_w_14353));
  bfr _b_12446(.a(_w_14348),.q(n1783));
  bfr _b_12444(.a(_w_14346),.q(_w_14347));
  bfr _b_12443(.a(_w_14345),.q(_w_14346));
  bfr _b_14105(.a(_w_16007),.q(_w_16008));
  bfr _b_12442(.a(_w_14344),.q(_w_14345));
  bfr _b_12441(.a(_w_14343),.q(_w_14344));
  bfr _b_12440(.a(_w_14342),.q(_w_14343));
  bfr _b_12439(.a(_w_14341),.q(_w_14342));
  bfr _b_14228(.a(_w_16130),.q(_w_16131));
  bfr _b_12437(.a(_w_14339),.q(n1770));
  bfr _b_12436(.a(_w_14338),.q(_w_14339));
  bfr _b_12434(.a(_w_14336),.q(_w_14337));
  bfr _b_12429(.a(_w_14331),.q(_w_14332));
  bfr _b_12428(.a(_w_14330),.q(_w_14331));
  bfr _b_12427(.a(_w_14329),.q(_w_14330));
  bfr _b_12426(.a(_w_14328),.q(_w_14329));
  bfr _b_13937(.a(_w_15839),.q(_w_15840));
  bfr _b_12425(.a(_w_14327),.q(_w_14328));
  bfr _b_12422(.a(_w_14324),.q(_w_14325));
  bfr _b_12421(.a(_w_14323),.q(_w_14324));
  bfr _b_12420(.a(_w_14322),.q(_w_14323));
  bfr _b_12419(.a(_w_14321),.q(_w_14322));
  bfr _b_12418(.a(_w_14320),.q(_w_14321));
  bfr _b_14014(.a(_w_15916),.q(_w_15917));
  bfr _b_12409(.a(_w_14311),.q(_w_14312));
  bfr _b_12408(.a(_w_14310),.q(_w_14311));
  bfr _b_12407(.a(_w_14309),.q(_w_14310));
  bfr _b_12404(.a(_w_14306),.q(n1763));
  bfr _b_12403(.a(_w_14305),.q(n308_2));
  bfr _b_12402(.a(_w_14304),.q(_w_14305));
  bfr _b_12401(.a(_w_14303),.q(n308_1));
  bfr _b_12400(.a(_w_14302),.q(_w_14303));
  bfr _b_12399(.a(_w_14301),.q(n1101_1));
  bfr _b_12397(.a(_w_14299),.q(_w_14300));
  bfr _b_14127(.a(_w_16029),.q(_w_16030));
  bfr _b_12396(.a(_w_14298),.q(_w_14299));
  bfr _b_12395(.a(_w_14297),.q(n736));
  bfr _b_12392(.a(_w_14294),.q(_w_14295));
  bfr _b_12391(.a(_w_14293),.q(_w_14294));
  bfr _b_12390(.a(_w_14292),.q(_w_14293));
  bfr _b_13305(.a(_w_15207),.q(_w_15208));
  bfr _b_12791(.a(_w_14693),.q(_w_14694));
  bfr _b_12389(.a(_w_14291),.q(n1757));
  bfr _b_12649(.a(_w_14551),.q(_w_14552));
  bfr _b_12388(.a(_w_14290),.q(n200));
  bfr _b_12387(.a(_w_14289),.q(n1754));
  bfr _b_12385(.a(_w_14287),.q(_w_14288));
  bfr _b_12383(.a(_w_14285),.q(_w_14286));
  bfr _b_12382(.a(_w_14284),.q(_w_14285));
  bfr _b_12381(.a(_w_14283),.q(_w_14284));
  bfr _b_12380(.a(_w_14282),.q(_w_14283));
  bfr _b_12377(.a(_w_14279),.q(_w_14280));
  bfr _b_12376(.a(_w_14278),.q(_w_14279));
  bfr _b_12373(.a(_w_14275),.q(n1846));
  bfr _b_12372(.a(_w_14274),.q(_w_14275));
  bfr _b_12371(.a(_w_14273),.q(_w_14274));
  bfr _b_12368(.a(_w_14270),.q(_w_14271));
  bfr _b_12367(.a(_w_14269),.q(_w_14270));
  bfr _b_12365(.a(_w_14267),.q(_w_14268));
  bfr _b_12363(.a(_w_14265),.q(_w_14266));
  bfr _b_12362(.a(_w_14264),.q(_w_14265));
  bfr _b_12361(.a(_w_14263),.q(_w_14264));
  bfr _b_12358(.a(_w_14260),.q(_w_14261));
  bfr _b_12357(.a(_w_14259),.q(_w_14260));
  bfr _b_12355(.a(_w_14257),.q(_w_14258));
  bfr _b_12354(.a(_w_14256),.q(_w_14257));
  bfr _b_12352(.a(_w_14254),.q(_w_14255));
  bfr _b_12351(.a(_w_14253),.q(_w_14254));
  bfr _b_13778(.a(_w_15680),.q(_w_15681));
  bfr _b_12347(.a(_w_14249),.q(_w_14250));
  bfr _b_12345(.a(_w_14247),.q(_w_14248));
  bfr _b_12344(.a(_w_14246),.q(_w_14247));
  bfr _b_12342(.a(_w_14244),.q(_w_14245));
  bfr _b_13795(.a(_w_15697),.q(_w_15698));
  bfr _b_12341(.a(_w_14243),.q(_w_14244));
  bfr _b_12340(.a(_w_14242),.q(_w_14243));
  bfr _b_12338(.a(_w_14240),.q(_w_14241));
  bfr _b_12337(.a(_w_14239),.q(_w_14240));
  bfr _b_12335(.a(_w_14237),.q(_w_14238));
  bfr _b_12334(.a(_w_14236),.q(_w_14237));
  bfr _b_12333(.a(_w_14235),.q(_w_14236));
  bfr _b_12326(.a(_w_14228),.q(_w_14229));
  bfr _b_12324(.a(_w_14226),.q(_w_14227));
  bfr _b_12323(.a(_w_14225),.q(n1734));
  bfr _b_12322(.a(_w_14224),.q(_w_14225));
  bfr _b_12321(.a(_w_14223),.q(_w_14224));
  bfr _b_12318(.a(_w_14220),.q(_w_14221));
  bfr _b_12316(.a(_w_14218),.q(_w_14219));
  bfr _b_12315(.a(_w_14217),.q(n568));
  bfr _b_12314(.a(_w_14216),.q(n1732));
  bfr _b_12312(.a(_w_14214),.q(_w_14215));
  bfr _b_12311(.a(_w_14213),.q(_w_14214));
  bfr _b_12310(.a(_w_14212),.q(_w_14213));
  bfr _b_12309(.a(_w_14211),.q(_w_14212));
  bfr _b_12308(.a(_w_14210),.q(_w_14211));
  bfr _b_12303(.a(_w_14205),.q(_w_14206));
  bfr _b_12302(.a(_w_14204),.q(_w_14205));
  bfr _b_12301(.a(_w_14203),.q(_w_14204));
  bfr _b_12300(.a(_w_14202),.q(_w_14203));
  bfr _b_12299(.a(_w_14201),.q(_w_14202));
  bfr _b_12298(.a(_w_14200),.q(n1730));
  bfr _b_12297(.a(_w_14199),.q(_w_14200));
  bfr _b_12295(.a(_w_14197),.q(_w_14198));
  bfr _b_14016(.a(_w_15918),.q(_w_15919));
  bfr _b_12294(.a(_w_14196),.q(_w_14197));
  bfr _b_12293(.a(_w_14195),.q(_w_14196));
  bfr _b_12292(.a(_w_14194),.q(_w_14195));
  bfr _b_12291(.a(_w_14193),.q(_w_14194));
  bfr _b_12287(.a(_w_14189),.q(_w_14190));
  bfr _b_13198(.a(_w_15100),.q(n1521_1));
  bfr _b_12285(.a(_w_14187),.q(_w_14188));
  bfr _b_12284(.a(_w_14186),.q(_w_14187));
  bfr _b_12283(.a(_w_14185),.q(_w_14186));
  bfr _b_12279(.a(_w_14181),.q(_w_14182));
  bfr _b_12278(.a(_w_14180),.q(_w_14181));
  bfr _b_12273(.a(_w_14175),.q(_w_14176));
  bfr _b_12270(.a(_w_14172),.q(_w_14173));
  bfr _b_12268(.a(_w_14170),.q(_w_14171));
  bfr _b_12267(.a(_w_14169),.q(_w_14170));
  bfr _b_12266(.a(_w_14168),.q(_w_14169));
  bfr _b_13158(.a(_w_15060),.q(_w_15061));
  bfr _b_12264(.a(_w_14166),.q(_w_14167));
  bfr _b_12263(.a(_w_14165),.q(_w_14166));
  bfr _b_12259(.a(_w_14161),.q(_w_14162));
  bfr _b_12257(.a(_w_14159),.q(_w_14160));
  bfr _b_12255(.a(_w_14157),.q(_w_14158));
  bfr _b_12254(.a(_w_14156),.q(_w_14157));
  bfr _b_12253(.a(_w_14155),.q(_w_14156));
  bfr _b_12252(.a(_w_14154),.q(_w_14155));
  bfr _b_12248(.a(_w_14150),.q(n1721));
  bfr _b_12246(.a(_w_14148),.q(_w_14149));
  bfr _b_12245(.a(_w_14147),.q(_w_14148));
  bfr _b_12242(.a(_w_14144),.q(_w_14145));
  bfr _b_12240(.a(_w_14142),.q(_w_14143));
  bfr _b_12239(.a(_w_14141),.q(_w_14142));
  bfr _b_12238(.a(_w_14140),.q(_w_14141));
  bfr _b_12235(.a(_w_14137),.q(_w_14138));
  bfr _b_12234(.a(_w_14136),.q(_w_14137));
  bfr _b_12233(.a(_w_14135),.q(_w_14136));
  bfr _b_12232(.a(_w_14134),.q(_w_14135));
  bfr _b_12231(.a(_w_14133),.q(_w_14134));
  bfr _b_12228(.a(_w_14130),.q(_w_14131));
  bfr _b_12227(.a(_w_14129),.q(_w_14130));
  bfr _b_12225(.a(_w_14127),.q(_w_14128));
  bfr _b_12222(.a(_w_14124),.q(_w_14125));
  bfr _b_12221(.a(_w_14123),.q(_w_14124));
  bfr _b_12218(.a(_w_14120),.q(_w_14121));
  bfr _b_12217(.a(_w_14119),.q(_w_14120));
  bfr _b_12215(.a(_w_14117),.q(n1705));
  bfr _b_12213(.a(_w_14115),.q(n1696));
  bfr _b_12212(.a(_w_14114),.q(n1693));
  bfr _b_12209(.a(_w_14111),.q(_w_14112));
  bfr _b_12208(.a(_w_14110),.q(_w_14111));
  bfr _b_12207(.a(_w_14109),.q(_w_14110));
  bfr _b_12206(.a(_w_14108),.q(n966));
  bfr _b_12204(.a(_w_14106),.q(n1879));
  bfr _b_12700(.a(_w_14602),.q(_w_14603));
  bfr _b_12203(.a(_w_14105),.q(_w_14106));
  bfr _b_12201(.a(_w_14103),.q(_w_14104));
  bfr _b_12200(.a(_w_14102),.q(_w_14103));
  bfr _b_12198(.a(_w_14100),.q(_w_14101));
  bfr _b_12194(.a(_w_14096),.q(_w_14097));
  bfr _b_12190(.a(_w_14092),.q(_w_14093));
  bfr _b_12189(.a(_w_14091),.q(_w_14092));
  bfr _b_12188(.a(_w_14090),.q(_w_14091));
  bfr _b_12186(.a(_w_14088),.q(_w_14089));
  bfr _b_12184(.a(_w_14086),.q(n1677));
  bfr _b_12182(.a(_w_14084),.q(_w_14085));
  bfr _b_12181(.a(_w_14083),.q(_w_14084));
  bfr _b_12180(.a(_w_14082),.q(_w_14083));
  bfr _b_12174(.a(_w_14076),.q(_w_14077));
  bfr _b_12170(.a(_w_14072),.q(_w_14073));
  bfr _b_13490(.a(_w_15392),.q(_w_15393));
  bfr _b_12168(.a(_w_14070),.q(_w_14071));
  bfr _b_12167(.a(_w_14069),.q(_w_14070));
  bfr _b_12165(.a(_w_14067),.q(_w_14068));
  bfr _b_12164(.a(_w_14066),.q(_w_14067));
  bfr _b_12163(.a(_w_14065),.q(_w_14066));
  bfr _b_12162(.a(_w_14064),.q(_w_14065));
  bfr _b_12161(.a(_w_14063),.q(_w_14064));
  bfr _b_13126(.a(_w_15028),.q(_w_15029));
  bfr _b_12159(.a(_w_14061),.q(_w_14062));
  bfr _b_12158(.a(_w_14060),.q(_w_14061));
  bfr _b_12155(.a(_w_14057),.q(n1675));
  bfr _b_12150(.a(_w_14052),.q(_w_14053));
  bfr _b_12149(.a(_w_14051),.q(_w_14052));
  bfr _b_12147(.a(_w_14049),.q(_w_14050));
  bfr _b_12142(.a(_w_14044),.q(_w_14045));
  bfr _b_12139(.a(_w_14041),.q(n754_1));
  bfr _b_12138(.a(_w_14040),.q(_w_14041));
  bfr _b_12136(.a(_w_14038),.q(_w_14039));
  bfr _b_12134(.a(_w_14036),.q(_w_14037));
  bfr _b_12133(.a(_w_14035),.q(_w_14036));
  bfr _b_12130(.a(_w_14032),.q(_w_14033));
  bfr _b_12121(.a(_w_14023),.q(_w_14024));
  bfr _b_12119(.a(_w_14021),.q(_w_14022));
  bfr _b_12118(.a(_w_14020),.q(_w_14021));
  bfr _b_12113(.a(_w_14015),.q(_w_14016));
  bfr _b_12112(.a(_w_14014),.q(_w_14015));
  bfr _b_12105(.a(_w_14007),.q(_w_14008));
  bfr _b_12103(.a(_w_14005),.q(_w_14006));
  bfr _b_12101(.a(_w_14003),.q(_w_14004));
  bfr _b_12100(.a(_w_14002),.q(_w_14003));
  bfr _b_12098(.a(_w_14000),.q(_w_14001));
  bfr _b_12097(.a(_w_13999),.q(_w_14000));
  bfr _b_12095(.a(_w_13997),.q(_w_13998));
  bfr _b_14259(.a(_w_16161),.q(_w_16162));
  bfr _b_14009(.a(_w_15911),.q(_w_15912));
  bfr _b_12756(.a(_w_14658),.q(_w_14659));
  bfr _b_12094(.a(_w_13996),.q(_w_13997));
  bfr _b_12092(.a(_w_13994),.q(_w_13995));
  bfr _b_12091(.a(_w_13993),.q(_w_13994));
  bfr _b_12089(.a(_w_13991),.q(_w_13992));
  bfr _b_12086(.a(_w_13988),.q(_w_13989));
  bfr _b_12085(.a(_w_13987),.q(_w_13988));
  bfr _b_12083(.a(_w_13985),.q(n1663));
  bfr _b_12081(.a(_w_13983),.q(n790_1));
  bfr _b_12080(.a(_w_13982),.q(_w_13983));
  bfr _b_12079(.a(_w_13981),.q(_w_13982));
  bfr _b_12070(.a(_w_13972),.q(_w_13973));
  bfr _b_12069(.a(_w_13971),.q(_w_13972));
  bfr _b_12066(.a(_w_13968),.q(_w_13969));
  bfr _b_12065(.a(_w_13967),.q(_w_13968));
  bfr _b_12064(.a(_w_13966),.q(_w_13967));
  bfr _b_12063(.a(_w_13965),.q(n1612));
  bfr _b_12060(.a(_w_13962),.q(_w_13963));
  bfr _b_12058(.a(_w_13960),.q(_w_13961));
  bfr _b_12057(.a(_w_13959),.q(_w_13960));
  bfr _b_12056(.a(_w_13958),.q(_w_13959));
  bfr _b_12055(.a(_w_13957),.q(n1598));
  bfr _b_12053(.a(_w_13955),.q(n430_1));
  bfr _b_12052(.a(_w_13954),.q(_w_13955));
  bfr _b_12050(.a(_w_13952),.q(_w_13953));
  bfr _b_12044(.a(_w_13946),.q(_w_13947));
  bfr _b_12043(.a(_w_13945),.q(_w_13946));
  bfr _b_12042(.a(_w_13944),.q(_w_13945));
  bfr _b_12039(.a(_w_13941),.q(n1574));
  bfr _b_12038(.a(_w_13940),.q(n1816));
  bfr _b_12036(.a(_w_13938),.q(n1565));
  bfr _b_12035(.a(_w_13937),.q(n1479_1));
  bfr _b_12033(.a(_w_13935),.q(_w_13936));
  bfr _b_12031(.a(_w_13933),.q(n1562));
  bfr _b_12030(.a(_w_13932),.q(n1556));
  bfr _b_12029(.a(_w_13931),.q(n1704_1));
  bfr _b_12027(.a(_w_13929),.q(_w_13930));
  bfr _b_12025(.a(_w_13927),.q(n1553));
  bfr _b_12024(.a(_w_13926),.q(n1545));
  bfr _b_12022(.a(_w_13924),.q(_w_13925));
  bfr _b_12016(.a(_w_13918),.q(_w_13919));
  bfr _b_12014(.a(_w_13916),.q(_w_13917));
  bfr _b_12011(.a(_w_13913),.q(_w_13914));
  bfr _b_12009(.a(_w_13911),.q(_w_13912));
  bfr _b_12008(.a(_w_13910),.q(_w_13911));
  bfr _b_12005(.a(_w_13907),.q(_w_13908));
  bfr _b_12004(.a(_w_13906),.q(n1014));
  bfr _b_12003(.a(_w_13905),.q(n1629_1));
  bfr _b_12002(.a(_w_13904),.q(_w_13905));
  bfr _b_12001(.a(_w_13903),.q(_w_13904));
  bfr _b_11999(.a(_w_13901),.q(n398));
  bfr _b_11997(.a(_w_13899),.q(_w_13900));
  bfr _b_11996(.a(_w_13898),.q(_w_13899));
  bfr _b_11994(.a(_w_13896),.q(_w_13897));
  bfr _b_11992(.a(_w_13894),.q(_w_13895));
  bfr _b_11991(.a(_w_13893),.q(_w_13894));
  bfr _b_11987(.a(_w_13889),.q(_w_13890));
  bfr _b_11986(.a(_w_13888),.q(_w_13889));
  bfr _b_11984(.a(_w_13886),.q(n1528));
  bfr _b_13101(.a(_w_15003),.q(_w_15004));
  bfr _b_11980(.a(_w_13882),.q(_w_13883));
  bfr _b_11979(.a(_w_13881),.q(_w_13882));
  bfr _b_11978(.a(_w_13880),.q(_w_13881));
  bfr _b_11977(.a(_w_13879),.q(_w_13880));
  bfr _b_11976(.a(_w_13878),.q(_w_13879));
  bfr _b_11975(.a(_w_13877),.q(_w_13878));
  bfr _b_11973(.a(_w_13875),.q(_w_13876));
  bfr _b_11971(.a(_w_13873),.q(n1522));
  bfr _b_11970(.a(_w_13872),.q(n570_1));
  bfr _b_12099(.a(_w_14001),.q(_w_14002));
  bfr _b_11969(.a(_w_13871),.q(_w_13872));
  bfr _b_11968(.a(_w_13870),.q(_w_13871));
  bfr _b_11965(.a(_w_13867),.q(n1095_1));
  bfr _b_11964(.a(_w_13866),.q(_w_13867));
  bfr _b_11962(.a(_w_13864),.q(_w_13865));
  bfr _b_11961(.a(_w_13863),.q(n1507));
  bfr _b_14190(.a(_w_16092),.q(_w_16093));
  bfr _b_11959(.a(_w_13861),.q(n460_1));
  bfr _b_11958(.a(_w_13860),.q(_w_13861));
  bfr _b_11956(.a(_w_13858),.q(_w_13859));
  bfr _b_11954(.a(_w_13856),.q(n1486));
  bfr _b_11953(.a(_w_13855),.q(n1480));
  bfr _b_11951(.a(_w_13853),.q(n46_1));
  bfr _b_11950(.a(_w_13852),.q(_w_13853));
  bfr _b_11949(.a(_w_13851),.q(_w_13852));
  bfr _b_13816(.a(_w_15718),.q(_w_15719));
  bfr _b_11948(.a(_w_13850),.q(_w_13851));
  bfr _b_11947(.a(_w_13849),.q(n1781));
  bfr _b_11945(.a(_w_13847),.q(_w_13848));
  bfr _b_11942(.a(_w_13844),.q(_w_13845));
  bfr _b_11940(.a(_w_13842),.q(_w_13843));
  bfr _b_11936(.a(_w_13838),.q(_w_13839));
  bfr _b_11935(.a(_w_13837),.q(_w_13838));
  bfr _b_11934(.a(_w_13836),.q(_w_13837));
  bfr _b_11933(.a(_w_13835),.q(_w_13836));
  bfr _b_11932(.a(_w_13834),.q(_w_13835));
  bfr _b_13294(.a(_w_15196),.q(_w_15197));
  bfr _b_11931(.a(_w_13833),.q(n1458));
  bfr _b_11930(.a(_w_13832),.q(_w_13833));
  bfr _b_11928(.a(_w_13830),.q(_w_13831));
  bfr _b_11927(.a(_w_13829),.q(_w_13830));
  bfr _b_11925(.a(_w_13827),.q(_w_13828));
  bfr _b_11924(.a(_w_13826),.q(_w_13827));
  bfr _b_11923(.a(_w_13825),.q(n1454));
  bfr _b_11922(.a(_w_13824),.q(_w_13825));
  bfr _b_11921(.a(_w_13823),.q(_w_13824));
  bfr _b_11918(.a(_w_13820),.q(_w_13821));
  bfr _b_11915(.a(_w_13817),.q(_w_13818));
  bfr _b_11914(.a(_w_13816),.q(_w_13817));
  bfr _b_11913(.a(_w_13815),.q(_w_13816));
  bfr _b_11912(.a(_w_13814),.q(_w_13815));
  bfr _b_12763(.a(_w_14665),.q(_w_14666));
  bfr _b_11910(.a(_w_13812),.q(_w_13813));
  bfr _b_11909(.a(_w_13811),.q(_w_13812));
  bfr _b_11908(.a(_w_13810),.q(_w_13811));
  bfr _b_11904(.a(_w_13806),.q(_w_13807));
  bfr _b_11903(.a(_w_13805),.q(_w_13806));
  bfr _b_11901(.a(_w_13803),.q(_w_13804));
  bfr _b_11897(.a(_w_13799),.q(_w_13800));
  bfr _b_11896(.a(_w_13798),.q(_w_13799));
  bfr _b_11895(.a(_w_13797),.q(_w_13798));
  bfr _b_11892(.a(_w_13794),.q(_w_13795));
  bfr _b_11891(.a(_w_13793),.q(_w_13794));
  bfr _b_12304(.a(_w_14206),.q(_w_14207));
  bfr _b_11889(.a(_w_13791),.q(_w_13792));
  bfr _b_11887(.a(_w_13789),.q(N103_14));
  bfr _b_11885(.a(_w_13787),.q(_w_13788));
  bfr _b_11884(.a(_w_13786),.q(_w_13787));
  bfr _b_11883(.a(_w_13785),.q(_w_13786));
  bfr _b_11880(.a(_w_13782),.q(_w_13783));
  bfr _b_11878(.a(_w_13780),.q(_w_13781));
  bfr _b_11876(.a(_w_13778),.q(_w_13779));
  bfr _b_11875(.a(_w_13777),.q(N103_13));
  bfr _b_11872(.a(_w_13774),.q(_w_13775));
  bfr _b_11870(.a(_w_13772),.q(_w_13773));
  bfr _b_11869(.a(_w_13771),.q(_w_13772));
  bfr _b_11868(.a(_w_13770),.q(_w_13771));
  bfr _b_14382(.a(_w_16284),.q(_w_16285));
  bfr _b_11865(.a(_w_13767),.q(_w_13768));
  bfr _b_13364(.a(_w_15266),.q(_w_15267));
  bfr _b_11863(.a(_w_13765),.q(_w_13766));
  bfr _b_13425(.a(_w_15327),.q(_w_15328));
  bfr _b_11862(.a(_w_13764),.q(_w_13765));
  bfr _b_11860(.a(_w_13762),.q(_w_13763));
  bfr _b_11858(.a(_w_13760),.q(_w_13761));
  bfr _b_11856(.a(_w_13758),.q(_w_13759));
  bfr _b_11853(.a(_w_13755),.q(n418_1));
  bfr _b_11850(.a(_w_13752),.q(_w_13753));
  bfr _b_11848(.a(_w_13750),.q(n1435));
  bfr _b_11846(.a(_w_13748),.q(_w_13749));
  bfr _b_11845(.a(_w_13747),.q(_w_13748));
  bfr _b_11844(.a(_w_13746),.q(_w_13747));
  bfr _b_11842(.a(_w_13744),.q(_w_13745));
  bfr _b_11837(.a(_w_13739),.q(_w_13740));
  bfr _b_11833(.a(_w_13735),.q(_w_13736));
  bfr _b_11832(.a(_w_13734),.q(_w_13735));
  bfr _b_11829(.a(_w_13731),.q(_w_13732));
  bfr _b_11828(.a(_w_13730),.q(_w_13731));
  bfr _b_11827(.a(_w_13729),.q(_w_13730));
  bfr _b_11825(.a(_w_13727),.q(_w_13728));
  bfr _b_11820(.a(_w_13722),.q(_w_13723));
  bfr _b_11867(.a(_w_13769),.q(n1450));
  bfr _b_11818(.a(_w_13720),.q(_w_13721));
  bfr _b_11817(.a(_w_13719),.q(_w_13720));
  bfr _b_11816(.a(_w_13718),.q(_w_13719));
  bfr _b_11812(.a(_w_13714),.q(_w_13715));
  bfr _b_11810(.a(_w_13712),.q(_w_13713));
  bfr _b_11805(.a(_w_13707),.q(_w_13708));
  bfr _b_11799(.a(_w_13701),.q(_w_13702));
  bfr _b_13423(.a(_w_15325),.q(_w_15326));
  bfr _b_11798(.a(_w_13700),.q(_w_13701));
  bfr _b_11795(.a(_w_13697),.q(_w_13698));
  bfr _b_11794(.a(_w_13696),.q(_w_13697));
  bfr _b_11791(.a(_w_13693),.q(_w_13694));
  bfr _b_11790(.a(_w_13692),.q(_w_13693));
  bfr _b_11789(.a(_w_13691),.q(_w_13692));
  bfr _b_11788(.a(_w_13690),.q(_w_13691));
  bfr _b_14083(.a(_w_15985),.q(_w_15986));
  bfr _b_11787(.a(_w_13689),.q(_w_13690));
  bfr _b_12282(.a(_w_14184),.q(_w_14185));
  bfr _b_11786(.a(_w_13688),.q(_w_13689));
  bfr _b_11785(.a(_w_13687),.q(_w_13688));
  bfr _b_11784(.a(_w_13686),.q(_w_13687));
  bfr _b_11783(.a(_w_13685),.q(_w_13686));
  bfr _b_14218(.a(_w_16120),.q(_w_16121));
  bfr _b_11782(.a(_w_13684),.q(_w_13685));
  bfr _b_11779(.a(_w_13681),.q(_w_13682));
  bfr _b_11778(.a(_w_13680),.q(_w_13681));
  bfr _b_12679(.a(_w_14581),.q(_w_14582));
  bfr _b_11776(.a(_w_13678),.q(_w_13679));
  bfr _b_11773(.a(_w_13675),.q(_w_13676));
  bfr _b_11772(.a(_w_13674),.q(_w_13675));
  bfr _b_11770(.a(_w_13672),.q(_w_13673));
  bfr _b_11767(.a(_w_13669),.q(_w_13670));
  bfr _b_11766(.a(_w_13668),.q(_w_13669));
  bfr _b_11764(.a(_w_13666),.q(_w_13667));
  bfr _b_11757(.a(_w_13659),.q(N1_2));
  bfr _b_11756(.a(_w_13658),.q(_w_13659));
  bfr _b_11755(.a(_w_13657),.q(_w_13658));
  bfr _b_11754(.a(_w_13656),.q(_w_13657));
  bfr _b_13482(.a(_w_15384),.q(_w_15385));
  bfr _b_11752(.a(_w_13654),.q(_w_13655));
  bfr _b_11750(.a(_w_13652),.q(_w_13653));
  bfr _b_11749(.a(_w_13651),.q(_w_13652));
  bfr _b_11748(.a(_w_13650),.q(_w_13651));
  bfr _b_11739(.a(_w_13641),.q(_w_13642));
  bfr _b_11738(.a(_w_13640),.q(_w_13641));
  bfr _b_12339(.a(_w_14241),.q(_w_14242));
  bfr _b_11735(.a(_w_13637),.q(_w_13638));
  bfr _b_12847(.a(_w_14749),.q(_w_14750));
  bfr _b_11734(.a(_w_13636),.q(_w_13637));
  bfr _b_11733(.a(_w_13635),.q(_w_13636));
  bfr _b_12453(.a(_w_14355),.q(_w_14356));
  bfr _b_11732(.a(_w_13634),.q(_w_13635));
  bfr _b_11731(.a(_w_13633),.q(_w_13634));
  bfr _b_11730(.a(_w_13632),.q(_w_13633));
  bfr _b_11729(.a(_w_13631),.q(_w_13632));
  bfr _b_12261(.a(_w_14163),.q(_w_14164));
  bfr _b_11726(.a(_w_13628),.q(_w_13629));
  bfr _b_11725(.a(_w_13627),.q(_w_13628));
  bfr _b_11724(.a(_w_13626),.q(_w_13627));
  bfr _b_11723(.a(_w_13625),.q(_w_13626));
  bfr _b_13150(.a(_w_15052),.q(n1748));
  bfr _b_11722(.a(_w_13624),.q(_w_13625));
  bfr _b_11720(.a(_w_13622),.q(_w_13623));
  bfr _b_12607(.a(_w_14509),.q(_w_14510));
  bfr _b_11718(.a(_w_13620),.q(_w_13621));
  bfr _b_11716(.a(_w_13618),.q(_w_13619));
  bfr _b_11715(.a(_w_13617),.q(_w_13618));
  bfr _b_11712(.a(_w_13614),.q(_w_13615));
  bfr _b_11711(.a(_w_13613),.q(_w_13614));
  bfr _b_12706(.a(_w_14608),.q(_w_14609));
  bfr _b_11710(.a(_w_13612),.q(_w_13613));
  bfr _b_11708(.a(_w_13610),.q(_w_13611));
  bfr _b_11707(.a(_w_13609),.q(_w_13610));
  bfr _b_11706(.a(_w_13608),.q(_w_13609));
  bfr _b_11705(.a(_w_13607),.q(_w_13608));
  bfr _b_11704(.a(_w_13606),.q(_w_13607));
  bfr _b_11703(.a(_w_13605),.q(N1_1));
  bfr _b_11702(.a(_w_13604),.q(_w_13605));
  bfr _b_11698(.a(_w_13600),.q(_w_13601));
  bfr _b_11695(.a(_w_13597),.q(_w_13598));
  bfr _b_11694(.a(_w_13596),.q(_w_13597));
  bfr _b_11692(.a(_w_13594),.q(_w_13595));
  bfr _b_11690(.a(_w_13592),.q(_w_13593));
  bfr _b_11686(.a(_w_13588),.q(_w_13589));
  bfr _b_11685(.a(_w_13587),.q(_w_13588));
  bfr _b_11684(.a(_w_13586),.q(_w_13587));
  bfr _b_11683(.a(_w_13585),.q(_w_13586));
  bfr _b_11681(.a(_w_13583),.q(n1426));
  bfr _b_11680(.a(_w_13582),.q(n1639));
  bfr _b_11679(.a(_w_13581),.q(n1420));
  bfr _b_11678(.a(_w_13580),.q(n1417));
  bfr _b_11675(.a(_w_13577),.q(n1402));
  bfr _b_11674(.a(_w_13576),.q(n40));
  bfr _b_13345(.a(_w_15247),.q(_w_15248));
  bfr _b_11673(.a(_w_13575),.q(_w_13576));
  bfr _b_11671(.a(_w_13573),.q(_w_13574));
  bfr _b_11668(.a(_w_13570),.q(n1393));
  bfr _b_11667(.a(_w_13569),.q(n1200_1));
  bfr _b_11665(.a(_w_13567),.q(_w_13568));
  bfr _b_11662(.a(_w_13564),.q(_w_13565));
  bfr _b_11659(.a(_w_13561),.q(n1390));
  bfr _b_11658(.a(_w_13560),.q(n1387));
  bfr _b_12571(.a(_w_14473),.q(_w_14474));
  bfr _b_11657(.a(_w_13559),.q(n1383));
  bfr _b_13058(.a(_w_14960),.q(_w_14961));
  bfr _b_11655(.a(_w_13557),.q(_w_13558));
  bfr _b_11654(.a(_w_13556),.q(_w_13557));
  bfr _b_11651(.a(_w_13553),.q(_w_13554));
  bfr _b_11649(.a(_w_13551),.q(_w_13552));
  bfr _b_11648(.a(_w_13550),.q(_w_13551));
  bfr _b_11647(.a(_w_13549),.q(_w_13550));
  bfr _b_11646(.a(_w_13548),.q(_w_13549));
  bfr _b_11645(.a(_w_13547),.q(_w_13548));
  bfr _b_11640(.a(_w_13542),.q(_w_13543));
  bfr _b_11638(.a(_w_13540),.q(_w_13541));
  bfr _b_13576(.a(_w_15478),.q(_w_15479));
  bfr _b_11637(.a(_w_13539),.q(n737_1));
  bfr _b_11634(.a(_w_13536),.q(n1373));
  bfr _b_11632(.a(_w_13534),.q(_w_13535));
  bfr _b_11629(.a(_w_13531),.q(_w_13532));
  bfr _b_11627(.a(_w_13529),.q(_w_13530));
  bfr _b_11622(.a(_w_13524),.q(n412_1));
  bfr _b_11621(.a(_w_13523),.q(_w_13524));
  bfr _b_11620(.a(_w_13522),.q(_w_13523));
  bfr _b_11617(.a(_w_13519),.q(_w_13520));
  bfr _b_11616(.a(_w_13518),.q(_w_13519));
  bfr _b_11611(.a(_w_13513),.q(_w_13514));
  bfr _b_11610(.a(_w_13512),.q(n1891));
  bfr _b_13231(.a(_w_15133),.q(_w_15134));
  bfr _b_11606(.a(_w_13508),.q(_w_13509));
  bfr _b_11605(.a(_w_13507),.q(_w_13508));
  bfr _b_11604(.a(_w_13506),.q(_w_13507));
  bfr _b_11602(.a(_w_13504),.q(_w_13505));
  bfr _b_11601(.a(_w_13503),.q(_w_13504));
  bfr _b_11600(.a(_w_13502),.q(_w_13503));
  bfr _b_11599(.a(_w_13501),.q(_w_13502));
  bfr _b_11598(.a(_w_13500),.q(_w_13501));
  bfr _b_11596(.a(_w_13498),.q(_w_13499));
  bfr _b_11595(.a(_w_13497),.q(_w_13498));
  bfr _b_11593(.a(_w_13495),.q(n406_1));
  bfr _b_11592(.a(_w_13494),.q(_w_13495));
  bfr _b_11591(.a(_w_13493),.q(_w_13494));
  bfr _b_11614(.a(_w_13516),.q(_w_13517));
  bfr _b_11590(.a(_w_13492),.q(_w_13493));
  bfr _b_13773(.a(_w_15675),.q(_w_15676));
  bfr _b_11589(.a(_w_13491),.q(N6180));
  bfr _b_11588(.a(_w_13490),.q(_w_13491));
  bfr _b_11587(.a(_w_13489),.q(_w_13490));
  bfr _b_11585(.a(_w_13487),.q(_w_13488));
  bfr _b_11584(.a(_w_13486),.q(_w_13487));
  bfr _b_12562(.a(_w_14464),.q(_w_14465));
  bfr _b_11578(.a(_w_13480),.q(_w_13481));
  bfr _b_11577(.a(_w_13479),.q(_w_13480));
  bfr _b_11575(.a(_w_13477),.q(_w_13478));
  bfr _b_11571(.a(_w_13473),.q(_w_13474));
  bfr _b_12241(.a(_w_14143),.q(_w_14144));
  bfr _b_11568(.a(_w_13470),.q(_w_13471));
  bfr _b_11567(.a(_w_13469),.q(_w_13470));
  bfr _b_11566(.a(_w_13468),.q(_w_13469));
  bfr _b_11564(.a(_w_13466),.q(_w_13467));
  bfr _b_11563(.a(_w_13465),.q(_w_13466));
  bfr _b_11562(.a(_w_13464),.q(_w_13465));
  bfr _b_13296(.a(_w_15198),.q(_w_15199));
  bfr _b_11560(.a(_w_13462),.q(_w_13463));
  bfr _b_11559(.a(_w_13461),.q(_w_13462));
  bfr _b_11557(.a(_w_13459),.q(_w_13460));
  bfr _b_11556(.a(_w_13458),.q(_w_13459));
  bfr _b_11554(.a(_w_13456),.q(_w_13457));
  bfr _b_11553(.a(_w_13455),.q(_w_13456));
  bfr _b_11551(.a(_w_13453),.q(_w_13454));
  bfr _b_11549(.a(_w_13451),.q(_w_13452));
  bfr _b_11548(.a(_w_13450),.q(_w_13451));
  bfr _b_12484(.a(_w_14386),.q(_w_14387));
  bfr _b_11547(.a(_w_13449),.q(_w_13450));
  bfr _b_11545(.a(_w_13447),.q(n1361));
  bfr _b_11543(.a(_w_13445),.q(_w_13446));
  bfr _b_11540(.a(_w_13442),.q(_w_13443));
  bfr _b_13706(.a(_w_15608),.q(_w_15609));
  bfr _b_11539(.a(_w_13441),.q(_w_13442));
  bfr _b_11538(.a(_w_13440),.q(_w_13441));
  bfr _b_13129(.a(_w_15031),.q(_w_15032));
  bfr _b_11536(.a(_w_13438),.q(_w_13439));
  bfr _b_11535(.a(_w_13437),.q(n1843));
  bfr _b_11534(.a(_w_13436),.q(n1772));
  bfr _b_11533(.a(_w_13435),.q(n1355));
  bfr _b_11531(.a(_w_13433),.q(n984));
  bfr _b_11530(.a(_w_13432),.q(n1346));
  bfr _b_11529(.a(_w_13431),.q(n1343));
  bfr _b_12305(.a(_w_14207),.q(_w_14208));
  bfr _b_11527(.a(_w_13429),.q(n484_1));
  bfr _b_11522(.a(_w_13424),.q(N6170));
  bfr _b_11521(.a(_w_13423),.q(_w_13424));
  bfr _b_11520(.a(_w_13422),.q(_w_13423));
  bfr _b_11519(.a(_w_13421),.q(_w_13422));
  bfr _b_11517(.a(_w_13419),.q(_w_13420));
  bfr _b_11821(.a(_w_13723),.q(_w_13724));
  bfr _b_11516(.a(_w_13418),.q(_w_13419));
  bfr _b_11513(.a(_w_13415),.q(_w_13416));
  bfr _b_11512(.a(_w_13414),.q(_w_13415));
  bfr _b_12494(.a(_w_14396),.q(_w_14397));
  bfr _b_11510(.a(_w_13412),.q(_w_13413));
  bfr _b_11508(.a(_w_13410),.q(_w_13411));
  bfr _b_11507(.a(_w_13409),.q(_w_13410));
  bfr _b_13614(.a(_w_15516),.q(_w_15517));
  bfr _b_11506(.a(_w_13408),.q(_w_13409));
  bfr _b_11504(.a(_w_13406),.q(_w_13407));
  bfr _b_11503(.a(_w_13405),.q(_w_13406));
  bfr _b_11502(.a(_w_13404),.q(_w_13405));
  bfr _b_11501(.a(_w_13403),.q(_w_13404));
  bfr _b_11499(.a(_w_13401),.q(_w_13402));
  bfr _b_11498(.a(_w_13400),.q(_w_13401));
  bfr _b_11497(.a(_w_13399),.q(_w_13400));
  bfr _b_13572(.a(_w_15474),.q(_w_15475));
  bfr _b_11496(.a(_w_13398),.q(_w_13399));
  bfr _b_11494(.a(_w_13396),.q(_w_13397));
  bfr _b_11493(.a(_w_13395),.q(_w_13396));
  bfr _b_11489(.a(_w_13391),.q(_w_13392));
  bfr _b_11485(.a(_w_13387),.q(_w_13388));
  bfr _b_11484(.a(_w_13386),.q(_w_13387));
  bfr _b_11481(.a(_w_13383),.q(_w_13384));
  bfr _b_11480(.a(_w_13382),.q(_w_13383));
  bfr _b_11476(.a(_w_13378),.q(_w_13379));
  bfr _b_11474(.a(_w_13376),.q(n1588_1));
  bfr _b_11473(.a(_w_13375),.q(_w_13376));
  bfr _b_11472(.a(_w_13374),.q(_w_13375));
  bfr _b_11471(.a(_w_13373),.q(_w_13374));
  bfr _b_13511(.a(_w_15413),.q(_w_15414));
  bfr _b_11801(.a(_w_13703),.q(_w_13704));
  bfr _b_11468(.a(_w_13370),.q(n268_1));
  bfr _b_11467(.a(_w_13369),.q(_w_13370));
  bfr _b_11466(.a(_w_13368),.q(_w_13369));
  bfr _b_11464(.a(_w_13366),.q(N256_8));
  bfr _b_11463(.a(_w_13365),.q(_w_13366));
  bfr _b_11462(.a(_w_13364),.q(_w_13365));
  bfr _b_11461(.a(_w_13363),.q(_w_13364));
  bfr _b_11460(.a(_w_13362),.q(_w_13363));
  bfr _b_11457(.a(_w_13359),.q(_w_13360));
  bfr _b_11456(.a(_w_13358),.q(_w_13359));
  bfr _b_11455(.a(_w_13357),.q(_w_13358));
  bfr _b_11450(.a(_w_13352),.q(_w_13353));
  bfr _b_11448(.a(_w_13350),.q(_w_13351));
  bfr _b_11751(.a(_w_13653),.q(_w_13654));
  bfr _b_11447(.a(_w_13349),.q(_w_13350));
  bfr _b_11445(.a(_w_13347),.q(_w_13348));
  bfr _b_11443(.a(_w_13345),.q(N2877));
  bfr _b_11442(.a(_w_13344),.q(_w_13345));
  bfr _b_11441(.a(_w_13343),.q(_w_13344));
  bfr _b_13008(.a(_w_14910),.q(_w_14911));
  bfr _b_11440(.a(_w_13342),.q(_w_13343));
  bfr _b_11437(.a(_w_13339),.q(_w_13340));
  bfr _b_12046(.a(_w_13948),.q(n547));
  bfr _b_11435(.a(_w_13337),.q(_w_13338));
  bfr _b_11434(.a(_w_13336),.q(_w_13337));
  bfr _b_11432(.a(_w_13334),.q(_w_13335));
  bfr _b_11431(.a(_w_13333),.q(_w_13334));
  bfr _b_11430(.a(_w_13332),.q(_w_13333));
  bfr _b_11424(.a(_w_13326),.q(_w_13327));
  bfr _b_12178(.a(_w_14080),.q(_w_14081));
  bfr _b_11423(.a(_w_13325),.q(_w_13326));
  bfr _b_12553(.a(_w_14455),.q(_w_14456));
  bfr _b_11421(.a(_w_13323),.q(_w_13324));
  bfr _b_11419(.a(_w_13321),.q(_w_13322));
  bfr _b_11417(.a(_w_13319),.q(_w_13320));
  bfr _b_11411(.a(_w_13313),.q(_w_13314));
  bfr _b_11410(.a(_w_13312),.q(_w_13313));
  bfr _b_11407(.a(_w_13309),.q(_w_13310));
  bfr _b_11406(.a(_w_13308),.q(_w_13309));
  bfr _b_11405(.a(_w_13307),.q(_w_13308));
  bfr _b_11404(.a(_w_13306),.q(_w_13307));
  bfr _b_11402(.a(_w_13304),.q(_w_13305));
  bfr _b_11398(.a(_w_13300),.q(_w_13301));
  bfr _b_11397(.a(_w_13299),.q(_w_13300));
  bfr _b_11396(.a(_w_13298),.q(_w_13299));
  bfr _b_11395(.a(_w_13297),.q(_w_13298));
  bfr _b_11394(.a(_w_13296),.q(_w_13297));
  bfr _b_11393(.a(_w_13295),.q(_w_13296));
  bfr _b_11391(.a(_w_13293),.q(_w_13294));
  bfr _b_11388(.a(_w_13290),.q(_w_13291));
  bfr _b_11387(.a(_w_13289),.q(_w_13290));
  bfr _b_11386(.a(_w_13288),.q(_w_13289));
  bfr _b_11385(.a(_w_13287),.q(_w_13288));
  bfr _b_11380(.a(_w_13282),.q(_w_13283));
  bfr _b_11938(.a(_w_13840),.q(_w_13841));
  bfr _b_11378(.a(_w_13280),.q(_w_13281));
  bfr _b_11377(.a(_w_13279),.q(_w_13280));
  bfr _b_14356(.a(_w_16258),.q(_w_16259));
  bfr _b_11373(.a(_w_13275),.q(_w_13276));
  bfr _b_13875(.a(_w_15777),.q(_w_15778));
  bfr _b_11372(.a(_w_13274),.q(_w_13275));
  bfr _b_11370(.a(_w_13272),.q(_w_13273));
  bfr _b_11368(.a(_w_13270),.q(_w_13271));
  bfr _b_11366(.a(_w_13268),.q(_w_13269));
  bfr _b_11364(.a(_w_13266),.q(_w_13267));
  bfr _b_11359(.a(_w_13261),.q(_w_13262));
  bfr _b_11357(.a(_w_13259),.q(_w_13260));
  bfr _b_11355(.a(_w_13257),.q(_w_13258));
  bfr _b_11354(.a(_w_13256),.q(_w_13257));
  bfr _b_11352(.a(_w_13254),.q(_w_13255));
  bfr _b_11349(.a(_w_13251),.q(_w_13252));
  bfr _b_11347(.a(_w_13249),.q(_w_13250));
  bfr _b_11346(.a(_w_13248),.q(_w_13249));
  bfr _b_11345(.a(_w_13247),.q(_w_13248));
  bfr _b_11344(.a(_w_13246),.q(_w_13247));
  bfr _b_11343(.a(_w_13245),.q(_w_13246));
  bfr _b_11341(.a(_w_13243),.q(_w_13244));
  bfr _b_11338(.a(_w_13240),.q(_w_13241));
  bfr _b_11337(.a(_w_13239),.q(_w_13240));
  bfr _b_11336(.a(_w_13238),.q(_w_13239));
  bfr _b_11335(.a(_w_13237),.q(_w_13238));
  bfr _b_11334(.a(_w_13236),.q(_w_13237));
  bfr _b_11333(.a(_w_13235),.q(_w_13236));
  bfr _b_11332(.a(_w_13234),.q(_w_13235));
  bfr _b_11331(.a(_w_13233),.q(_w_13234));
  bfr _b_11330(.a(_w_13232),.q(_w_13233));
  bfr _b_11329(.a(_w_13231),.q(_w_13232));
  bfr _b_11328(.a(_w_13230),.q(_w_13231));
  bfr _b_11324(.a(_w_13226),.q(_w_13227));
  bfr _b_11322(.a(_w_13224),.q(_w_13225));
  bfr _b_11321(.a(_w_13223),.q(_w_13224));
  bfr _b_11320(.a(_w_13222),.q(_w_13223));
  bfr _b_11318(.a(_w_13220),.q(_w_13221));
  bfr _b_11317(.a(_w_13219),.q(_w_13220));
  bfr _b_11314(.a(_w_13216),.q(_w_13217));
  bfr _b_11313(.a(_w_13215),.q(_w_13216));
  bfr _b_11311(.a(_w_13213),.q(_w_13214));
  bfr _b_11309(.a(_w_13211),.q(_w_13212));
  bfr _b_11308(.a(_w_13210),.q(_w_13211));
  bfr _b_11307(.a(_w_13209),.q(_w_13210));
  bfr _b_11306(.a(_w_13208),.q(_w_13209));
  bfr _b_11305(.a(_w_13207),.q(_w_13208));
  bfr _b_11303(.a(_w_13205),.q(n1307));
  bfr _b_11301(.a(_w_13203),.q(n472_1));
  bfr _b_11298(.a(_w_13200),.q(_w_13201));
  bfr _b_11297(.a(_w_13199),.q(n1292));
  bfr _b_11294(.a(_w_13196),.q(_w_13197));
  bfr _b_11293(.a(_w_13195),.q(_w_13196));
  bfr _b_13554(.a(_w_15456),.q(_w_15457));
  bfr _b_11291(.a(_w_13193),.q(_w_13194));
  bfr _b_11290(.a(_w_13192),.q(_w_13193));
  bfr _b_11289(.a(_w_13191),.q(_w_13192));
  bfr _b_11287(.a(_w_13189),.q(_w_13190));
  bfr _b_11286(.a(_w_13188),.q(_w_13189));
  bfr _b_11737(.a(_w_13639),.q(_w_13640));
  bfr _b_11285(.a(_w_13187),.q(_w_13188));
  bfr _b_11283(.a(_w_13185),.q(_w_13186));
  bfr _b_11281(.a(_w_13183),.q(_w_13184));
  bfr _b_11280(.a(_w_13182),.q(_w_13183));
  bfr _b_13841(.a(_w_15743),.q(_w_15744));
  bfr _b_11279(.a(_w_13181),.q(_w_13182));
  bfr _b_11277(.a(_w_13179),.q(_w_13180));
  bfr _b_11275(.a(_w_13177),.q(_w_13178));
  bfr _b_11274(.a(_w_13176),.q(_w_13177));
  bfr _b_11271(.a(_w_13173),.q(n1289));
  bfr _b_11269(.a(_w_13171),.q(_w_13172));
  bfr _b_11267(.a(_w_13169),.q(n618));
  bfr _b_11265(.a(_w_13167),.q(_w_13168));
  bfr _b_11263(.a(_w_13165),.q(n1286));
  bfr _b_11262(.a(_w_13164),.q(_w_13165));
  bfr _b_11261(.a(_w_13163),.q(_w_13164));
  bfr _b_11257(.a(_w_13159),.q(_w_13160));
  bfr _b_11256(.a(_w_13158),.q(_w_13159));
  bfr _b_11255(.a(_w_13157),.q(_w_13158));
  bfr _b_11254(.a(_w_13156),.q(_w_13157));
  bfr _b_11253(.a(_w_13155),.q(_w_13156));
  bfr _b_11251(.a(_w_13153),.q(_w_13154));
  bfr _b_11249(.a(_w_13151),.q(_w_13152));
  bfr _b_11248(.a(_w_13150),.q(_w_13151));
  bfr _b_11247(.a(_w_13149),.q(n1789));
  bfr _b_11245(.a(_w_13147),.q(_w_13148));
  bfr _b_11244(.a(_w_13146),.q(_w_13147));
  bfr _b_11243(.a(_w_13145),.q(_w_13146));
  bfr _b_11242(.a(_w_13144),.q(_w_13145));
  bfr _b_11241(.a(_w_13143),.q(_w_13144));
  bfr _b_11240(.a(_w_13142),.q(_w_13143));
  bfr _b_11239(.a(_w_13141),.q(_w_13142));
  bfr _b_11236(.a(_w_13138),.q(_w_13139));
  bfr _b_11235(.a(_w_13137),.q(_w_13138));
  bfr _b_11234(.a(_w_13136),.q(n1812));
  bfr _b_11231(.a(_w_13133),.q(_w_13134));
  bfr _b_11230(.a(_w_13132),.q(_w_13133));
  bfr _b_11229(.a(_w_13131),.q(_w_13132));
  bfr _b_11228(.a(_w_13130),.q(_w_13131));
  bfr _b_13503(.a(_w_15405),.q(_w_15406));
  bfr _b_11227(.a(_w_13129),.q(_w_13130));
  bfr _b_11225(.a(_w_13127),.q(_w_13128));
  bfr _b_11224(.a(_w_13126),.q(_w_13127));
  bfr _b_11223(.a(_w_13125),.q(_w_13126));
  bfr _b_11222(.a(_w_13124),.q(_w_13125));
  bfr _b_12451(.a(_w_14353),.q(_w_14354));
  bfr _b_11218(.a(_w_13120),.q(_w_13121));
  bfr _b_11216(.a(_w_13118),.q(_w_13119));
  bfr _b_11214(.a(_w_13116),.q(_w_13117));
  bfr _b_11213(.a(_w_13115),.q(_w_13116));
  bfr _b_11212(.a(_w_13114),.q(_w_13115));
  bfr _b_11208(.a(_w_13110),.q(_w_13111));
  bfr _b_11206(.a(_w_13108),.q(_w_13109));
  bfr _b_11205(.a(_w_13107),.q(_w_13108));
  bfr _b_12889(.a(_w_14791),.q(_w_14792));
  bfr _b_11200(.a(_w_13102),.q(_w_13103));
  bfr _b_11486(.a(_w_13388),.q(_w_13389));
  bfr _b_11199(.a(_w_13101),.q(_w_13102));
  bfr _b_11194(.a(_w_13096),.q(n334));
  bfr _b_11193(.a(_w_13095),.q(n1741_1));
  bfr _b_13119(.a(_w_15021),.q(_w_15022));
  bfr _b_11192(.a(_w_13094),.q(_w_13095));
  bfr _b_11190(.a(_w_13092),.q(_w_13093));
  bfr _b_11189(.a(_w_13091),.q(n1592));
  bfr _b_11188(.a(_w_13090),.q(n388_1));
  bfr _b_11187(.a(_w_13089),.q(_w_13090));
  bfr _b_11409(.a(_w_13311),.q(_w_13312));
  bfr _b_11185(.a(_w_13087),.q(_w_13088));
  bfr _b_11183(.a(_w_13085),.q(_w_13086));
  bfr _b_11177(.a(_w_13079),.q(_w_13080));
  bfr _b_11176(.a(_w_13078),.q(n1270));
  bfr _b_11175(.a(_w_13077),.q(_w_13078));
  bfr _b_11174(.a(_w_13076),.q(_w_13077));
  bfr _b_11173(.a(_w_13075),.q(_w_13076));
  bfr _b_11171(.a(_w_13073),.q(_w_13074));
  bfr _b_11170(.a(_w_13072),.q(_w_13073));
  bfr _b_11179(.a(_w_13081),.q(_w_13082));
  bfr _b_11169(.a(_w_13071),.q(_w_13072));
  bfr _b_11168(.a(_w_13070),.q(_w_13071));
  bfr _b_12084(.a(_w_13986),.q(_w_13987));
  bfr _b_11166(.a(_w_13068),.q(_w_13069));
  bfr _b_11164(.a(_w_13066),.q(_w_13067));
  bfr _b_11163(.a(_w_13065),.q(_w_13066));
  bfr _b_11161(.a(_w_13063),.q(_w_13064));
  bfr _b_11160(.a(_w_13062),.q(N6270));
  bfr _b_11159(.a(_w_13061),.q(_w_13062));
  bfr _b_11156(.a(_w_13058),.q(_w_13059));
  bfr _b_14061(.a(_w_15963),.q(_w_15964));
  bfr _b_11155(.a(_w_13057),.q(_w_13058));
  bfr _b_11153(.a(_w_13055),.q(_w_13056));
  bfr _b_11152(.a(_w_13054),.q(n244));
  bfr _b_11148(.a(_w_13050),.q(_w_13051));
  bfr _b_11147(.a(_w_13049),.q(_w_13050));
  bfr _b_14019(.a(_w_15921),.q(_w_15922));
  bfr _b_11145(.a(_w_13047),.q(n760_1));
  bfr _b_13313(.a(_w_15215),.q(_w_15216));
  bfr _b_11144(.a(_w_13046),.q(_w_13047));
  bfr _b_11143(.a(_w_13045),.q(_w_13046));
  bfr _b_11142(.a(_w_13044),.q(_w_13045));
  bfr _b_11141(.a(_w_13043),.q(n1261));
  bfr _b_11136(.a(_w_13038),.q(n704));
  bfr _b_11135(.a(_w_13037),.q(n1255));
  bfr _b_11134(.a(_w_13036),.q(n1570_1));
  bfr _b_11133(.a(_w_13035),.q(_w_13036));
  bfr _b_11132(.a(_w_13034),.q(_w_13035));
  bfr _b_11131(.a(_w_13033),.q(_w_13034));
  bfr _b_11130(.a(_w_13032),.q(n1252));
  bfr _b_11129(.a(_w_13031),.q(n1529));
  bfr _b_11128(.a(_w_13030),.q(_w_13031));
  bfr _b_11127(.a(_w_13029),.q(_w_13030));
  bfr _b_11126(.a(_w_13028),.q(_w_13029));
  bfr _b_11125(.a(_w_13027),.q(_w_13028));
  bfr _b_12177(.a(_w_14079),.q(_w_14080));
  bfr _b_11124(.a(_w_13026),.q(_w_13027));
  bfr _b_12944(.a(_w_14846),.q(_w_14847));
  bfr _b_11123(.a(_w_13025),.q(_w_13026));
  bfr _b_11122(.a(_w_13024),.q(_w_13025));
  bfr _b_11120(.a(_w_13022),.q(_w_13023));
  bfr _b_13512(.a(_w_15414),.q(_w_15415));
  bfr _b_11118(.a(_w_13020),.q(_w_13021));
  bfr _b_11117(.a(_w_13019),.q(_w_13020));
  bfr _b_11113(.a(_w_13015),.q(n1331));
  bfr _b_11112(.a(_w_13014),.q(n1249));
  bfr _b_11111(.a(_w_13013),.q(n1714));
  bfr _b_11109(.a(_w_13011),.q(n788));
  bfr _b_11107(.a(_w_13009),.q(n881_1));
  bfr _b_11106(.a(_w_13008),.q(_w_13009));
  bfr _b_11105(.a(_w_13007),.q(_w_13008));
  bfr _b_11104(.a(_w_13006),.q(_w_13007));
  bfr _b_11103(.a(_w_13005),.q(n1222));
  bfr _b_11102(.a(_w_13004),.q(n1219));
  bfr _b_11101(.a(_w_13003),.q(n739));
  bfr _b_11095(.a(_w_12997),.q(_w_12998));
  bfr _b_11093(.a(_w_12995),.q(_w_12996));
  bfr _b_11091(.a(_w_12993),.q(_w_12994));
  bfr _b_11090(.a(_w_12992),.q(_w_12993));
  bfr _b_11089(.a(_w_12991),.q(_w_12992));
  bfr _b_11088(.a(_w_12990),.q(_w_12991));
  bfr _b_11085(.a(_w_12987),.q(_w_12988));
  bfr _b_11084(.a(_w_12986),.q(_w_12987));
  bfr _b_11083(.a(_w_12985),.q(_w_12986));
  bfr _b_11080(.a(_w_12982),.q(_w_12983));
  bfr _b_11079(.a(_w_12981),.q(_w_12982));
  bfr _b_11076(.a(_w_12978),.q(n1186));
  bfr _b_11075(.a(_w_12977),.q(_w_12978));
  bfr _b_11074(.a(_w_12976),.q(_w_12977));
  bfr _b_11073(.a(_w_12975),.q(_w_12976));
  bfr _b_11072(.a(_w_12974),.q(_w_12975));
  bfr _b_11071(.a(_w_12973),.q(_w_12974));
  bfr _b_11797(.a(_w_13699),.q(_w_13700));
  bfr _b_11070(.a(_w_12972),.q(_w_12973));
  bfr _b_11067(.a(_w_12969),.q(_w_12970));
  bfr _b_11066(.a(_w_12968),.q(_w_12969));
  bfr _b_12258(.a(_w_14160),.q(_w_14161));
  bfr _b_11064(.a(_w_12966),.q(_w_12967));
  bfr _b_11058(.a(_w_12960),.q(_w_12961));
  bfr _b_13759(.a(_w_15661),.q(_w_15662));
  bfr _b_12715(.a(_w_14617),.q(_w_14618));
  bfr _b_11893(.a(_w_13795),.q(_w_13796));
  bfr _b_11055(.a(_w_12957),.q(_w_12958));
  bfr _b_11052(.a(_w_12954),.q(_w_12955));
  bfr _b_11051(.a(_w_12953),.q(_w_12954));
  bfr _b_11047(.a(_w_12949),.q(_w_12950));
  bfr _b_11046(.a(_w_12948),.q(_w_12949));
  bfr _b_11045(.a(_w_12947),.q(_w_12948));
  bfr _b_11044(.a(_w_12946),.q(_w_12947));
  bfr _b_11043(.a(_w_12945),.q(_w_12946));
  bfr _b_11042(.a(_w_12944),.q(_w_12945));
  bfr _b_11041(.a(_w_12943),.q(_w_12944));
  bfr _b_11040(.a(_w_12942),.q(_w_12943));
  bfr _b_11037(.a(_w_12939),.q(_w_12940));
  bfr _b_11032(.a(_w_12934),.q(_w_12935));
  bfr _b_11031(.a(_w_12933),.q(_w_12934));
  bfr _b_11030(.a(_w_12932),.q(_w_12933));
  bfr _b_11029(.a(_w_12931),.q(_w_12932));
  bfr _b_11028(.a(_w_12930),.q(_w_12931));
  bfr _b_11025(.a(_w_12927),.q(_w_12928));
  bfr _b_12411(.a(_w_14313),.q(_w_14314));
  bfr _b_11024(.a(_w_12926),.q(_w_12927));
  bfr _b_11023(.a(_w_12925),.q(_w_12926));
  bfr _b_11182(.a(_w_13084),.q(_w_13085));
  bfr _b_11020(.a(_w_12922),.q(_w_12923));
  bfr _b_11017(.a(_w_12919),.q(_w_12920));
  bfr _b_11015(.a(_w_12917),.q(_w_12918));
  bfr _b_11013(.a(_w_12915),.q(_w_12916));
  bfr _b_11011(.a(_w_12913),.q(n1310));
  bfr _b_12672(.a(_w_14574),.q(_w_14575));
  bfr _b_11009(.a(_w_12911),.q(_w_12912));
  bfr _b_11034(.a(_w_12936),.q(_w_12937));
  bfr _b_11007(.a(_w_12909),.q(_w_12910));
  bfr _b_11005(.a(_w_12907),.q(_w_12908));
  bfr _b_11004(.a(_w_12906),.q(_w_12907));
  bfr _b_11003(.a(_w_12905),.q(_w_12906));
  bfr _b_11000(.a(_w_12902),.q(_w_12903));
  bfr _b_10998(.a(_w_12900),.q(_w_12901));
  bfr _b_10996(.a(_w_12898),.q(_w_12899));
  bfr _b_10993(.a(_w_12895),.q(_w_12896));
  bfr _b_12755(.a(_w_14657),.q(n1852));
  bfr _b_10991(.a(_w_12893),.q(_w_12894));
  bfr _b_10990(.a(_w_12892),.q(_w_12893));
  bfr _b_10989(.a(_w_12891),.q(_w_12892));
  bfr _b_10988(.a(_w_12890),.q(_w_12891));
  bfr _b_10987(.a(_w_12889),.q(_w_12890));
  bfr _b_10984(.a(_w_12886),.q(_w_12887));
  bfr _b_10982(.a(_w_12884),.q(_w_12885));
  bfr _b_10981(.a(_w_12883),.q(_w_12884));
  bfr _b_13413(.a(_w_15315),.q(n342_1));
  bfr _b_10980(.a(_w_12882),.q(_w_12883));
  bfr _b_10978(.a(_w_12880),.q(_w_12881));
  bfr _b_10976(.a(_w_12878),.q(_w_12879));
  bfr _b_10972(.a(_w_12874),.q(_w_12875));
  bfr _b_11146(.a(_w_13048),.q(n1264));
  bfr _b_10971(.a(_w_12873),.q(_w_12874));
  bfr _b_10969(.a(_w_12871),.q(_w_12872));
  bfr _b_10967(.a(_w_12869),.q(_w_12870));
  bfr _b_13607(.a(_w_15509),.q(_w_15510));
  bfr _b_10966(.a(_w_12868),.q(_w_12869));
  bfr _b_14252(.a(_w_16154),.q(_w_16155));
  bfr _b_10964(.a(_w_12866),.q(_w_12867));
  bfr _b_10961(.a(_w_12863),.q(n1156));
  bfr _b_10959(.a(_w_12861),.q(_w_12862));
  bfr _b_10958(.a(_w_12860),.q(N86_6));
  bfr _b_10957(.a(_w_12859),.q(_w_12860));
  bfr _b_10956(.a(_w_12858),.q(n1153));
  bfr _b_11721(.a(_w_13623),.q(_w_13624));
  bfr _b_10955(.a(_w_12857),.q(n1501));
  bfr _b_10952(.a(_w_12854),.q(n1392_1));
  bfr _b_12489(.a(_w_14391),.q(_w_14392));
  bfr _b_10951(.a(_w_12853),.q(_w_12854));
  bfr _b_10949(.a(_w_12851),.q(_w_12852));
  bfr _b_10948(.a(_w_12850),.q(n1144));
  bfr _b_10947(.a(_w_12849),.q(n464));
  bfr _b_10945(.a(_w_12847),.q(_w_12848));
  bfr _b_10943(.a(_w_12845),.q(_w_12846));
  bfr _b_13672(.a(_w_15574),.q(_w_15575));
  bfr _b_10942(.a(_w_12844),.q(_w_12845));
  bfr _b_10940(.a(_w_12842),.q(_w_12843));
  bfr _b_10938(.a(_w_12840),.q(n571));
  bfr _b_10934(.a(_w_12836),.q(_w_12837));
  bfr _b_10931(.a(_w_12833),.q(_w_12834));
  bfr _b_10930(.a(_w_12832),.q(_w_12833));
  bfr _b_10929(.a(_w_12831),.q(_w_12832));
  bfr _b_10926(.a(_w_12828),.q(_w_12829));
  bfr _b_10925(.a(_w_12827),.q(_w_12828));
  bfr _b_10923(.a(_w_12825),.q(n903));
  bfr _b_10922(.a(_w_12824),.q(n1828));
  bfr _b_13818(.a(_w_15720),.q(_w_15721));
  bfr _b_10921(.a(_w_12823),.q(n1509_1));
  bfr _b_10920(.a(_w_12822),.q(_w_12823));
  bfr _b_11211(.a(_w_13113),.q(_w_13114));
  bfr _b_10919(.a(_w_12821),.q(_w_12822));
  bfr _b_10917(.a(_w_12819),.q(N5308));
  bfr _b_10916(.a(_w_12818),.q(_w_12819));
  bfr _b_10913(.a(_w_12815),.q(_w_12816));
  bfr _b_10910(.a(_w_12812),.q(_w_12813));
  bfr _b_11579(.a(_w_13481),.q(_w_13482));
  bfr _b_10909(.a(_w_12811),.q(_w_12812));
  bfr _b_10908(.a(_w_12810),.q(_w_12811));
  bfr _b_10903(.a(_w_12805),.q(_w_12806));
  bfr _b_10902(.a(_w_12804),.q(_w_12805));
  bfr _b_10901(.a(_w_12803),.q(_w_12804));
  bfr _b_10894(.a(_w_12796),.q(_w_12797));
  bfr _b_10893(.a(_w_12795),.q(_w_12796));
  bfr _b_10892(.a(_w_12794),.q(_w_12795));
  bfr _b_10992(.a(_w_12894),.q(_w_12895));
  bfr _b_10891(.a(_w_12793),.q(_w_12794));
  bfr _b_10889(.a(_w_12791),.q(_w_12792));
  bfr _b_10888(.a(_w_12790),.q(_w_12791));
  bfr _b_10886(.a(_w_12788),.q(_w_12789));
  bfr _b_10885(.a(_w_12787),.q(_w_12788));
  bfr _b_10883(.a(_w_12785),.q(_w_12786));
  bfr _b_10882(.a(_w_12784),.q(_w_12785));
  bfr _b_13255(.a(_w_15157),.q(_w_15158));
  bfr _b_12077(.a(_w_13979),.q(n1651));
  bfr _b_10881(.a(_w_12783),.q(_w_12784));
  bfr _b_10880(.a(_w_12782),.q(_w_12783));
  bfr _b_10877(.a(_w_12779),.q(_w_12780));
  bfr _b_11570(.a(_w_13472),.q(_w_13473));
  bfr _b_10876(.a(_w_12778),.q(_w_12779));
  bfr _b_10875(.a(_w_12777),.q(_w_12778));
  bfr _b_10873(.a(_w_12775),.q(_w_12776));
  bfr _b_10870(.a(_w_12772),.q(_w_12773));
  bfr _b_10869(.a(_w_12771),.q(_w_12772));
  bfr _b_10868(.a(_w_12770),.q(_w_12771));
  bfr _b_10866(.a(_w_12768),.q(_w_12769));
  bfr _b_10863(.a(_w_12765),.q(_w_12766));
  bfr _b_10862(.a(_w_12764),.q(_w_12765));
  bfr _b_10860(.a(_w_12762),.q(_w_12763));
  bfr _b_10859(.a(_w_12761),.q(_w_12762));
  bfr _b_11197(.a(_w_13099),.q(_w_13100));
  bfr _b_10858(.a(_w_12760),.q(_w_12761));
  bfr _b_10857(.a(_w_12759),.q(_w_12760));
  bfr _b_10854(.a(_w_12756),.q(_w_12757));
  bfr _b_10853(.a(_w_12755),.q(_w_12756));
  bfr _b_10852(.a(_w_12754),.q(_w_12755));
  bfr _b_10851(.a(_w_12753),.q(_w_12754));
  bfr _b_10847(.a(_w_12749),.q(_w_12750));
  bfr _b_10845(.a(_w_12747),.q(_w_12748));
  bfr _b_10843(.a(_w_12745),.q(_w_12746));
  bfr _b_12578(.a(_w_14480),.q(_w_14481));
  bfr _b_10842(.a(_w_12744),.q(_w_12745));
  bfr _b_11371(.a(_w_13273),.q(_w_13274));
  bfr _b_10841(.a(_w_12743),.q(_w_12744));
  bfr _b_10840(.a(_w_12742),.q(_w_12743));
  bfr _b_10838(.a(_w_12740),.q(_w_12741));
  bfr _b_10836(.a(_w_12738),.q(_w_12739));
  bfr _b_11682(.a(_w_13584),.q(_w_13585));
  bfr _b_10833(.a(_w_12735),.q(N273_19));
  bfr _b_10832(.a(_w_12734),.q(_w_12735));
  bfr _b_10831(.a(_w_12733),.q(_w_12734));
  bfr _b_10830(.a(_w_12732),.q(n404));
  bfr _b_10829(.a(_w_12731),.q(n550));
  bfr _b_10826(.a(_w_12728),.q(n534));
  bfr _b_10824(.a(_w_12726),.q(_w_12727));
  bfr _b_10822(.a(_w_12724),.q(_w_12725));
  bfr _b_10821(.a(_w_12723),.q(_w_12724));
  bfr _b_10817(.a(_w_12719),.q(_w_12720));
  bfr _b_10816(.a(_w_12718),.q(_w_12719));
  bfr _b_10815(.a(_w_12717),.q(_w_12718));
  bfr _b_10811(.a(_w_12713),.q(_w_12714));
  bfr _b_10809(.a(_w_12711),.q(_w_12712));
  bfr _b_10808(.a(_w_12710),.q(_w_12711));
  bfr _b_10807(.a(_w_12709),.q(_w_12710));
  bfr _b_10805(.a(_w_12707),.q(_w_12708));
  bfr _b_10804(.a(_w_12706),.q(_w_12707));
  bfr _b_11663(.a(_w_13565),.q(n1297_1));
  bfr _b_10803(.a(_w_12705),.q(_w_12706));
  bfr _b_10801(.a(_w_12703),.q(_w_12704));
  bfr _b_10799(.a(_w_12701),.q(_w_12702));
  bfr _b_10797(.a(_w_12699),.q(_w_12700));
  bfr _b_10796(.a(_w_12698),.q(_w_12699));
  bfr _b_12757(.a(_w_14659),.q(_w_14660));
  bfr _b_10795(.a(_w_12697),.q(_w_12698));
  bfr _b_10794(.a(_w_12696),.q(N86_13));
  bfr _b_12040(.a(_w_13942),.q(n1577));
  bfr _b_10792(.a(_w_12694),.q(_w_12695));
  bfr _b_10786(.a(_w_12688),.q(N6123));
  bfr _b_14245(.a(_w_16147),.q(_w_16148));
  bfr _b_10785(.a(_w_12687),.q(_w_12688));
  bfr _b_10783(.a(_w_12685),.q(_w_12686));
  bfr _b_10782(.a(_w_12684),.q(_w_12685));
  bfr _b_10781(.a(_w_12683),.q(_w_12684));
  bfr _b_10778(.a(_w_12680),.q(_w_12681));
  bfr _b_10777(.a(_w_12679),.q(_w_12680));
  bfr _b_10775(.a(_w_12677),.q(_w_12678));
  bfr _b_10773(.a(_w_12675),.q(_w_12676));
  bfr _b_10770(.a(_w_12672),.q(_w_12673));
  bfr _b_10769(.a(_w_12671),.q(_w_12672));
  bfr _b_10767(.a(_w_12669),.q(_w_12670));
  bfr _b_10765(.a(_w_12667),.q(_w_12668));
  bfr _b_10763(.a(_w_12665),.q(_w_12666));
  bfr _b_10760(.a(_w_12662),.q(_w_12663));
  bfr _b_10759(.a(_w_12661),.q(_w_12662));
  bfr _b_10756(.a(_w_12658),.q(_w_12659));
  bfr _b_10754(.a(_w_12656),.q(_w_12657));
  bfr _b_10751(.a(_w_12653),.q(_w_12654));
  bfr _b_10750(.a(_w_12652),.q(_w_12653));
  bfr _b_10749(.a(_w_12651),.q(_w_12652));
  bfr _b_10748(.a(_w_12650),.q(_w_12651));
  bfr _b_10747(.a(_w_12649),.q(_w_12650));
  bfr _b_10746(.a(_w_12648),.q(_w_12649));
  bfr _b_10758(.a(_w_12660),.q(_w_12661));
  bfr _b_10745(.a(_w_12647),.q(_w_12648));
  bfr _b_10744(.a(_w_12646),.q(_w_12647));
  bfr _b_10741(.a(_w_12643),.q(_w_12644));
  bfr _b_10740(.a(_w_12642),.q(_w_12643));
  bfr _b_10739(.a(_w_12641),.q(_w_12642));
  bfr _b_10736(.a(_w_12638),.q(_w_12639));
  bfr _b_10735(.a(_w_12637),.q(_w_12638));
  bfr _b_10734(.a(_w_12636),.q(_w_12637));
  bfr _b_10731(.a(_w_12633),.q(_w_12634));
  bfr _b_10730(.a(_w_12632),.q(_w_12633));
  bfr _b_10729(.a(_w_12631),.q(_w_12632));
  bfr _b_10725(.a(_w_12627),.q(_w_12628));
  bfr _b_12566(.a(_w_14468),.q(_w_14469));
  bfr _b_10724(.a(_w_12626),.q(_w_12627));
  bfr _b_10723(.a(_w_12625),.q(_w_12626));
  bfr _b_10722(.a(_w_12624),.q(_w_12625));
  bfr _b_11509(.a(_w_13411),.q(_w_13412));
  bfr _b_10721(.a(_w_12623),.q(_w_12624));
  bfr _b_10720(.a(_w_12622),.q(_w_12623));
  bfr _b_10719(.a(_w_12621),.q(_w_12622));
  bfr _b_10715(.a(_w_12617),.q(_w_12618));
  bfr _b_10714(.a(_w_12616),.q(n800));
  bfr _b_10713(.a(_w_12615),.q(N4946));
  bfr _b_10711(.a(_w_12613),.q(_w_12614));
  bfr _b_10710(.a(_w_12612),.q(_w_12613));
  bfr _b_10709(.a(_w_12611),.q(_w_12612));
  bfr _b_13110(.a(_w_15012),.q(_w_15013));
  bfr _b_10706(.a(_w_12608),.q(_w_12609));
  bfr _b_10705(.a(_w_12607),.q(_w_12608));
  bfr _b_10704(.a(_w_12606),.q(_w_12607));
  bfr _b_10702(.a(_w_12604),.q(_w_12605));
  bfr _b_10700(.a(_w_12602),.q(_w_12603));
  bfr _b_10698(.a(_w_12600),.q(_w_12601));
  bfr _b_10697(.a(_w_12599),.q(_w_12600));
  bfr _b_10696(.a(_w_12598),.q(_w_12599));
  bfr _b_10694(.a(_w_12596),.q(_w_12597));
  bfr _b_14186(.a(_w_16088),.q(_w_16089));
  bfr _b_10692(.a(_w_12594),.q(_w_12595));
  bfr _b_10691(.a(_w_12593),.q(_w_12594));
  bfr _b_13218(.a(_w_15120),.q(_w_15121));
  bfr _b_10689(.a(_w_12591),.q(_w_12592));
  bfr _b_10686(.a(_w_12588),.q(_w_12589));
  bfr _b_10682(.a(_w_12584),.q(_w_12585));
  bfr _b_10681(.a(_w_12583),.q(_w_12584));
  bfr _b_10679(.a(_w_12581),.q(_w_12582));
  bfr _b_10677(.a(_w_12579),.q(_w_12580));
  bfr _b_10676(.a(_w_12578),.q(_w_12579));
  bfr _b_10674(.a(_w_12576),.q(_w_12577));
  bfr _b_12598(.a(_w_14500),.q(_w_14501));
  bfr _b_10673(.a(_w_12575),.q(_w_12576));
  bfr _b_10672(.a(_w_12574),.q(_w_12575));
  bfr _b_10671(.a(_w_12573),.q(_w_12574));
  bfr _b_12964(.a(_w_14866),.q(_w_14867));
  bfr _b_10668(.a(_w_12570),.q(_w_12571));
  bfr _b_10666(.a(_w_12568),.q(_w_12569));
  bfr _b_10665(.a(_w_12567),.q(_w_12568));
  bfr _b_10663(.a(_w_12565),.q(_w_12566));
  bfr _b_10662(.a(_w_12564),.q(_w_12565));
  bfr _b_10660(.a(_w_12562),.q(_w_12563));
  bfr _b_10659(.a(_w_12561),.q(_w_12562));
  bfr _b_10655(.a(_w_12557),.q(_w_12558));
  bfr _b_10654(.a(_w_12556),.q(_w_12557));
  bfr _b_10652(.a(_w_12554),.q(_w_12555));
  bfr _b_10651(.a(_w_12553),.q(_w_12554));
  bfr _b_10650(.a(_w_12552),.q(_w_12553));
  bfr _b_11717(.a(_w_13619),.q(_w_13620));
  bfr _b_10647(.a(_w_12549),.q(_w_12550));
  bfr _b_10646(.a(_w_12548),.q(_w_12549));
  bfr _b_10645(.a(_w_12547),.q(_w_12548));
  bfr _b_10643(.a(_w_12545),.q(_w_12546));
  bfr _b_10640(.a(_w_12542),.q(_w_12543));
  bfr _b_10639(.a(_w_12541),.q(_w_12542));
  bfr _b_10637(.a(_w_12539),.q(_w_12540));
  bfr _b_10636(.a(_w_12538),.q(_w_12539));
  bfr _b_10635(.a(_w_12537),.q(_w_12538));
  bfr _b_10630(.a(_w_12532),.q(_w_12533));
  bfr _b_10628(.a(_w_12530),.q(_w_12531));
  bfr _b_10627(.a(_w_12529),.q(_w_12530));
  bfr _b_10626(.a(_w_12528),.q(_w_12529));
  bfr _b_10625(.a(_w_12527),.q(_w_12528));
  bfr _b_10624(.a(_w_12526),.q(_w_12527));
  bfr _b_10623(.a(_w_12525),.q(_w_12526));
  bfr _b_10619(.a(_w_12521),.q(_w_12522));
  bfr _b_10617(.a(_w_12519),.q(_w_12520));
  bfr _b_10615(.a(_w_12517),.q(n95));
  bfr _b_10613(.a(_w_12515),.q(n319));
  bfr _b_10612(.a(_w_12514),.q(n1798));
  bfr _b_10611(.a(_w_12513),.q(n996));
  bfr _b_10610(.a(_w_12512),.q(n503));
  bfr _b_10608(.a(_w_12510),.q(_w_12511));
  bfr _b_10607(.a(_w_12509),.q(_w_12510));
  bfr _b_10604(.a(_w_12506),.q(n446));
  bfr _b_10603(.a(_w_12505),.q(_w_12506));
  bfr _b_10602(.a(_w_12504),.q(_w_12505));
  bfr _b_10737(.a(_w_12639),.q(_w_12640));
  bfr _b_10599(.a(_w_12501),.q(_w_12502));
  bfr _b_10597(.a(_w_12499),.q(_w_12500));
  bfr _b_10596(.a(_w_12498),.q(_w_12499));
  bfr _b_11433(.a(_w_13335),.q(_w_13336));
  bfr _b_10595(.a(_w_12497),.q(_w_12498));
  bfr _b_13048(.a(_w_14950),.q(n1881_1));
  bfr _b_10594(.a(_w_12496),.q(_w_12497));
  bfr _b_10593(.a(_w_12495),.q(_w_12496));
  bfr _b_10590(.a(_w_12492),.q(_w_12493));
  bfr _b_10586(.a(_w_12488),.q(n230));
  bfr _b_10585(.a(_w_12487),.q(n58));
  bfr _b_10584(.a(_w_12486),.q(n458));
  bfr _b_10582(.a(_w_12484),.q(_w_12485));
  bfr _b_10578(.a(_w_12480),.q(_w_12481));
  bfr _b_10638(.a(_w_12540),.q(_w_12541));
  bfr _b_10576(.a(_w_12478),.q(_w_12479));
  bfr _b_10575(.a(_w_12477),.q(N35_15));
  bfr _b_10572(.a(_w_12474),.q(_w_12475));
  bfr _b_10570(.a(_w_12472),.q(_w_12473));
  bfr _b_10569(.a(_w_12471),.q(_w_12472));
  bfr _b_14288(.a(_w_16190),.q(_w_16191));
  bfr _b_10568(.a(_w_12470),.q(_w_12471));
  bfr _b_10567(.a(_w_12469),.q(_w_12470));
  bfr _b_10566(.a(_w_12468),.q(_w_12469));
  bfr _b_10565(.a(_w_12467),.q(_w_12468));
  bfr _b_10564(.a(_w_12466),.q(_w_12467));
  bfr _b_10937(.a(_w_12839),.q(n909));
  bfr _b_10563(.a(_w_12465),.q(N35_14));
  bfr _b_10562(.a(_w_12464),.q(_w_12465));
  bfr _b_10560(.a(_w_12462),.q(_w_12463));
  bfr _b_10559(.a(_w_12461),.q(_w_12462));
  bfr _b_10558(.a(_w_12460),.q(_w_12461));
  bfr _b_10557(.a(_w_12459),.q(_w_12460));
  bfr _b_10556(.a(_w_12458),.q(_w_12459));
  bfr _b_10555(.a(_w_12457),.q(_w_12458));
  bfr _b_10554(.a(_w_12456),.q(_w_12457));
  bfr _b_10553(.a(_w_12455),.q(_w_12456));
  bfr _b_10551(.a(_w_12453),.q(N35_13));
  bfr _b_10550(.a(_w_12452),.q(_w_12453));
  bfr _b_10548(.a(_w_12450),.q(_w_12451));
  bfr _b_10545(.a(_w_12447),.q(_w_12448));
  bfr _b_10543(.a(_w_12445),.q(n1321_1));
  bfr _b_10542(.a(_w_12444),.q(_w_12445));
  bfr _b_10539(.a(_w_12441),.q(n448));
  bfr _b_12878(.a(_w_14780),.q(_w_14781));
  bfr _b_10536(.a(_w_12438),.q(_w_12439));
  bfr _b_10534(.a(_w_12436),.q(_w_12437));
  bfr _b_11157(.a(_w_13059),.q(_w_13060));
  bfr _b_10533(.a(_w_12435),.q(_w_12436));
  bfr _b_10532(.a(_w_12434),.q(_w_12435));
  bfr _b_10531(.a(_w_12433),.q(n318_1));
  bfr _b_10529(.a(_w_12431),.q(_w_12432));
  bfr _b_10528(.a(_w_12430),.q(_w_12431));
  bfr _b_10527(.a(_w_12429),.q(n336_1));
  bfr _b_10526(.a(_w_12428),.q(_w_12429));
  bfr _b_10525(.a(_w_12427),.q(_w_12428));
  bfr _b_13999(.a(_w_15901),.q(_w_15902));
  bfr _b_10524(.a(_w_12426),.q(_w_12427));
  bfr _b_10521(.a(_w_12423),.q(n1276));
  bfr _b_10519(.a(_w_12421),.q(_w_12422));
  bfr _b_10518(.a(_w_12420),.q(_w_12421));
  bfr _b_13084(.a(_w_14986),.q(_w_14987));
  bfr _b_10517(.a(_w_12419),.q(_w_12420));
  bfr _b_10513(.a(_w_12415),.q(_w_12416));
  bfr _b_10512(.a(_w_12414),.q(_w_12415));
  bfr _b_10511(.a(_w_12413),.q(_w_12414));
  bfr _b_10509(.a(_w_12411),.q(n83));
  bfr _b_10508(.a(_w_12410),.q(n1441));
  bfr _b_10507(.a(_w_12409),.q(n490_1));
  bfr _b_10506(.a(_w_12408),.q(_w_12409));
  bfr _b_10503(.a(_w_12405),.q(n425));
  bfr _b_12698(.a(_w_14600),.q(_w_14601));
  bfr _b_10501(.a(_w_12403),.q(_w_12404));
  bfr _b_10500(.a(_w_12402),.q(_w_12403));
  bfr _b_10498(.a(_w_12400),.q(n1683));
  bfr _b_10497(.a(_w_12399),.q(_w_12400));
  bfr _b_10496(.a(_w_12398),.q(_w_12399));
  bfr _b_10494(.a(_w_12396),.q(n981));
  bfr _b_10492(.a(_w_12394),.q(_w_12395));
  bfr _b_10491(.a(_w_12393),.q(_w_12394));
  bfr _b_10490(.a(_w_12392),.q(_w_12393));
  bfr _b_13357(.a(_w_15259),.q(_w_15260));
  bfr _b_10488(.a(_w_12390),.q(_w_12391));
  bfr _b_10487(.a(_w_12389),.q(_w_12390));
  bfr _b_10486(.a(_w_12388),.q(_w_12389));
  bfr _b_11807(.a(_w_13709),.q(_w_13710));
  bfr _b_10484(.a(_w_12386),.q(_w_12387));
  bfr _b_10483(.a(_w_12385),.q(_w_12386));
  bfr _b_13866(.a(_w_15768),.q(_w_15769));
  bfr _b_10480(.a(_w_12382),.q(_w_12383));
  bfr _b_10479(.a(_w_12381),.q(_w_12382));
  bfr _b_10477(.a(_w_12379),.q(_w_12380));
  bfr _b_10476(.a(_w_12378),.q(_w_12379));
  bfr _b_10475(.a(_w_12377),.q(_w_12378));
  bfr _b_10474(.a(_w_12376),.q(_w_12377));
  bfr _b_10473(.a(_w_12375),.q(_w_12376));
  bfr _b_10468(.a(_w_12370),.q(_w_12371));
  bfr _b_10466(.a(_w_12368),.q(_w_12369));
  bfr _b_10464(.a(_w_12366),.q(n850));
  bfr _b_10462(.a(_w_12364),.q(n491));
  bfr _b_14292(.a(_w_16194),.q(_w_16195));
  bfr _b_13648(.a(_w_15550),.q(_w_15551));
  bfr _b_10460(.a(_w_12362),.q(_w_12363));
  bfr _b_10459(.a(_w_12361),.q(_w_12362));
  bfr _b_10457(.a(_w_12359),.q(n1082));
  bfr _b_13567(.a(_w_15469),.q(_w_15470));
  bfr _b_10456(.a(_w_12358),.q(_w_12359));
  bfr _b_10455(.a(_w_12357),.q(_w_12358));
  bfr _b_10454(.a(_w_12356),.q(n1699));
  bfr _b_10451(.a(_w_12353),.q(_w_12354));
  bfr _b_10449(.a(_w_12351),.q(_w_12352));
  bfr _b_10448(.a(_w_12350),.q(_w_12351));
  bfr _b_10447(.a(_w_12349),.q(_w_12350));
  bfr _b_10446(.a(_w_12348),.q(_w_12349));
  bfr _b_10443(.a(_w_12345),.q(_w_12346));
  bfr _b_10440(.a(_w_12342),.q(_w_12343));
  bfr _b_13027(.a(_w_14929),.q(_w_14930));
  bfr _b_12151(.a(_w_14053),.q(_w_14054));
  bfr _b_10437(.a(_w_12339),.q(_w_12340));
  bfr _b_10436(.a(_w_12338),.q(_w_12339));
  bfr _b_10434(.a(_w_12336),.q(_w_12337));
  bfr _b_10432(.a(_w_12334),.q(n1216));
  bfr _b_13779(.a(_w_15681),.q(_w_15682));
  bfr _b_11018(.a(_w_12920),.q(_w_12921));
  bfr _b_10439(.a(_w_12341),.q(_w_12342));
  bfr _b_10430(.a(_w_12332),.q(n242));
  bfr _b_12793(.a(_w_14695),.q(_w_14696));
  bfr _b_10429(.a(_w_12331),.q(_w_12332));
  bfr _b_10427(.a(_w_12329),.q(_w_12330));
  bfr _b_10426(.a(_w_12328),.q(_w_12329));
  bfr _b_10423(.a(_w_12325),.q(_w_12326));
  bfr _b_10421(.a(_w_12323),.q(_w_12324));
  bfr _b_10420(.a(_w_12322),.q(_w_12323));
  bfr _b_10416(.a(_w_12318),.q(n370));
  bfr _b_10693(.a(_w_12595),.q(_w_12596));
  bfr _b_10415(.a(_w_12317),.q(_w_12318));
  bfr _b_10413(.a(_w_12315),.q(_w_12316));
  bfr _b_14209(.a(_w_16111),.q(_w_16112));
  bfr _b_10412(.a(_w_12314),.q(_w_12315));
  bfr _b_10411(.a(_w_12313),.q(_w_12314));
  bfr _b_12336(.a(_w_14238),.q(_w_14239));
  bfr _b_10410(.a(_w_12312),.q(_w_12313));
  bfr _b_10409(.a(_w_12311),.q(_w_12312));
  bfr _b_10406(.a(_w_12308),.q(_w_12309));
  bfr _b_10405(.a(_w_12307),.q(_w_12308));
  bfr _b_10403(.a(_w_12305),.q(_w_12306));
  bfr _b_10401(.a(_w_12303),.q(_w_12304));
  bfr _b_12462(.a(_w_14364),.q(n1786));
  bfr _b_10400(.a(_w_12302),.q(_w_12303));
  bfr _b_10399(.a(_w_12301),.q(n978));
  bfr _b_10397(.a(_w_12299),.q(_w_12300));
  bfr _b_10394(.a(_w_12296),.q(n368));
  bfr _b_10392(.a(_w_12294),.q(_w_12295));
  bfr _b_10391(.a(_w_12293),.q(_w_12294));
  bfr _b_10390(.a(_w_12292),.q(_w_12293));
  bfr _b_10389(.a(_w_12291),.q(_w_12292));
  bfr _b_13656(.a(_w_15558),.q(_w_15559));
  bfr _b_10388(.a(_w_12290),.q(_w_12291));
  bfr _b_10387(.a(_w_12289),.q(_w_12290));
  bfr _b_10385(.a(_w_12287),.q(_w_12288));
  bfr _b_13903(.a(_w_15805),.q(_w_15806));
  bfr _b_10384(.a(_w_12286),.q(_w_12287));
  bfr _b_10382(.a(_w_12284),.q(_w_12285));
  bfr _b_10380(.a(_w_12282),.q(_w_12283));
  bfr _b_10378(.a(_w_12280),.q(n524));
  bfr _b_13307(.a(_w_15209),.q(_w_15210));
  bfr _b_10377(.a(_w_12279),.q(_w_12280));
  bfr _b_12733(.a(_w_14635),.q(_w_14636));
  bfr _b_10609(.a(_w_12511),.q(n1464));
  bfr _b_10375(.a(_w_12277),.q(_w_12278));
  bfr _b_10374(.a(_w_12276),.q(N6200));
  bfr _b_10373(.a(_w_12275),.q(_w_12276));
  bfr _b_10372(.a(_w_12274),.q(_w_12275));
  bfr _b_12015(.a(_w_13917),.q(_w_13918));
  bfr _b_10371(.a(_w_12273),.q(_w_12274));
  bfr _b_10370(.a(_w_12272),.q(_w_12273));
  bfr _b_10368(.a(_w_12270),.q(_w_12271));
  bfr _b_10367(.a(_w_12269),.q(_w_12270));
  bfr _b_10366(.a(_w_12268),.q(_w_12269));
  bfr _b_10360(.a(_w_12262),.q(_w_12263));
  bfr _b_10359(.a(_w_12261),.q(_w_12262));
  bfr _b_10356(.a(_w_12258),.q(_w_12259));
  bfr _b_10355(.a(_w_12257),.q(_w_12258));
  bfr _b_10354(.a(_w_12256),.q(_w_12257));
  bfr _b_10353(.a(_w_12255),.q(_w_12256));
  bfr _b_10350(.a(_w_12252),.q(_w_12253));
  bfr _b_13606(.a(_w_15508),.q(N18_14));
  bfr _b_10347(.a(_w_12249),.q(_w_12250));
  bfr _b_12269(.a(_w_14171),.q(_w_14172));
  bfr _b_10346(.a(_w_12248),.q(_w_12249));
  bfr _b_10341(.a(_w_12243),.q(_w_12244));
  bfr _b_10339(.a(_w_12241),.q(_w_12242));
  bfr _b_10337(.a(_w_12239),.q(_w_12240));
  bfr _b_10336(.a(_w_12238),.q(_w_12239));
  bfr _b_10335(.a(_w_12237),.q(_w_12238));
  bfr _b_10332(.a(_w_12234),.q(_w_12235));
  bfr _b_10330(.a(_w_12232),.q(_w_12233));
  bfr _b_14088(.a(_w_15990),.q(_w_15991));
  bfr _b_10327(.a(_w_12229),.q(_w_12230));
  bfr _b_10326(.a(_w_12228),.q(_w_12229));
  bfr _b_10325(.a(_w_12227),.q(_w_12228));
  bfr _b_10323(.a(_w_12225),.q(_w_12226));
  bfr _b_10322(.a(_w_12224),.q(_w_12225));
  bfr _b_10320(.a(_w_12222),.q(_w_12223));
  bfr _b_10318(.a(_w_12220),.q(_w_12221));
  bfr _b_10316(.a(_w_12218),.q(_w_12219));
  bfr _b_14375(.a(_w_16277),.q(_w_16278));
  bfr _b_14312(.a(_w_16214),.q(_w_16215));
  bfr _b_10314(.a(_w_12216),.q(n1396));
  bfr _b_10313(.a(_w_12215),.q(n1004_1));
  bfr _b_10312(.a(_w_12214),.q(_w_12215));
  bfr _b_10310(.a(_w_12212),.q(_w_12213));
  bfr _b_10308(.a(_w_12210),.q(n354_1));
  bfr _b_10307(.a(_w_12209),.q(_w_12210));
  bfr _b_11415(.a(_w_13317),.q(_w_13318));
  bfr _b_10306(.a(_w_12208),.q(_w_12209));
  bfr _b_10305(.a(_w_12207),.q(_w_12208));
  bfr _b_10303(.a(_w_12205),.q(N4241));
  bfr _b_10302(.a(_w_12204),.q(_w_12205));
  bfr _b_13687(.a(_w_15589),.q(_w_15590));
  bfr _b_10728(.a(_w_12630),.q(_w_12631));
  bfr _b_10299(.a(_w_12201),.q(_w_12202));
  bfr _b_10298(.a(_w_12200),.q(_w_12201));
  bfr _b_10296(.a(_w_12198),.q(_w_12199));
  bfr _b_10293(.a(_w_12195),.q(_w_12196));
  bfr _b_10292(.a(_w_12194),.q(_w_12195));
  bfr _b_10290(.a(_w_12192),.q(_w_12193));
  bfr _b_10289(.a(_w_12191),.q(_w_12192));
  bfr _b_10288(.a(_w_12190),.q(_w_12191));
  bfr _b_10286(.a(_w_12188),.q(_w_12189));
  bfr _b_10284(.a(_w_12186),.q(_w_12187));
  bfr _b_10283(.a(_w_12185),.q(_w_12186));
  bfr _b_11310(.a(_w_13212),.q(_w_13213));
  bfr _b_10282(.a(_w_12184),.q(_w_12185));
  bfr _b_10281(.a(_w_12183),.q(_w_12184));
  bfr _b_10280(.a(_w_12182),.q(_w_12183));
  bfr _b_10279(.a(_w_12181),.q(_w_12182));
  bfr _b_10278(.a(_w_12180),.q(_w_12181));
  bfr _b_10277(.a(_w_12179),.q(_w_12180));
  bfr _b_10275(.a(_w_12177),.q(_w_12178));
  bfr _b_10274(.a(_w_12176),.q(_w_12177));
  bfr _b_5086(.a(_w_6988),.q(_w_6989));
  bfr _b_8624(.a(_w_10526),.q(_w_10527));
  bfr _b_5079(.a(_w_6981),.q(_w_6982));
  bfr _b_9071(.a(_w_10973),.q(_w_10974));
  bfr _b_5078(.a(_w_6980),.q(_w_6981));
  bfr _b_9116(.a(_w_11018),.q(_w_11019));
  bfr _b_3640(.a(_w_5542),.q(n1698_1));
  bfr _b_8836(.a(_w_10738),.q(_w_10739));
  bfr _b_5069(.a(_w_6971),.q(_w_6972));
  bfr _b_5064(.a(_w_6966),.q(_w_6967));
  bfr _b_5059(.a(_w_6961),.q(_w_6962));
  bfr _b_5057(.a(_w_6959),.q(_w_6960));
  bfr _b_5055(.a(_w_6957),.q(_w_6958));
  bfr _b_6340(.a(_w_8242),.q(_w_8243));
  bfr _b_5041(.a(_w_6943),.q(_w_6944));
  bfr _b_8789(.a(_w_10691),.q(_w_10692));
  bfr _b_5080(.a(_w_6982),.q(_w_6983));
  spl4L N205_s_1(.a(N205_0),.q0(N205_4),.q1(N205_5),.q2(_w_8020),.q3(_w_8022));
  bfr _b_5035(.a(_w_6937),.q(_w_6938));
  bfr _b_5073(.a(_w_6975),.q(_w_6976));
  bfr _b_5032(.a(_w_6934),.q(_w_6935));
  spl4L N154_s_4(.a(N154_3),.q0(N154_16),.q1(N154_17),.q2(N154_18),.q3(N154_19));
  bfr _b_9699(.a(_w_11601),.q(n434));
  bfr _b_5011(.a(_w_6913),.q(_w_6914));
  bfr _b_6563(.a(_w_8465),.q(_w_8466));
  bfr _b_5003(.a(_w_6905),.q(_w_6906));
  bfr _b_5000(.a(_w_6902),.q(_w_6903));
  bfr _b_13832(.a(_w_15734),.q(_w_15735));
  and_bi g804(.a(n802_0),.b(n803),.q(n804));
  bfr _b_6920(.a(_w_8822),.q(_w_8823));
  bfr _b_4991(.a(_w_6893),.q(_w_6894));
  bfr _b_4990(.a(_w_6892),.q(_w_6893));
  and_bi g420(.a(n418_0),.b(n419),.q(n420));
  bfr _b_4987(.a(_w_6889),.q(_w_6890));
  bfr _b_4983(.a(_w_6885),.q(N103_7));
  bfr _b_4978(.a(_w_6880),.q(_w_6881));
  spl2 g1517_s_0(.a(n1517),.q0(n1517_0),.q1(n1517_1));
  and_bi g1607(.a(n1594_1),.b(n1597_1),.q(n1607));
  bfr _b_4977(.a(_w_6879),.q(_w_6880));
  bfr _b_4976(.a(_w_6878),.q(_w_6879));
  bfr _b_4974(.a(_w_6876),.q(_w_6877));
  bfr _b_12417(.a(_w_14319),.q(_w_14320));
  bfr _b_4972(.a(_w_6874),.q(_w_6875));
  bfr _b_4971(.a(_w_6873),.q(_w_6874));
  bfr _b_12810(.a(_w_14712),.q(_w_14713));
  spl2 g1879_s_0(.a(n1879),.q0(n1879_0),.q1(n1879_1));
  bfr _b_4968(.a(_w_6870),.q(_w_6871));
  bfr _b_4967(.a(_w_6869),.q(_w_6870));
  bfr _b_4961(.a(_w_6863),.q(_w_6864));
  bfr _b_12346(.a(_w_14248),.q(_w_14249));
  bfr _b_5306(.a(_w_7208),.q(_w_7209));
  bfr _b_5484(.a(_w_7386),.q(_w_7387));
  bfr _b_9362(.a(_w_11264),.q(_w_11265));
  bfr _b_10176(.a(_w_12078),.q(n809));
  bfr _b_4958(.a(_w_6860),.q(_w_6861));
  bfr _b_4956(.a(_w_6858),.q(_w_6859));
  bfr _b_10285(.a(_w_12187),.q(_w_12188));
  spl2 g622_s_0(.a(n622),.q0(n622_0),.q1(n622_1));
  bfr _b_5287(.a(_w_7189),.q(_w_7190));
  bfr _b_4952(.a(_w_6854),.q(_w_6855));
  bfr _b_4948(.a(_w_6850),.q(_w_6851));
  and_bi g392(.a(n374_1),.b(n390_1),.q(_w_11598));
  bfr _b_4946(.a(_w_6848),.q(_w_6849));
  bfr _b_7317(.a(_w_9219),.q(n647));
  bfr _b_4943(.a(_w_6845),.q(_w_6846));
  bfr _b_11483(.a(_w_13385),.q(_w_13386));
  bfr _b_4942(.a(_w_6844),.q(_w_6845));
  bfr _b_4941(.a(_w_6843),.q(_w_6844));
  bfr _b_4936(.a(_w_6838),.q(_w_6839));
  bfr _b_4250(.a(_w_6152),.q(N171_7));
  bfr _b_6442(.a(_w_8344),.q(_w_8345));
  spl2 g545_s_0(.a(n545),.q0(n545_0),.q1(n545_1));
  bfr _b_4933(.a(_w_6835),.q(_w_6836));
  bfr _b_12288(.a(_w_14190),.q(_w_14191));
  spl2 g753_s_0(.a(n753),.q0(n753_0),.q1(n753_1));
  bfr _b_8579(.a(_w_10481),.q(_w_10482));
  and_bi g854(.a(n853_0),.b(n846_0),.q(n854));
  bfr _b_10333(.a(_w_12235),.q(_w_12236));
  bfr _b_5034(.a(_w_6936),.q(_w_6937));
  bfr _b_5774(.a(_w_7676),.q(_w_7677));
  bfr _b_4927(.a(_w_6829),.q(_w_6830));
  bfr _b_4924(.a(_w_6826),.q(_w_6827));
  bfr _b_8474(.a(_w_10376),.q(_w_10377));
  bfr _b_4917(.a(_w_6819),.q(_w_6820));
  bfr _b_4912(.a(_w_6814),.q(_w_6815));
  bfr _b_10472(.a(_w_12374),.q(_w_12375));
  and_bb g308(.a(n247_1),.b(n307_0),.q(n308));
  bfr _b_4981(.a(_w_6883),.q(N103_6));
  bfr _b_8604(.a(_w_10506),.q(_w_10507));
  bfr _b_4911(.a(_w_6813),.q(_w_6814));
  bfr _b_4910(.a(_w_6812),.q(_w_6813));
  bfr _b_14081(.a(_w_15983),.q(_w_15984));
  bfr _b_4905(.a(_w_6807),.q(_w_6808));
  bfr _b_9795(.a(_w_11697),.q(_w_11698));
  bfr _b_4893(.a(_w_6795),.q(_w_6796));
  bfr _b_4887(.a(_w_6789),.q(N137_2));
  and_bb g144(.a(N307_8),.b(N69_6),.q(_w_9623));
  bfr _b_4886(.a(_w_6788),.q(_w_6789));
  bfr _b_13601(.a(_w_15503),.q(_w_15504));
  bfr _b_7180(.a(_w_9082),.q(_w_9083));
  bfr _b_13894(.a(_w_15796),.q(_w_15797));
  bfr _b_8963(.a(_w_10865),.q(_w_10866));
  bfr _b_6832(.a(_w_8734),.q(_w_8735));
  bfr _b_4883(.a(_w_6785),.q(_w_6786));
  and_bi g64(.a(n54_1),.b(n62_1),.q(_w_8564));
  bfr _b_10417(.a(_w_12319),.q(_w_12320));
  bfr _b_6647(.a(_w_8549),.q(_w_8550));
  bfr _b_4876(.a(_w_6778),.q(_w_6779));
  spl2 g1799_s_0(.a(n1799),.q0(n1799_0),.q1(n1799_1));
  bfr _b_6016(.a(_w_7918),.q(_w_7919));
  bfr _b_10936(.a(_w_12838),.q(n718));
  bfr _b_10376(.a(_w_12278),.q(_w_12279));
  bfr _b_4874(.a(_w_6776),.q(_w_6777));
  bfr _b_12117(.a(_w_14019),.q(_w_14020));
  spl2 g1194_s_0(.a(n1194),.q0(n1194_0),.q1(_w_6181));
  bfr _b_11911(.a(_w_13813),.q(_w_13814));
  bfr _b_9485(.a(_w_11387),.q(_w_11388));
  bfr _b_4873(.a(_w_6775),.q(_w_6776));
  bfr _b_11302(.a(_w_13204),.q(n1135));
  bfr _b_4870(.a(_w_6772),.q(_w_6773));
  bfr _b_11800(.a(_w_13702),.q(_w_13703));
  and_bi g914(.a(n913_0),.b(n826_0),.q(n914));
  bfr _b_4868(.a(_w_6770),.q(_w_6771));
  bfr _b_8459(.a(_w_10361),.q(_w_10362));
  bfr _b_6281(.a(_w_8183),.q(_w_8184));
  bfr _b_4861(.a(_w_6763),.q(_w_6764));
  spl2 g1448_s_0(.a(n1448),.q0(n1448_0),.q1(n1448_1));
  bfr _b_4858(.a(_w_6760),.q(_w_6761));
  bfr _b_4303(.a(_w_6205),.q(_w_6206));
  bfr _b_4856(.a(_w_6758),.q(_w_6759));
  bfr _b_4853(.a(_w_6755),.q(_w_6756));
  bfr _b_4847(.a(_w_6749),.q(_w_6750));
  spl2 g693_s_0(.a(n693),.q0(n693_0),.q1(n693_1));
  and_bb g232(.a(N1_12),.b(N409_4),.q(n232));
  bfr _b_14177(.a(_w_16079),.q(_w_16080));
  bfr _b_4841(.a(_w_6743),.q(_w_6744));
  bfr _b_7366(.a(_w_9268),.q(_w_9269));
  bfr _b_4838(.a(_w_6740),.q(_w_6741));
  bfr _b_4837(.a(_w_6739),.q(_w_6740));
  bfr _b_5017(.a(_w_6919),.q(_w_6920));
  bfr _b_10121(.a(_w_12023),.q(_w_12024));
  bfr _b_14365(.a(_w_16267),.q(_w_16268));
  bfr _b_4835(.a(_w_6737),.q(_w_6738));
  bfr _b_7351(.a(_w_9253),.q(_w_9254));
  bfr _b_7398(.a(_w_9300),.q(_w_9301));
  bfr _b_4871(.a(_w_6773),.q(_w_6774));
  or_bb g1600(.a(n1534_0),.b(n1599_0),.q(_w_12980));
  bfr _b_4834(.a(_w_6736),.q(_w_6737));
  bfr _b_4833(.a(_w_6735),.q(_w_6736));
  bfr _b_8307(.a(_w_10209),.q(_w_10210));
  bfr _b_10453(.a(_w_12355),.q(n1192));
  bfr _b_4832(.a(_w_6734),.q(_w_6735));
  bfr _b_4285(.a(_w_6187),.q(n738_1));
  and_bi g837(.a(n766_1),.b(n769_1),.q(n837));
  bfr _b_5047(.a(_w_6949),.q(_w_6950));
  bfr _b_10800(.a(_w_12702),.q(_w_12703));
  bfr _b_9518(.a(_w_11420),.q(_w_11421));
  bfr _b_4826(.a(_w_6728),.q(_w_6729));
  bfr _b_5001(.a(_w_6903),.q(_w_6904));
  bfr _b_4824(.a(_w_6726),.q(_w_6727));
  bfr _b_4818(.a(_w_6720),.q(_w_6721));
  bfr _b_14305(.a(_w_16207),.q(_w_16208));
  bfr _b_6846(.a(_w_8748),.q(n1047));
  bfr _b_4814(.a(_w_6716),.q(_w_6717));
  spl2 g1612_s_0(.a(n1612),.q0(n1612_0),.q1(n1612_1));
  bfr _b_12640(.a(_w_14542),.q(_w_14543));
  bfr _b_11426(.a(_w_13328),.q(_w_13329));
  bfr _b_4811(.a(_w_6713),.q(_w_6714));
  bfr _b_4830(.a(_w_6732),.q(_w_6733));
  bfr _b_5023(.a(_w_6925),.q(_w_6926));
  bfr _b_4807(.a(_w_6709),.q(n1303_1));
  bfr _b_5522(.a(_w_7424),.q(_w_7425));
  or_bb g1433(.a(n1431_0),.b(n1432),.q(n1433));
  bfr _b_6233(.a(_w_8135),.q(_w_8136));
  bfr _b_4801(.a(_w_6703),.q(_w_6704));
  bfr _b_4800(.a(_w_6702),.q(_w_6703));
  bfr _b_7304(.a(_w_9206),.q(_w_9207));
  bfr _b_4799(.a(_w_6701),.q(n1224_1));
  bfr _b_11087(.a(_w_12989),.q(_w_12990));
  spl2 g1061_s_0(.a(n1061),.q0(n1061_0),.q1(n1061_1));
  bfr _b_4793(.a(_w_6695),.q(n192_1));
  bfr _b_13646(.a(_w_15548),.q(_w_15549));
  bfr _b_4790(.a(_w_6692),.q(_w_6693));
  bfr _b_6021(.a(_w_7923),.q(_w_7924));
  bfr _b_4787(.a(_w_6689),.q(N1_11));
  bfr _b_12249(.a(_w_14151),.q(n1723));
  bfr _b_4783(.a(_w_6685),.q(_w_6686));
  bfr _b_4778(.a(_w_6680),.q(_w_6681));
  bfr _b_4775(.a(_w_6677),.q(_w_6678));
  bfr _b_9590(.a(_w_11492),.q(_w_11493));
  bfr _b_4774(.a(_w_6676),.q(_w_6677));
  bfr _b_12144(.a(_w_14046),.q(_w_14047));
  bfr _b_11165(.a(_w_13067),.q(_w_13068));
  bfr _b_4497(.a(_w_6399),.q(_w_6400));
  bfr _b_4769(.a(_w_6671),.q(_w_6672));
  bfr _b_4768(.a(_w_6670),.q(_w_6671));
  bfr _b_4959(.a(_w_6861),.q(_w_6862));
  bfr _b_13846(.a(_w_15748),.q(_w_15749));
  bfr _b_4581(.a(_w_6483),.q(_w_6484));
  bfr _b_6780(.a(_w_8682),.q(_w_8683));
  bfr _b_4757(.a(_w_6659),.q(_w_6660));
  or_bb g784(.a(n723_0),.b(n783_0),.q(n784));
  bfr _b_5920(.a(_w_7822),.q(_w_7823));
  bfr _b_4753(.a(_w_6655),.q(_w_6656));
  bfr _b_4744(.a(_w_6646),.q(_w_6647));
  or_bb g675(.a(n673_0),.b(n674),.q(n675));
  bfr _b_4742(.a(_w_6644),.q(_w_6645));
  bfr _b_8400(.a(_w_10302),.q(_w_10303));
  bfr _b_4740(.a(_w_6642),.q(_w_6643));
  bfr _b_4738(.a(_w_6640),.q(_w_6641));
  and_bb g936(.a(N18_19),.b(N528_5),.q(_w_8595));
  bfr _b_5221(.a(_w_7123),.q(_w_7124));
  bfr _b_4736(.a(_w_6638),.q(_w_6639));
  bfr _b_4732(.a(_w_6634),.q(_w_6635));
  bfr _b_12447(.a(_w_14349),.q(_w_14350));
  and_bb g377(.a(N171_4),.b(N290_14),.q(n377));
  bfr _b_4730(.a(_w_6632),.q(_w_6633));
  bfr _b_12018(.a(_w_13920),.q(_w_13921));
  and_bi g692(.a(n618_1),.b(n690_1),.q(_w_9220));
  bfr _b_4722(.a(_w_6624),.q(_w_6625));
  bfr _b_12320(.a(_w_14222),.q(_w_14223));
  bfr _b_11381(.a(_w_13283),.q(_w_13284));
  bfr _b_4717(.a(_w_6619),.q(_w_6620));
  spl2 g177_s_0(.a(n177),.q0(n177_0),.q1(n177_1));
  bfr _b_4716(.a(_w_6618),.q(_w_6619));
  spl2 g1276_s_0(.a(n1276),.q0(n1276_0),.q1(n1276_1));
  bfr _b_5918(.a(_w_7820),.q(_w_7821));
  bfr _b_12468(.a(_w_14370),.q(_w_14371));
  and_bi g1087(.a(n1072_1),.b(n1085_1),.q(_w_8389));
  bfr _b_4712(.a(_w_6614),.q(_w_6615));
  bfr _b_12406(.a(_w_14308),.q(_w_14309));
  spl2 g842_s_0(.a(n842),.q0(n842_0),.q1(n842_1));
  bfr _b_11840(.a(_w_13742),.q(_w_13743));
  and_bi g1606(.a(n1600_1),.b(n1603_1),.q(n1606));
  bfr _b_5809(.a(_w_7711),.q(_w_7712));
  bfr _b_4706(.a(_w_6608),.q(_w_6609));
  bfr _b_12999(.a(_w_14901),.q(_w_14902));
  bfr _b_4702(.a(_w_6604),.q(_w_6605));
  bfr _b_4700(.a(_w_6602),.q(_w_6603));
  spl2 g241_s_0(.a(n241),.q0(n241_0),.q1(n241_1));
  bfr _b_4696(.a(_w_6598),.q(_w_6599));
  bfr _b_4888(.a(_w_6790),.q(_w_6791));
  bfr _b_5031(.a(_w_6933),.q(_w_6934));
  bfr _b_4690(.a(_w_6592),.q(_w_6593));
  bfr _b_14139(.a(_w_16041),.q(_w_16042));
  bfr _b_4689(.a(_w_6591),.q(_w_6592));
  bfr _b_6894(.a(_w_8796),.q(_w_8797));
  bfr _b_4683(.a(_w_6585),.q(_w_6586));
  bfr _b_4681(.a(_w_6583),.q(_w_6584));
  bfr _b_11528(.a(_w_13430),.q(n1295));
  bfr _b_6487(.a(_w_8389),.q(n1087));
  bfr _b_4680(.a(_w_6582),.q(_w_6583));
  bfr _b_4851(.a(_w_6753),.q(_w_6754));
  bfr _b_4676(.a(_w_6578),.q(_w_6579));
  bfr _b_13965(.a(_w_15867),.q(_w_15868));
  bfr _b_11769(.a(_w_13671),.q(_w_13672));
  bfr _b_5452(.a(_w_7354),.q(_w_7355));
  bfr _b_9667(.a(_w_11569),.q(_w_11570));
  bfr _b_4686(.a(_w_6588),.q(_w_6589));
  spl2 g1463_s_0(.a(n1463),.q0(n1463_0),.q1(n1463_1));
  bfr _b_4660(.a(_w_6562),.q(_w_6563));
  and_bi g865(.a(n863_0),.b(n864),.q(n865));
  bfr _b_4016(.a(_w_5918),.q(_w_5919));
  bfr _b_7346(.a(_w_9248),.q(n677));
  bfr _b_4658(.a(_w_6560),.q(_w_6561));
  bfr _b_7248(.a(_w_9150),.q(_w_9151));
  bfr _b_4655(.a(_w_6557),.q(_w_6558));
  or_bb g1149(.a(n1051_0),.b(n1148_0),.q(n1149));
  bfr _b_9278(.a(_w_11180),.q(_w_11181));
  bfr _b_13418(.a(_w_15320),.q(_w_15321));
  bfr _b_4650(.a(_w_6552),.q(_w_6553));
  bfr _b_12655(.a(_w_14557),.q(_w_14558));
  or_bb g1833(.a(n1823_0),.b(n1832_0),.q(n1833));
  or_bb g329(.a(n327_0),.b(n328),.q(n329));
  bfr _b_12384(.a(_w_14286),.q(_w_14287));
  spl2 g127_s_0(.a(n127),.q0(n127_0),.q1(n127_1));
  spl2 g1899_s_0(.a(n1899),.q0(n1899_0),.q1(n1899_1));
  bfr _b_6029(.a(_w_7931),.q(_w_7932));
  bfr _b_11780(.a(_w_13682),.q(_w_13683));
  bfr _b_9720(.a(_w_11622),.q(_w_11623));
  bfr _b_8248(.a(_w_10150),.q(_w_10151));
  bfr _b_9969(.a(_w_11871),.q(_w_11872));
  bfr _b_4642(.a(_w_6544),.q(_w_6545));
  spl2 g90_s_0(.a(n90),.q0(n90_0),.q1(n90_1));
  bfr _b_13093(.a(_w_14995),.q(_w_14996));
  bfr _b_12805(.a(_w_14707),.q(_w_14708));
  bfr _b_5924(.a(_w_7826),.q(_w_7827));
  bfr _b_9755(.a(_w_11657),.q(_w_11658));
  bfr _b_4639(.a(_w_6541),.q(_w_6542));
  bfr _b_4637(.a(_w_6539),.q(_w_6540));
  bfr _b_3858(.a(_w_5760),.q(_w_5761));
  bfr _b_14106(.a(_w_16008),.q(_w_16009));
  bfr _b_12146(.a(_w_14048),.q(_w_14049));
  bfr _b_4636(.a(_w_6538),.q(_w_6539));
  spl2 g1476_s_0(.a(n1476),.q0(n1476_0),.q1(n1476_1));
  bfr _b_7378(.a(_w_9280),.q(_w_9281));
  bfr _b_4635(.a(_w_6537),.q(_w_6538));
  bfr _b_5160(.a(_w_7062),.q(_w_7063));
  bfr _b_4634(.a(_w_6536),.q(_w_6537));
  bfr _b_12216(.a(_w_14118),.q(_w_14119));
  bfr _b_4630(.a(_w_6532),.q(_w_6533));
  bfr _b_12271(.a(_w_14173),.q(_w_14174));
  bfr _b_4629(.a(_w_6531),.q(_w_6532));
  bfr _b_4627(.a(_w_6529),.q(_w_6530));
  bfr _b_4623(.a(_w_6525),.q(_w_6526));
  bfr _b_9633(.a(_w_11535),.q(_w_11536));
  bfr _b_9957(.a(_w_11859),.q(_w_11860));
  bfr _b_4621(.a(_w_6523),.q(_w_6524));
  or_bb g1727(.a(n1725_0),.b(n1726),.q(_w_8155));
  bfr _b_11367(.a(_w_13269),.q(_w_13270));
  bfr _b_4619(.a(_w_6521),.q(_w_6522));
  bfr _b_3741(.a(_w_5643),.q(_w_5644));
  bfr _b_5213(.a(_w_7115),.q(_w_7116));
  bfr _b_4784(.a(_w_6686),.q(_w_6687));
  or_bb g1558(.a(n1548_0),.b(n1557_0),.q(n1558));
  bfr _b_6341(.a(_w_8243),.q(_w_8244));
  bfr _b_5076(.a(_w_6978),.q(_w_6979));
  bfr _b_8113(.a(_w_10015),.q(_w_10016));
  bfr _b_14340(.a(_w_16242),.q(_w_16243));
  bfr _b_4613(.a(_w_6515),.q(_w_6516));
  bfr _b_6842(.a(_w_8744),.q(_w_8745));
  bfr _b_4607(.a(_w_6509),.q(_w_6510));
  spl2 g1060_s_0(.a(n1060),.q0(n1060_0),.q1(n1060_1));
  bfr _b_4731(.a(_w_6633),.q(N154_3));
  and_bi g1735(.a(n1698_1),.b(n1701_1),.q(n1735));
  bfr _b_11871(.a(_w_13773),.q(_w_13774));
  bfr _b_4602(.a(_w_6504),.q(_w_6505));
  bfr _b_4973(.a(_w_6875),.q(_w_6876));
  bfr _b_4599(.a(_w_6501),.q(_w_6502));
  bfr _b_11100(.a(_w_13002),.q(n1210));
  bfr _b_4588(.a(_w_6490),.q(_w_6491));
  bfr _b_5170(.a(_w_7072),.q(_w_7073));
  bfr _b_10588(.a(_w_12490),.q(n251));
  bfr _b_4572(.a(_w_6474),.q(_w_6475));
  bfr _b_4568(.a(_w_6470),.q(_w_6471));
  bfr _b_4567(.a(_w_6469),.q(_w_6470));
  bfr _b_4565(.a(_w_6467),.q(_w_6468));
  bfr _b_4552(.a(_w_6454),.q(_w_6455));
  bfr _b_10895(.a(_w_12797),.q(_w_12798));
  bfr _b_4955(.a(_w_6857),.q(_w_6858));
  bfr _b_4538(.a(_w_6440),.q(_w_6441));
  bfr _b_4563(.a(_w_6465),.q(N154_7));
  bfr _b_4533(.a(_w_6435),.q(_w_6436));
  bfr _b_11955(.a(_w_13857),.q(n1492));
  and_bb g722(.a(N426_9),.b(N86_13),.q(n722));
  and_bi g1823(.a(n1794_1),.b(n1797_1),.q(n1823));
  bfr _b_9964(.a(_w_11866),.q(_w_11867));
  bfr _b_4530(.a(_w_6432),.q(_w_6433));
  bfr _b_3676(.a(_w_5578),.q(_w_5579));
  bfr _b_4528(.a(_w_6430),.q(_w_6431));
  bfr _b_8875(.a(_w_10777),.q(N3895));
  bfr _b_13900(.a(_w_15802),.q(_w_15803));
  bfr _b_11803(.a(_w_13705),.q(_w_13706));
  bfr _b_4656(.a(_w_6558),.q(_w_6559));
  bfr _b_11882(.a(_w_13784),.q(_w_13785));
  bfr _b_5911(.a(_w_7813),.q(_w_7814));
  bfr _b_5273(.a(_w_7175),.q(_w_7176));
  bfr _b_14085(.a(_w_15987),.q(_w_15988));
  bfr _b_4523(.a(_w_6425),.q(N137_15));
  bfr _b_6662(.a(_w_8564),.q(n64));
  bfr _b_4522(.a(_w_6424),.q(_w_6425));
  bfr _b_11035(.a(_w_12937),.q(n1167));
  bfr _b_4521(.a(_w_6423),.q(_w_6424));
  and_bi g533(.a(n478_1),.b(n481_1),.q(n533));
  bfr _b_10918(.a(_w_12820),.q(_w_12821));
  bfr _b_8554(.a(_w_10456),.q(_w_10457));
  bfr _b_4517(.a(_w_6419),.q(_w_6420));
  bfr _b_3421(.a(_w_5323),.q(_w_5324));
  bfr _b_4511(.a(_w_6413),.q(N137_14));
  bfr _b_4638(.a(_w_6540),.q(_w_6541));
  bfr _b_6433(.a(_w_8335),.q(_w_8336));
  bfr _b_4507(.a(_w_6409),.q(_w_6410));
  bfr _b_4506(.a(_w_6408),.q(_w_6409));
  bfr _b_4505(.a(_w_6407),.q(_w_6408));
  bfr _b_4501(.a(_w_6403),.q(_w_6404));
  bfr _b_4012(.a(_w_5914),.q(_w_5915));
  bfr _b_4499(.a(_w_6401),.q(N137_13));
  bfr _b_4498(.a(_w_6400),.q(_w_6401));
  bfr _b_4496(.a(_w_6398),.q(_w_6399));
  spl2 g1052_s_0(.a(n1052),.q0(n1052_0),.q1(n1052_1));
  bfr _b_12749(.a(_w_14651),.q(_w_14652));
  bfr _b_4494(.a(_w_6396),.q(_w_6397));
  bfr _b_10441(.a(_w_12343),.q(_w_12344));
  bfr _b_6269(.a(_w_8171),.q(_w_8172));
  bfr _b_4601(.a(_w_6503),.q(_w_6504));
  bfr _b_6136(.a(_w_8038),.q(_w_8039));
  bfr _b_4492(.a(_w_6394),.q(_w_6395));
  bfr _b_4491(.a(_w_6393),.q(n256_1));
  bfr _b_4482(.a(_w_6384),.q(_w_6385));
  bfr _b_4477(.a(_w_6379),.q(n42_1));
  bfr _b_5450(.a(_w_7352),.q(_w_7353));
  bfr _b_11479(.a(_w_13381),.q(_w_13382));
  bfr _b_4473(.a(_w_6375),.q(_w_6376));
  bfr _b_12871(.a(_w_14773),.q(_w_14774));
  and_bi g49(.a(n48_0),.b(n40_0),.q(n49));
  bfr _b_10393(.a(_w_12295),.q(_w_12296));
  bfr _b_4468(.a(_w_6370),.q(_w_6371));
  bfr _b_4466(.a(_w_6368),.q(_w_6369));
  bfr _b_11062(.a(_w_12964),.q(_w_12965));
  and_bb g718(.a(N460_7),.b(N52_15),.q(_w_12827));
  bfr _b_5877(.a(_w_7779),.q(_w_7780));
  bfr _b_4463(.a(_w_6365),.q(n168_1));
  bfr _b_7735(.a(_w_9637),.q(n589));
  bfr _b_4462(.a(_w_6364),.q(_w_6365));
  spl2 g963_s_0(.a(n963),.q0(n963_0),.q1(n963_1));
  bfr _b_12020(.a(_w_13922),.q(n1537));
  bfr _b_5242(.a(_w_7144),.q(_w_7145));
  bfr _b_4461(.a(_w_6363),.q(_w_6364));
  bfr _b_9772(.a(_w_11674),.q(_w_11675));
  bfr _b_4458(.a(_w_6360),.q(_w_6361));
  bfr _b_4457(.a(_w_6359),.q(_w_6360));
  bfr _b_8088(.a(_w_9990),.q(_w_9991));
  bfr _b_7060(.a(_w_8962),.q(_w_8963));
  bfr _b_4748(.a(_w_6650),.q(_w_6651));
  bfr _b_4483(.a(_w_6385),.q(n968_1));
  bfr _b_3749(.a(_w_5651),.q(_w_5652));
  bfr _b_4450(.a(_w_6352),.q(_w_6353));
  spl2 g1247_s_0(.a(n1247),.q0(n1247_0),.q1(n1247_1));
  bfr _b_4899(.a(_w_6801),.q(_w_6802));
  bfr _b_7623(.a(_w_9525),.q(_w_9526));
  spl2 g1312_s_0(.a(n1312),.q0(n1312_0),.q1(n1312_1));
  bfr _b_4445(.a(_w_6347),.q(_w_6348));
  bfr _b_13732(.a(_w_15634),.q(_w_15635));
  bfr _b_5539(.a(_w_7441),.q(_w_7442));
  bfr _b_4444(.a(_w_6346),.q(_w_6347));
  spl4L N460_s_1(.a(N460_0),.q0(N460_4),.q1(N460_5),.q2(N460_6),.q3(N460_7));
  spl4L N171_s_4(.a(N171_3),.q0(N171_16),.q1(N171_17),.q2(N171_18),.q3(N171_19));
  bfr _b_12692(.a(_w_14594),.q(_w_14595));
  bfr _b_4435(.a(_w_6337),.q(n162_1));
  bfr _b_4429(.a(_w_6331),.q(_w_6332));
  bfr _b_9722(.a(_w_11624),.q(_w_11625));
  bfr _b_11744(.a(_w_13646),.q(_w_13647));
  bfr _b_8529(.a(_w_10431),.q(_w_10432));
  bfr _b_4423(.a(_w_6325),.q(_w_6326));
  or_bb g1309(.a(n1283_0),.b(n1308_0),.q(n1309));
  bfr _b_4421(.a(_w_6323),.q(_w_6324));
  bfr _b_13980(.a(_w_15882),.q(_w_15883));
  bfr _b_13624(.a(N120),.q(_w_15526));
  bfr _b_5474(.a(_w_7376),.q(_w_7377));
  bfr _b_10661(.a(_w_12563),.q(_w_12564));
  bfr _b_8763(.a(_w_10665),.q(_w_10666));
  bfr _b_4685(.a(_w_6587),.q(_w_6588));
  bfr _b_4419(.a(_w_6321),.q(_w_6322));
  bfr _b_4409(.a(_w_6311),.q(_w_6312));
  bfr _b_7097(.a(_w_8999),.q(_w_9000));
  bfr _b_11916(.a(_w_13818),.q(_w_13819));
  bfr _b_9411(.a(_w_11313),.q(_w_11314));
  bfr _b_11701(.a(_w_13603),.q(_w_13604));
  bfr _b_4406(.a(_w_6308),.q(n606_1));
  bfr _b_4405(.a(_w_6307),.q(_w_6308));
  bfr _b_3631(.a(_w_5533),.q(_w_5534));
  bfr _b_4714(.a(_w_6616),.q(_w_6617));
  bfr _b_4139(.a(_w_6041),.q(_w_6042));
  bfr _b_3955(.a(_w_5857),.q(_w_5858));
  bfr _b_6032(.a(_w_7934),.q(_w_7935));
  bfr _b_4400(.a(_w_6302),.q(_w_6303));
  bfr _b_7913(.a(_w_9815),.q(_w_9816));
  bfr _b_11389(.a(_w_13291),.q(_w_13292));
  bfr _b_4398(.a(_w_6300),.q(_w_6301));
  bfr _b_4397(.a(_w_6299),.q(n1806_1));
  bfr _b_4395(.a(_w_6297),.q(_w_6298));
  bfr _b_4393(.a(_w_6295),.q(n582_1));
  bfr _b_12687(.a(_w_14589),.q(_w_14590));
  bfr _b_7702(.a(_w_9604),.q(_w_9605));
  bfr _b_4391(.a(_w_6293),.q(_w_6294));
  bfr _b_3613(.a(_w_5515),.q(_w_5516));
  bfr _b_4387(.a(_w_6289),.q(_w_6290));
  bfr _b_4386(.a(_w_6288),.q(_w_6289));
  bfr _b_4032(.a(_w_5934),.q(_w_5935));
  bfr _b_10779(.a(_w_12681),.q(_w_12682));
  bfr _b_4695(.a(_w_6597),.q(_w_6598));
  bfr _b_4375(.a(_w_6277),.q(_w_6278));
  bfr _b_10848(.a(_w_12750),.q(_w_12751));
  bfr _b_4372(.a(_w_6274),.q(_w_6275));
  bfr _b_10667(.a(_w_12569),.q(_w_12570));
  spl2 g853_s_0(.a(n853),.q0(n853_0),.q1(n853_1));
  bfr _b_7695(.a(_w_9597),.q(_w_9598));
  bfr _b_3709(.a(_w_5611),.q(_w_5612));
  bfr _b_4280(.a(_w_6182),.q(_w_6183));
  bfr _b_4356(.a(_w_6258),.q(_w_6259));
  bfr _b_4632(.a(_w_6534),.q(_w_6535));
  bfr _b_4432(.a(_w_6334),.q(_w_6335));
  bfr _b_4355(.a(_w_6257),.q(_w_6258));
  bfr _b_12115(.a(_w_14017),.q(_w_14018));
  bfr _b_4354(.a(_w_6256),.q(_w_6257));
  and_bb g612(.a(N1_17),.b(N494_4),.q(_w_11052));
  bfr _b_4353(.a(_w_6255),.q(_w_6256));
  bfr _b_4668(.a(_w_6570),.q(_w_6571));
  bfr _b_10250(.a(_w_12152),.q(_w_12153));
  bfr _b_4388(.a(_w_6290),.q(_w_6291));
  bfr _b_6644(.a(_w_8546),.q(_w_8547));
  bfr _b_8342(.a(_w_10244),.q(_w_10245));
  bfr _b_10237(.a(_w_12139),.q(_w_12140));
  bfr _b_4204(.a(_w_6106),.q(_w_6107));
  and_bb g695(.a(n617_1),.b(n693_1),.q(_w_11836));
  bfr _b_4345(.a(_w_6247),.q(_w_6248));
  bfr _b_7547(.a(_w_9449),.q(_w_9450));
  bfr _b_4344(.a(_w_6246),.q(_w_6247));
  bfr _b_4343(.a(_w_6245),.q(_w_6246));
  bfr _b_10802(.a(_w_12704),.q(_w_12705));
  bfr _b_4342(.a(_w_6244),.q(_w_6245));
  bfr _b_6752(.a(_w_8654),.q(_w_8655));
  bfr _b_9751(.a(_w_11653),.q(_w_11654));
  bfr _b_12286(.a(_w_14188),.q(_w_14189));
  bfr _b_4315(.a(_w_6217),.q(_w_6218));
  bfr _b_4340(.a(_w_6242),.q(_w_6243));
  bfr _b_3786(.a(_w_5688),.q(_w_5689));
  bfr _b_7185(.a(_w_9087),.q(_w_9088));
  bfr _b_4863(.a(_w_6765),.q(_w_6766));
  bfr _b_4339(.a(_w_6241),.q(_w_6242));
  bfr _b_6034(.a(_w_7936),.q(_w_7937));
  bfr _b_4336(.a(_w_6238),.q(_w_6239));
  spl2 g1224_s_0(.a(n1224),.q0(n1224_0),.q1(_w_6698));
  bfr _b_7589(.a(_w_9491),.q(_w_9492));
  bfr _b_4332(.a(_w_6234),.q(_w_6235));
  bfr _b_9170(.a(_w_11072),.q(_w_11073));
  bfr _b_4328(.a(_w_6230),.q(_w_6231));
  bfr _b_6972(.a(_w_8874),.q(_w_8875));
  bfr _b_11469(.a(_w_13371),.q(n212));
  bfr _b_4326(.a(_w_6228),.q(_w_6229));
  or_bb g646(.a(n633_0),.b(n645_0),.q(n646));
  bfr _b_10520(.a(_w_12422),.q(_w_12423));
  bfr _b_8962(.a(_w_10864),.q(_w_10865));
  bfr _b_12549(.a(_w_14451),.q(_w_14452));
  bfr _b_10605(.a(_w_12507),.q(n488));
  bfr _b_10223(.a(_w_12125),.q(_w_12126));
  bfr _b_13454(.a(_w_15356),.q(_w_15357));
  bfr _b_4323(.a(_w_6225),.q(_w_6226));
  bfr _b_4316(.a(_w_6218),.q(_w_6219));
  bfr _b_10683(.a(_w_12585),.q(_w_12586));
  bfr _b_4641(.a(_w_6543),.q(_w_6544));
  bfr _b_13976(.a(_w_15878),.q(_w_15879));
  and_bb g1456(.a(N120_18),.b(N511_11),.q(_w_10843));
  bfr _b_4554(.a(_w_6456),.q(_w_6457));
  bfr _b_4314(.a(_w_6216),.q(_w_6217));
  bfr _b_13114(.a(_w_15016),.q(_w_15017));
  bfr _b_4688(.a(_w_6590),.q(_w_6591));
  bfr _b_3586(.a(_w_5488),.q(_w_5489));
  spl2 g354_s_0(.a(n354),.q0(n354_0),.q1(_w_12207));
  and_bi g403(.a(n402_0),.b(n370_0),.q(n403));
  bfr _b_4311(.a(_w_6213),.q(_w_6214));
  or_bb g898(.a(n896_0),.b(n897),.q(n898));
  bfr _b_6570(.a(_w_8472),.q(_w_8473));
  bfr _b_6818(.a(_w_8720),.q(_w_8721));
  bfr _b_4913(.a(_w_6815),.q(_w_6816));
  bfr _b_4305(.a(_w_6207),.q(n670_1));
  bfr _b_6930(.a(_w_8832),.q(n820));
  bfr _b_14115(.a(_w_16017),.q(_w_16018));
  bfr _b_11656(.a(_w_13558),.q(_w_13559));
  bfr _b_8925(.a(_w_10827),.q(_w_10828));
  bfr _b_4304(.a(_w_6206),.q(_w_6207));
  bfr _b_11793(.a(_w_13695),.q(_w_13696));
  bfr _b_3836(.a(_w_5738),.q(_w_5739));
  bfr _b_11068(.a(_w_12970),.q(_w_12971));
  spl4L N358_s_3(.a(N358_2),.q0(N358_12),.q1(N358_13),.q2(N358_14),.q3(N358_15));
  bfr _b_6901(.a(_w_8803),.q(_w_8804));
  bfr _b_10924(.a(_w_12826),.q(n876));
  and_bb g543(.a(N205_5),.b(N273_16),.q(n543));
  bfr _b_9336(.a(_w_11238),.q(_w_11239));
  bfr _b_4301(.a(_w_6203),.q(n676_1));
  or_bb g997(.a(n995_0),.b(n996),.q(n997));
  spl2 g1368_s_0(.a(n1368),.q0(n1368_0),.q1(n1368_1));
  bfr _b_4294(.a(_w_6196),.q(_w_6197));
  bfr _b_14183(.a(_w_16085),.q(_w_16086));
  bfr _b_4292(.a(_w_6194),.q(_w_6195));
  bfr _b_4290(.a(_w_6192),.q(_w_6193));
  bfr _b_6383(.a(_w_8285),.q(_w_8286));
  bfr _b_7819(.a(_w_9721),.q(_w_9722));
  bfr _b_4289(.a(_w_6191),.q(n706_1));
  bfr _b_4550(.a(_w_6452),.q(_w_6453));
  bfr _b_7250(.a(_w_9152),.q(_w_9153));
  bfr _b_4284(.a(_w_6186),.q(_w_6187));
  bfr _b_6871(.a(_w_8773),.q(n1301));
  bfr _b_4282(.a(_w_6184),.q(n1194_1));
  bfr _b_4281(.a(_w_6183),.q(_w_6184));
  bfr _b_4384(.a(_w_6286),.q(_w_6287));
  bfr _b_4279(.a(_w_6181),.q(_w_6182));
  bfr _b_14326(.a(_w_16228),.q(_w_16229));
  bfr _b_4357(.a(_w_6259),.q(_w_6260));
  and_bb g635(.a(N222_13),.b(N290_17),.q(n635));
  bfr _b_11555(.a(_w_13457),.q(_w_13458));
  bfr _b_7261(.a(_w_9163),.q(_w_9164));
  bfr _b_4276(.a(_w_6178),.q(_w_6179));
  bfr _b_4751(.a(_w_6653),.q(N1_14));
  bfr _b_4274(.a(_w_6176),.q(n112_1));
  spl2 g814_s_0(.a(n814),.q0(n814_0),.q1(_w_7463));
  bfr _b_5005(.a(_w_6907),.q(_w_6908));
  bfr _b_4268(.a(_w_6170),.q(_w_6171));
  bfr _b_5935(.a(_w_7837),.q(_w_7838));
  bfr _b_11920(.a(_w_13822),.q(_w_13823));
  bfr _b_4266(.a(_w_6168),.q(n742_1));
  bfr _b_14234(.a(_w_16136),.q(_w_16137));
  bfr _b_6878(.a(_w_8780),.q(n861));
  bfr _b_14278(.a(_w_16180),.q(_w_16181));
  bfr _b_4320(.a(_w_6222),.q(_w_6223));
  bfr _b_4257(.a(_w_6159),.q(_w_6160));
  bfr _b_4254(.a(_w_6156),.q(n1686_1));
  bfr _b_4253(.a(_w_6155),.q(_w_6156));
  bfr _b_4251(.a(_w_6153),.q(_w_6154));
  bfr _b_4246(.a(_w_6148),.q(N171_11));
  bfr _b_9799(.a(_w_11701),.q(_w_11702));
  bfr _b_5864(.a(_w_7766),.q(_w_7767));
  bfr _b_4231(.a(_w_6133),.q(_w_6134));
  bfr _b_8035(.a(_w_9937),.q(_w_9938));
  bfr _b_4227(.a(_w_6129),.q(_w_6130));
  bfr _b_11178(.a(_w_13080),.q(_w_13081));
  or_bb g1230(.a(n1172_0),.b(n1229_0),.q(n1230));
  bfr _b_4224(.a(_w_6126),.q(_w_6127));
  bfr _b_4219(.a(_w_6121),.q(_w_6122));
  bfr _b_4212(.a(_w_6114),.q(_w_6115));
  spl2 g1388_s_0(.a(n1388),.q0(n1388_0),.q1(n1388_1));
  bfr _b_4822(.a(_w_6724),.q(_w_6725));
  and_bi g774(.a(n772_0),.b(n773),.q(n774));
  bfr _b_4211(.a(_w_6113),.q(_w_6114));
  bfr _b_4209(.a(_w_6111),.q(_w_6112));
  spl4L N324_s_2(.a(N324_1),.q0(N324_8),.q1(N324_9),.q2(N324_10),.q3(N324_11));
  bfr _b_4208(.a(_w_6110),.q(_w_6111));
  bfr _b_11151(.a(_w_13053),.q(_w_13054));
  and_bi g744(.a(n742_0),.b(n743),.q(n744));
  bfr _b_9901(.a(_w_11803),.q(_w_11804));
  bfr _b_4206(.a(_w_6108),.q(_w_6109));
  bfr _b_4205(.a(_w_6107),.q(_w_6108));
  bfr _b_4984(.a(_w_6886),.q(_w_6887));
  bfr _b_4199(.a(_w_6101),.q(_w_6102));
  bfr _b_13266(.a(_w_15168),.q(_w_15169));
  bfr _b_4382(.a(_w_6284),.q(_w_6285));
  bfr _b_13223(.a(_w_15125),.q(_w_15126));
  bfr _b_3910(.a(_w_5812),.q(_w_5813));
  bfr _b_5181(.a(_w_7083),.q(_w_7084));
  bfr _b_4193(.a(_w_6095),.q(_w_6096));
  bfr _b_4191(.a(_w_6093),.q(_w_6094));
  bfr _b_7358(.a(_w_9260),.q(n1659_1));
  and_bb g1387(.a(n1384_1),.b(n1385_1),.q(_w_13560));
  bfr _b_4186(.a(_w_6088),.q(n852_1));
  bfr _b_4263(.a(_w_6165),.q(_w_6166));
  spl2 g210_s_0(.a(n210),.q0(n210_0),.q1(n210_1));
  bfr _b_4184(.a(_w_6086),.q(_w_6087));
  bfr _b_5159(.a(_w_7061),.q(n796_1));
  bfr _b_7873(.a(_w_9775),.q(_w_9776));
  bfr _b_4183(.a(_w_6085),.q(_w_6086));
  bfr _b_7462(.a(_w_9364),.q(_w_9365));
  bfr _b_8960(.a(_w_10862),.q(_w_10863));
  bfr _b_4182(.a(_w_6084),.q(n875_1));
  bfr _b_13473(.a(_w_15375),.q(_w_15376));
  bfr _b_4786(.a(_w_6688),.q(_w_6689));
  or_bb g1752(.a(n1750_0),.b(n1751),.q(n1752));
  bfr _b_4175(.a(_w_6077),.q(_w_6078));
  bfr _b_4172(.a(_w_6074),.q(_w_6075));
  bfr _b_3697(.a(_w_5599),.q(_w_5600));
  spl2 g459_s_0(.a(n459),.q0(n459_0),.q1(n459_1));
  and_bb g944(.a(N460_9),.b(N86_15),.q(_w_11134));
  bfr _b_9245(.a(_w_11147),.q(_w_11148));
  bfr _b_4541(.a(_w_6443),.q(_w_6444));
  spl2 g762_s_0(.a(n762),.q0(n762_0),.q1(n762_1));
  bfr _b_14053(.a(_w_15955),.q(_w_15956));
  bfr _b_4166(.a(_w_6068),.q(_w_6069));
  bfr _b_7863(.a(_w_9765),.q(_w_9766));
  bfr _b_8291(.a(_w_10193),.q(_w_10194));
  bfr _b_4160(.a(_w_6062),.q(_w_6063));
  bfr _b_4158(.a(_w_6060),.q(_w_6061));
  and_bi g1729(.a(n1716_1),.b(n1719_1),.q(_w_10149));
  bfr _b_4587(.a(_w_6489),.q(N154_1));
  bfr _b_4154(.a(_w_6056),.q(_w_6057));
  bfr _b_4147(.a(_w_6049),.q(_w_6050));
  bfr _b_3986(.a(_w_5888),.q(_w_5889));
  bfr _b_9259(.a(_w_11161),.q(_w_11162));
  bfr _b_4145(.a(_w_6047),.q(_w_6048));
  bfr _b_9095(.a(_w_10997),.q(_w_10998));
  bfr _b_4142(.a(_w_6044),.q(_w_6045));
  and_bi g1147(.a(n1052_1),.b(n1145_1),.q(_w_11577));
  bfr _b_4862(.a(_w_6764),.q(_w_6765));
  bfr _b_4133(.a(_w_6035),.q(_w_6036));
  bfr _b_4132(.a(_w_6034),.q(_w_6035));
  bfr _b_4131(.a(_w_6033),.q(_w_6034));
  bfr _b_4931(.a(_w_6833),.q(_w_6834));
  bfr _b_4122(.a(_w_6024),.q(_w_6025));
  bfr _b_3778(.a(_w_5680),.q(_w_5681));
  bfr _b_4114(.a(_w_6016),.q(_w_6017));
  bfr _b_4112(.a(_w_6014),.q(_w_6015));
  bfr _b_4109(.a(_w_6011),.q(_w_6012));
  bfr _b_4108(.a(_w_6010),.q(_w_6011));
  bfr _b_4104(.a(_w_6006),.q(_w_6007));
  and_bi g1689(.a(n1688_0),.b(n1683_0),.q(n1689));
  bfr _b_4103(.a(_w_6005),.q(_w_6006));
  bfr _b_4102(.a(_w_6004),.q(_w_6005));
  bfr _b_4089(.a(_w_5991),.q(_w_5992));
  bfr _b_4349(.a(_w_6251),.q(_w_6252));
  spl2 g502_s_0(.a(n502),.q0(n502_0),.q1(_w_7881));
  bfr _b_8853(.a(_w_10755),.q(_w_10756));
  bfr _b_4087(.a(_w_5989),.q(_w_5990));
  spl2 g170_s_0(.a(n170),.q0(n170_0),.q1(n170_1));
  bfr _b_4085(.a(_w_5987),.q(_w_5988));
  or_bb g412(.a(n367_0),.b(n411_0),.q(n412));
  bfr _b_11478(.a(_w_13380),.q(_w_13381));
  bfr _b_10761(.a(_w_12663),.q(_w_12664));
  bfr _b_10738(.a(_w_12640),.q(_w_12641));
  bfr _b_8567(.a(_w_10469),.q(_w_10470));
  bfr _b_4081(.a(_w_5983),.q(_w_5984));
  bfr _b_14199(.a(_w_16101),.q(_w_16102));
  bfr _b_4076(.a(_w_5978),.q(_w_5979));
  bfr _b_10444(.a(_w_12346),.q(n1058));
  or_bb g1746(.a(n1744_0),.b(n1745),.q(n1746));
  bfr _b_4075(.a(_w_5977),.q(_w_5978));
  bfr _b_4070(.a(_w_5972),.q(_w_5973));
  spl2 g841_s_0(.a(n841),.q0(n841_0),.q1(n841_1));
  bfr _b_4061(.a(_w_5963),.q(_w_5964));
  bfr _b_14034(.a(_w_15936),.q(_w_15937));
  bfr _b_4058(.a(_w_5960),.q(_w_5961));
  bfr _b_4051(.a(_w_5953),.q(_w_5954));
  bfr _b_5013(.a(_w_6915),.q(_w_6916));
  bfr _b_4047(.a(_w_5949),.q(_w_5950));
  bfr _b_4044(.a(_w_5946),.q(_w_5947));
  and_bi g1450(.a(n1363_1),.b(n1448_1),.q(_w_13769));
  and_bi g1287(.a(n1194_1),.b(n1197_1),.q(n1287));
  bfr _b_4043(.a(_w_5945),.q(_w_5946));
  bfr _b_7205(.a(_w_9107),.q(_w_9108));
  bfr _b_4038(.a(_w_5940),.q(_w_5941));
  bfr _b_4037(.a(_w_5939),.q(_w_5940));
  bfr _b_4036(.a(_w_5938),.q(_w_5939));
  bfr _b_4527(.a(_w_6429),.q(N137_7));
  bfr _b_4034(.a(_w_5936),.q(N239_1));
  bfr _b_4385(.a(_w_6287),.q(n202_1));
  bfr _b_4033(.a(_w_5935),.q(_w_5936));
  bfr _b_4472(.a(_w_6374),.q(_w_6375));
  bfr _b_11823(.a(_w_13725),.q(_w_13726));
  or_bb g65(.a(n63_0),.b(n64),.q(n65));
  bfr _b_4030(.a(_w_5932),.q(_w_5933));
  bfr _b_4026(.a(_w_5928),.q(_w_5929));
  bfr _b_14104(.a(_w_16006),.q(_w_16007));
  bfr _b_12479(.a(_w_14381),.q(_w_14382));
  bfr _b_8143(.a(_w_10045),.q(_w_10046));
  bfr _b_4021(.a(_w_5923),.q(_w_5924));
  bfr _b_13013(.a(_w_14915),.q(_w_14916));
  bfr _b_4019(.a(_w_5921),.q(_w_5922));
  bfr _b_3416(.a(_w_5318),.q(_w_5319));
  bfr _b_10253(.a(_w_12155),.q(_w_12156));
  bfr _b_4005(.a(_w_5907),.q(_w_5908));
  bfr _b_13550(.a(_w_15452),.q(_w_15453));
  bfr _b_5908(.a(_w_7810),.q(_w_7811));
  bfr _b_4433(.a(_w_6335),.q(_w_6336));
  bfr _b_4651(.a(_w_6553),.q(_w_6554));
  spl2 g893_s_0(.a(n893),.q0(n893_0),.q1(_w_6157));
  bfr _b_12006(.a(_w_13908),.q(_w_13909));
  bfr _b_3996(.a(_w_5898),.q(_w_5899));
  bfr _b_3995(.a(_w_5897),.q(_w_5898));
  bfr _b_3993(.a(_w_5895),.q(_w_5896));
  bfr _b_12017(.a(_w_13919),.q(_w_13920));
  bfr _b_3987(.a(_w_5889),.q(_w_5890));
  bfr _b_6982(.a(_w_8884),.q(_w_8885));
  bfr _b_3983(.a(_w_5885),.q(_w_5886));
  and_bi g1632(.a(n1631_0),.b(n1618_0),.q(n1632));
  bfr _b_9026(.a(_w_10928),.q(_w_10929));
  spl4L N256_s_3(.a(N256_2),.q0(_w_8036),.q1(N256_13),.q2(_w_8085),.q3(_w_8102));
  bfr _b_6154(.a(_w_8056),.q(_w_8057));
  bfr _b_3980(.a(_w_5882),.q(_w_5883));
  bfr _b_5066(.a(_w_6968),.q(_w_6969));
  bfr _b_3979(.a(_w_5881),.q(_w_5882));
  bfr _b_9741(.a(_w_11643),.q(_w_11644));
  bfr _b_13317(.a(_w_15219),.q(_w_15220));
  bfr _b_4394(.a(_w_6296),.q(_w_6297));
  bfr _b_3975(.a(_w_5877),.q(_w_5878));
  spl4L N86_s_4(.a(N86_3),.q0(N86_16),.q1(N86_17),.q2(N86_18),.q3(N86_19));
  bfr _b_3973(.a(_w_5875),.q(_w_5876));
  bfr _b_3494(.a(_w_5396),.q(_w_5397));
  bfr _b_4244(.a(_w_6146),.q(_w_6147));
  bfr _b_7583(.a(_w_9485),.q(_w_9486));
  bfr _b_3972(.a(_w_5874),.q(_w_5875));
  bfr _b_3971(.a(_w_5873),.q(_w_5874));
  bfr _b_3969(.a(_w_5871),.q(_w_5872));
  bfr _b_3966(.a(_w_5868),.q(_w_5869));
  spl2 g1478_s_0(.a(n1478),.q0(n1478_0),.q1(n1478_1));
  bfr _b_10904(.a(_w_12806),.q(_w_12807));
  bfr _b_4950(.a(_w_6852),.q(_w_6853));
  or_bb g342(.a(n297_0),.b(n341_0),.q(n342));
  bfr _b_3961(.a(_w_5863),.q(_w_5864));
  bfr _b_3539(.a(_w_5441),.q(_w_5442));
  bfr _b_3994(.a(_w_5896),.q(_w_5897));
  bfr _b_3958(.a(_w_5860),.q(N239_13));
  bfr _b_13410(.a(_w_15312),.q(_w_15313));
  bfr _b_4806(.a(_w_6708),.q(_w_6709));
  bfr _b_3957(.a(_w_5859),.q(_w_5860));
  bfr _b_3956(.a(_w_5858),.q(_w_5859));
  bfr _b_10006(.a(_w_11908),.q(_w_11909));
  bfr _b_3954(.a(_w_5856),.q(_w_5857));
  bfr _b_4258(.a(_w_6160),.q(n893_1));
  and_bi g338(.a(n336_0),.b(n337),.q(n338));
  bfr _b_8593(.a(_w_10495),.q(_w_10496));
  bfr _b_11636(.a(_w_13538),.q(_w_13539));
  bfr _b_3953(.a(_w_5855),.q(_w_5856));
  bfr _b_3951(.a(_w_5853),.q(_w_5854));
  bfr _b_6316(.a(_w_8218),.q(_w_8219));
  bfr _b_3947(.a(_w_5849),.q(_w_5850));
  bfr _b_8697(.a(_w_10599),.q(n546_1));
  bfr _b_9400(.a(_w_11302),.q(_w_11303));
  bfr _b_3940(.a(_w_5842),.q(_w_5843));
  bfr _b_3590(.a(_w_5492),.q(_w_5493));
  bfr _b_9942(.a(_w_11844),.q(_w_11845));
  bfr _b_3935(.a(_w_5837),.q(_w_5838));
  spl2 g1118_s_0(.a(n1118),.q0(n1118_0),.q1(n1118_1));
  bfr _b_7053(.a(_w_8955),.q(n782));
  bfr _b_4471(.a(_w_6373),.q(n784_1));
  bfr _b_7439(.a(_w_9341),.q(_w_9342));
  bfr _b_4107(.a(_w_6009),.q(_w_6010));
  spl2 g1164_s_0(.a(n1164),.q0(n1164_0),.q1(n1164_1));
  bfr _b_11361(.a(_w_13263),.q(_w_13264));
  bfr _b_5195(.a(_w_7097),.q(_w_7098));
  bfr _b_3928(.a(_w_5830),.q(n980_1));
  bfr _b_4317(.a(_w_6219),.q(N120_13));
  and_bb g1855(.a(N239_18),.b(N511_18),.q(_w_14658));
  bfr _b_11813(.a(_w_13715),.q(_w_13716));
  bfr _b_10061(.a(_w_11963),.q(_w_11964));
  bfr _b_8304(.a(_w_10206),.q(n157));
  bfr _b_3923(.a(_w_5825),.q(_w_5826));
  bfr _b_3920(.a(_w_5822),.q(_w_5823));
  bfr _b_13641(.a(_w_15543),.q(_w_15544));
  bfr _b_5177(.a(_w_7079),.q(_w_7080));
  bfr _b_3917(.a(_w_5819),.q(N256_2));
  bfr _b_4176(.a(_w_6078),.q(_w_6079));
  spl2 g1274_s_0(.a(n1274),.q0(n1274_0),.q1(n1274_1));
  bfr _b_4604(.a(_w_6506),.q(_w_6507));
  bfr _b_10634(.a(_w_12536),.q(_w_12537));
  bfr _b_3915(.a(_w_5817),.q(_w_5818));
  bfr _b_3913(.a(_w_5815),.q(_w_5816));
  bfr _b_6406(.a(_w_8308),.q(_w_8309));
  bfr _b_11670(.a(_w_13572),.q(_w_13573));
  bfr _b_3909(.a(_w_5811),.q(_w_5812));
  bfr _b_9900(.a(_w_11802),.q(_w_11803));
  bfr _b_14144(.a(_w_16046),.q(_w_16047));
  bfr _b_3907(.a(_w_5809),.q(_w_5810));
  bfr _b_5071(.a(_w_6973),.q(_w_6974));
  bfr _b_13990(.a(_w_15892),.q(_w_15893));
  bfr _b_11974(.a(_w_13876),.q(_w_13877));
  bfr _b_3906(.a(_w_5808),.q(_w_5809));
  bfr _b_9255(.a(_w_11157),.q(n1543));
  bfr _b_3902(.a(_w_5804),.q(_w_5805));
  bfr _b_3901(.a(_w_5803),.q(_w_5804));
  bfr _b_3900(.a(_w_5802),.q(_w_5803));
  bfr _b_3895(.a(_w_5797),.q(_w_5798));
  bfr _b_4123(.a(_w_6025),.q(_w_6026));
  bfr _b_3890(.a(_w_5792),.q(_w_5793));
  bfr _b_3458(.a(_w_5360),.q(_w_5361));
  bfr _b_3887(.a(_w_5789),.q(_w_5790));
  bfr _b_4940(.a(_w_6842),.q(_w_6843));
  bfr _b_11139(.a(_w_13041),.q(_w_13042));
  bfr _b_3886(.a(_w_5788),.q(_w_5789));
  bfr _b_3884(.a(_w_5786),.q(_w_5787));
  bfr _b_11857(.a(_w_13759),.q(_w_13760));
  bfr _b_3882(.a(_w_5784),.q(_w_5785));
  spl2 g920_s_0(.a(n920),.q0(n920_0),.q1(n920_1));
  bfr _b_4412(.a(_w_6314),.q(_w_6315));
  bfr _b_7204(.a(_w_9106),.q(_w_9107));
  bfr _b_11761(.a(_w_13663),.q(_w_13664));
  bfr _b_4007(.a(_w_5909),.q(_w_5910));
  bfr _b_3877(.a(_w_5779),.q(_w_5780));
  and_bi g1390(.a(n1383_1),.b(n1388_1),.q(_w_13561));
  bfr _b_8619(.a(_w_10521),.q(_w_10522));
  bfr _b_3873(.a(_w_5775),.q(_w_5776));
  bfr _b_4434(.a(_w_6336),.q(_w_6337));
  and_bi g1733(.a(n1704_1),.b(n1707_1),.q(n1733));
  bfr _b_3867(.a(_w_5769),.q(_w_5770));
  bfr _b_3865(.a(_w_5767),.q(_w_5768));
  bfr _b_4100(.a(_w_6002),.q(_w_6003));
  bfr _b_3855(.a(_w_5757),.q(_w_5758));
  bfr _b_9046(.a(_w_10948),.q(_w_10949));
  bfr _b_3850(.a(_w_5752),.q(_w_5753));
  and_bb g1060(.a(N120_14),.b(N443_11),.q(_w_9368));
  and_bi g1372(.a(n1327_1),.b(n1330_1),.q(n1372));
  bfr _b_3842(.a(_w_5744),.q(_w_5745));
  bfr _b_3779(.a(_w_5681),.q(_w_5682));
  bfr _b_7375(.a(_w_9277),.q(n1434_1));
  bfr _b_8592(.a(_w_10494),.q(_w_10495));
  bfr _b_3841(.a(_w_5743),.q(_w_5744));
  bfr _b_10598(.a(_w_12500),.q(_w_12501));
  bfr _b_3840(.a(_w_5742),.q(_w_5743));
  or_bb g1703(.a(n1701_0),.b(n1702),.q(n1703));
  bfr _b_4001(.a(_w_5903),.q(_w_5904));
  bfr _b_4679(.a(_w_6581),.q(_w_6582));
  bfr _b_3831(.a(_w_5733),.q(_w_5734));
  bfr _b_8466(.a(_w_10368),.q(_w_10369));
  bfr _b_11691(.a(_w_13593),.q(_w_13594));
  bfr _b_3827(.a(_w_5729),.q(_w_5730));
  and_bb g960(.a(N222_17),.b(N324_17),.q(_w_9739));
  bfr _b_3825(.a(_w_5727),.q(_w_5728));
  spl2 g441_s_0(.a(n441),.q0(n441_0),.q1(n441_1));
  bfr _b_5157(.a(_w_7059),.q(_w_7060));
  bfr _b_3821(.a(_w_5723),.q(_w_5724));
  and_bb g737(.a(N239_4),.b(N290_18),.q(n737));
  bfr _b_5626(.a(_w_7528),.q(_w_7529));
  bfr _b_12577(.a(_w_14479),.q(_w_14480));
  bfr _b_3817(.a(_w_5719),.q(_w_5720));
  bfr _b_3813(.a(_w_5715),.q(_w_5716));
  bfr _b_6087(.a(_w_7989),.q(_w_7990));
  bfr _b_13928(.a(_w_15830),.q(_w_15831));
  bfr _b_4134(.a(_w_6036),.q(_w_6037));
  bfr _b_3811(.a(_w_5713),.q(_w_5714));
  bfr _b_12547(.a(_w_14449),.q(_w_14450));
  bfr _b_3810(.a(_w_5712),.q(_w_5713));
  bfr _b_13039(.a(_w_14941),.q(_w_14942));
  bfr _b_3807(.a(_w_5709),.q(_w_5710));
  bfr _b_11150(.a(_w_13052),.q(_w_13053));
  bfr _b_9562(.a(_w_11464),.q(_w_11465));
  bfr _b_11374(.a(_w_13276),.q(_w_13277));
  bfr _b_3804(.a(_w_5706),.q(_w_5707));
  bfr _b_4020(.a(_w_5922),.q(_w_5923));
  bfr _b_11278(.a(_w_13180),.q(_w_13181));
  bfr _b_10879(.a(_w_12781),.q(_w_12782));
  bfr _b_10058(.a(_w_11960),.q(_w_11961));
  bfr _b_3800(.a(_w_5702),.q(_w_5703));
  bfr _b_3799(.a(_w_5701),.q(_w_5702));
  bfr _b_3798(.a(_w_5700),.q(_w_5701));
  bfr _b_11339(.a(_w_13241),.q(_w_13242));
  bfr _b_3796(.a(_w_5698),.q(N256_7));
  spl2 g1092_s_0(.a(n1092),.q0(n1092_0),.q1(n1092_1));
  and_bb g419(.a(n365_1),.b(n417_1),.q(_w_9685));
  bfr _b_3792(.a(_w_5694),.q(_w_5695));
  and_bi g821(.a(n814_1),.b(n817_1),.q(n821));
  and_bi g1626(.a(n1625_0),.b(n1620_0),.q(n1626));
  bfr _b_3784(.a(_w_5686),.q(_w_5687));
  bfr _b_12068(.a(_w_13970),.q(n1624));
  bfr _b_3781(.a(_w_5683),.q(_w_5684));
  bfr _b_3777(.a(_w_5679),.q(_w_5680));
  bfr _b_3776(.a(_w_5678),.q(_w_5679));
  spl2 g1700_s_0(.a(n1700),.q0(n1700_0),.q1(n1700_1));
  bfr _b_3773(.a(_w_5675),.q(_w_5676));
  and_bi g1568(.a(n1545_1),.b(n1566_1),.q(_w_14968));
  bfr _b_3770(.a(_w_5672),.q(_w_5673));
  bfr _b_4440(.a(_w_6342),.q(_w_6343));
  spl2 g868_s_0(.a(n868),.q0(n868_0),.q1(n868_1));
  spl2 g1436_s_0(.a(n1436),.q0(n1436_0),.q1(n1436_1));
  bfr _b_13399(.a(_w_15301),.q(_w_15302));
  bfr _b_4267(.a(_w_6169),.q(_w_6170));
  bfr _b_8784(.a(_w_10686),.q(_w_10687));
  bfr _b_11014(.a(_w_12916),.q(_w_12917));
  bfr _b_3765(.a(_w_5667),.q(_w_5668));
  bfr _b_9131(.a(_w_11033),.q(_w_11034));
  bfr _b_3762(.a(_w_5664),.q(_w_5665));
  bfr _b_3761(.a(_w_5663),.q(_w_5664));
  bfr _b_4197(.a(_w_6099),.q(_w_6100));
  bfr _b_3760(.a(_w_5662),.q(N256_6));
  bfr _b_3899(.a(_w_5801),.q(_w_5802));
  bfr _b_3837(.a(_w_5739),.q(_w_5740));
  bfr _b_13363(.a(_w_15265),.q(_w_15266));
  bfr _b_11026(.a(_w_12928),.q(_w_12929));
  bfr _b_3754(.a(_w_5656),.q(_w_5657));
  bfr _b_3753(.a(_w_5655),.q(_w_5656));
  bfr _b_3747(.a(_w_5649),.q(_w_5650));
  bfr _b_4300(.a(_w_6202),.q(_w_6203));
  spl2 g1034_s_0(.a(n1034),.q0(n1034_0),.q1(_w_5555));
  and_bi g548(.a(n546_0),.b(n547),.q(n548));
  bfr _b_3745(.a(_w_5647),.q(_w_5648));
  bfr _b_4006(.a(_w_5908),.q(N239_11));
  bfr _b_3571(.a(_w_5473),.q(_w_5474));
  bfr _b_13750(.a(_w_15652),.q(_w_15653));
  spl2 g820_s_0(.a(n820),.q0(n820_0),.q1(n820_1));
  bfr _b_3742(.a(_w_5644),.q(_w_5645));
  bfr _b_4721(.a(_w_6623),.q(_w_6624));
  or_bb g1326(.a(n1324_0),.b(n1325),.q(n1326));
  bfr _b_3739(.a(_w_5641),.q(_w_5642));
  bfr _b_9718(.a(_w_11620),.q(_w_11621));
  or_bb g1333(.a(n1275_0),.b(n1332_0),.q(n1333));
  bfr _b_8532(.a(_w_10434),.q(_w_10435));
  bfr _b_10899(.a(_w_12801),.q(_w_12802));
  bfr _b_3736(.a(_w_5638),.q(_w_5639));
  bfr _b_4194(.a(_w_6096),.q(_w_6097));
  bfr _b_3602(.a(_w_5504),.q(_w_5505));
  bfr _b_13405(.a(_w_15307),.q(_w_15308));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  or_bb g219(.a(n217_0),.b(n218),.q(n219));
  bfr _b_4746(.a(_w_6648),.q(_w_6649));
  bfr _b_5016(.a(_w_6918),.q(_w_6919));
  bfr _b_3669(.a(_w_5571),.q(_w_5572));
  bfr _b_3727(.a(_w_5629),.q(_w_5630));
  bfr _b_3714(.a(_w_5616),.q(_w_5617));
  bfr _b_5093(.a(_w_6995),.q(_w_6996));
  bfr _b_10552(.a(_w_12454),.q(_w_12455));
  bfr _b_6877(.a(_w_8779),.q(n912));
  bfr _b_3706(.a(_w_5608),.q(_w_5609));
  bfr _b_3703(.a(_w_5605),.q(_w_5606));
  bfr _b_12683(.a(_w_14585),.q(_w_14586));
  bfr _b_4121(.a(_w_6023),.q(_w_6024));
  spl2 g793_s_0(.a(n793),.q0(n793_0),.q1(n793_1));
  bfr _b_3702(.a(_w_5604),.q(_w_5605));
  bfr _b_3701(.a(_w_5603),.q(_w_5604));
  bfr _b_10690(.a(_w_12592),.q(_w_12593));
  bfr _b_5868(.a(_w_7770),.q(_w_7771));
  bfr _b_8594(.a(_w_10496),.q(_w_10497));
  bfr _b_8677(.a(_w_10579),.q(_w_10580));
  bfr _b_13901(.a(_w_15803),.q(_w_15804));
  bfr _b_11033(.a(_w_12935),.q(_w_12936));
  bfr _b_3695(.a(_w_5597),.q(_w_5598));
  bfr _b_4476(.a(_w_6378),.q(_w_6379));
  spl2 g1395_s_0(.a(n1395),.q0(n1395_0),.q1(n1395_1));
  bfr _b_3691(.a(_w_5593),.q(_w_5594));
  bfr _b_7744(.a(_w_9646),.q(_w_9647));
  bfr _b_5027(.a(_w_6929),.q(_w_6930));
  bfr _b_11849(.a(_w_13751),.q(n580));
  spl2 g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1));
  bfr _b_10270(.a(_w_12172),.q(_w_12173));
  bfr _b_3681(.a(_w_5583),.q(_w_5584));
  spl2 g890_s_0(.a(n890),.q0(n890_0),.q1(n890_1));
  bfr _b_5775(.a(_w_7677),.q(_w_7678));
  bfr _b_3678(.a(_w_5580),.q(_w_5581));
  bfr _b_7051(.a(_w_8953),.q(_w_8954));
  bfr _b_3677(.a(_w_5579),.q(_w_5580));
  bfr _b_7794(.a(_w_9696),.q(_w_9697));
  bfr _b_5576(.a(_w_7478),.q(n82_1));
  bfr _b_10104(.a(_w_12006),.q(_w_12007));
  bfr _b_3670(.a(_w_5572),.q(_w_5573));
  bfr _b_3668(.a(_w_5570),.q(_w_5571));
  bfr _b_3667(.a(_w_5569),.q(_w_5570));
  and_bb g671(.a(n625_1),.b(n669_1),.q(_w_8774));
  or_bb g1142(.a(n1140_0),.b(n1141),.q(n1142));
  bfr _b_3661(.a(_w_5563),.q(_w_5564));
  bfr _b_13667(.a(_w_15569),.q(_w_15545));
  or_bb g1265(.a(n1263_0),.b(n1264),.q(_w_13377));
  bfr _b_3658(.a(_w_5560),.q(n33_0));
  bfr _b_13666(.a(_w_15568),.q(_w_15569));
  bfr _b_6512(.a(_w_8414),.q(N205_1));
  bfr _b_3651(.a(_w_5553),.q(_w_5554));
  and_bi g468(.a(n466_0),.b(n467),.q(n468));
  spl2 g954_s_0(.a(n954),.q0(n954_0),.q1(n954_1));
  bfr _b_3643(.a(_w_5545),.q(_w_5546));
  and_bi g685(.a(n684_0),.b(n620_0),.q(n685));
  bfr _b_5700(.a(_w_7602),.q(_w_7603));
  bfr _b_11296(.a(_w_13198),.q(n80));
  and_bi g649(.a(n648_0),.b(n632_0),.q(n649));
  bfr _b_5112(.a(_w_7014),.q(_w_7015));
  bfr _b_9827(.a(_w_11729),.q(_w_11730));
  bfr _b_3637(.a(_w_5539),.q(_w_5540));
  bfr _b_3633(.a(_w_5535),.q(_w_5536));
  bfr _b_3630(.a(_w_5532),.q(_w_5533));
  bfr _b_3629(.a(_w_5531),.q(_w_5532));
  and_bi g1238(.a(n1236_0),.b(n1237),.q(n1238));
  bfr _b_4934(.a(_w_6836),.q(_w_6837));
  bfr _b_3624(.a(_w_5526),.q(_w_5527));
  spl4L N426_s_0(.a(_w_15727),.q0(N426_0),.q1(N426_1),.q2(N426_2),.q3(N426_3));
  bfr _b_6291(.a(_w_8193),.q(_w_8194));
  bfr _b_11763(.a(_w_13665),.q(_w_13666));
  bfr _b_6245(.a(_w_8147),.q(_w_8148));
  bfr _b_3619(.a(_w_5521),.q(_w_5522));
  bfr _b_8274(.a(_w_10176),.q(_w_10177));
  bfr _b_3617(.a(_w_5519),.q(_w_5520));
  bfr _b_9159(.a(_w_11061),.q(n128));
  bfr _b_3616(.a(_w_5518),.q(_w_5519));
  bfr _b_3615(.a(_w_5517),.q(_w_5518));
  bfr _b_4376(.a(_w_6278),.q(_w_6279));
  bfr _b_3614(.a(_w_5516),.q(_w_5517));
  spl2 g385_s_0(.a(n385),.q0(n385_0),.q1(n385_1));
  bfr _b_3611(.a(_w_5513),.q(_w_5514));
  bfr _b_3607(.a(_w_5509),.q(_w_5510));
  bfr _b_12989(.a(_w_14891),.q(_w_14892));
  bfr _b_3606(.a(_w_5508),.q(_w_5509));
  bfr _b_3598(.a(_w_5500),.q(_w_5501));
  bfr _b_6499(.a(_w_8401),.q(_w_8402));
  bfr _b_3594(.a(_w_5496),.q(_w_5497));
  bfr _b_3593(.a(_w_5495),.q(_w_5496));
  bfr _b_3592(.a(_w_5494),.q(_w_5495));
  and_bb g292(.a(N1_13),.b(N426_4),.q(n292));
  bfr _b_11995(.a(_w_13897),.q(_w_13898));
  bfr _b_10907(.a(_w_12809),.q(_w_12810));
  bfr _b_9494(.a(_w_11396),.q(_w_11397));
  bfr _b_3585(.a(_w_5487),.q(_w_5488));
  spl2 g907_s_0(.a(n907),.q0(n907_0),.q1(n907_1));
  bfr _b_14124(.a(_w_16026),.q(_w_16027));
  bfr _b_8402(.a(_w_10304),.q(n634));
  bfr _b_3583(.a(_w_5485),.q(_w_5486));
  bfr _b_11490(.a(_w_13392),.q(_w_13393));
  bfr _b_3582(.a(_w_5484),.q(_w_5485));
  bfr _b_10962(.a(_w_12864),.q(_w_12865));
  bfr _b_4684(.a(_w_6586),.q(_w_6587));
  bfr _b_5024(.a(_w_6926),.q(_w_6927));
  spl2 g309_s_0(.a(n309),.q0(n309_0),.q1(n309_1));
  bfr _b_10251(.a(_w_12153),.q(_w_12154));
  bfr _b_3575(.a(_w_5477),.q(_w_5478));
  and_bi g453(.a(n382_1),.b(n385_1),.q(n453));
  bfr _b_4896(.a(_w_6798),.q(_w_6799));
  or_bb g1594(.a(n1536_0),.b(n1593_0),.q(n1594));
  bfr _b_10363(.a(_w_12265),.q(_w_12266));
  bfr _b_3659(.a(_w_5561),.q(_w_5562));
  bfr _b_12536(.a(_w_14438),.q(_w_14439));
  or_bb g1223(.a(n1221_0),.b(n1222),.q(n1223));
  bfr _b_3569(.a(_w_5471),.q(_w_5472));
  bfr _b_12120(.a(_w_14022),.q(_w_14023));
  bfr _b_10408(.a(_w_12310),.q(n337));
  bfr _b_3846(.a(_w_5748),.q(N256_0));
  bfr _b_14215(.a(_w_16117),.q(_w_16118));
  bfr _b_5381(.a(_w_7283),.q(_w_7284));
  bfr _b_6707(.a(_w_8609),.q(_w_8610));
  bfr _b_8295(.a(_w_10197),.q(_w_10198));
  bfr _b_8578(.a(_w_10480),.q(_w_10481));
  bfr _b_3566(.a(_w_5468),.q(_w_5469));
  and_bi g1554(.a(n1552_0),.b(n1553),.q(n1554));
  bfr _b_3564(.a(_w_5466),.q(_w_5467));
  bfr _b_3853(.a(_w_5755),.q(_w_5756));
  bfr _b_3562(.a(_w_5464),.q(_w_5465));
  bfr _b_3561(.a(_w_5463),.q(_w_5464));
  and_bb g1681(.a(N222_9),.b(N460_17),.q(_w_13137));
  bfr _b_6916(.a(_w_8818),.q(_w_8819));
  bfr _b_7199(.a(_w_9101),.q(_w_9102));
  bfr _b_5067(.a(_w_6969),.q(_w_6970));
  bfr _b_3556(.a(_w_5458),.q(_w_5459));
  or_bb g1160(.a(n1158_0),.b(n1159),.q(_w_11174));
  and_bb g147(.a(N103_5),.b(N273_10),.q(n147));
  bfr _b_6958(.a(_w_8860),.q(_w_8861));
  and_bi g1475(.a(n1473_0),.b(n1474),.q(n1475));
  bfr _b_3548(.a(_w_5450),.q(N52_2));
  bfr _b_10297(.a(_w_12199),.q(_w_12200));
  bfr _b_4667(.a(_w_6569),.q(_w_6570));
  bfr _b_4575(.a(_w_6477),.q(_w_6478));
  bfr _b_3544(.a(_w_5446),.q(_w_5447));
  bfr _b_12552(.a(_w_14454),.q(_w_14455));
  bfr _b_10658(.a(_w_12560),.q(_w_12561));
  bfr _b_3543(.a(_w_5445),.q(_w_5446));
  bfr _b_11736(.a(_w_13638),.q(_w_13639));
  bfr _b_5261(.a(_w_7163),.q(_w_7164));
  bfr _b_13006(.a(_w_14908),.q(_w_14909));
  bfr _b_7431(.a(_w_9333),.q(_w_9334));
  bfr _b_7762(.a(_w_9664),.q(_w_9665));
  bfr _b_3533(.a(_w_5435),.q(_w_5436));
  bfr _b_3532(.a(_w_5434),.q(_w_5435));
  and_bi g590(.a(n588_0),.b(n589),.q(n590));
  bfr _b_4704(.a(_w_6606),.q(_w_6607));
  bfr _b_8001(.a(_w_9903),.q(_w_9904));
  bfr _b_3529(.a(_w_5431),.q(_w_5432));
  bfr _b_10210(.a(_w_12112),.q(_w_12113));
  bfr _b_3528(.a(_w_5430),.q(_w_5431));
  or_bb g1077(.a(n1075_0),.b(n1076_0),.q(n1077));
  bfr _b_3525(.a(_w_5427),.q(_w_5428));
  bfr _b_5457(.a(_w_7359),.q(_w_7360));
  bfr _b_3523(.a(_w_5425),.q(_w_5426));
  bfr _b_3521(.a(_w_5423),.q(_w_5424));
  bfr _b_11065(.a(_w_12967),.q(_w_12968));
  and_bi g1069(.a(n980_1),.b(n983_1),.q(n1069));
  bfr _b_5228(.a(_w_7130),.q(_w_7131));
  bfr _b_3520(.a(_w_5422),.q(_w_5423));
  bfr _b_3834(.a(_w_5736),.q(_w_5737));
  bfr _b_3680(.a(_w_5582),.q(_w_5583));
  bfr _b_6236(.a(_w_8138),.q(n424_1));
  bfr _b_3516(.a(_w_5418),.q(_w_5419));
  spl2 g1186_s_0(.a(n1186),.q0(n1186_0),.q1(n1186_1));
  and_bi g1385(.a(n1291_1),.b(n1294_1),.q(n1385));
  bfr _b_3515(.a(_w_5417),.q(_w_5418));
  bfr _b_3514(.a(_w_5416),.q(_w_5417));
  spl2 g1193_s_0(.a(n1193),.q0(n1193_0),.q1(n1193_1));
  bfr _b_6538(.a(_w_8440),.q(_w_8441));
  bfr _b_10695(.a(_w_12597),.q(_w_12598));
  or_bb g1863(.a(n1861_0),.b(n1862),.q(n1863));
  bfr _b_3513(.a(_w_5415),.q(_w_5416));
  bfr _b_3512(.a(_w_5414),.q(_w_5415));
  bfr _b_4529(.a(_w_6431),.q(_w_6432));
  and_bi g1848(.a(n1847_0),.b(n1818_0),.q(n1848));
  bfr _b_6815(.a(_w_8717),.q(_w_8718));
  bfr _b_3507(.a(_w_5409),.q(_w_5410));
  bfr _b_3506(.a(_w_5408),.q(_w_5409));
  bfr _b_4743(.a(_w_6645),.q(_w_6646));
  bfr _b_13555(.a(_w_15457),.q(_w_15458));
  bfr _b_11390(.a(_w_13292),.q(_w_13293));
  bfr _b_11114(.a(_w_13016),.q(_w_13017));
  spl2 g1110_s_0(.a(n1110),.q0(n1110_0),.q1(n1110_1));
  bfr _b_5622(.a(_w_7524),.q(_w_7525));
  spl2 g1856_s_0(.a(n1856),.q0(n1856_0),.q1(n1856_1));
  bfr _b_10493(.a(_w_12395),.q(n1893));
  bfr _b_3510(.a(_w_5412),.q(_w_5413));
  bfr _b_3502(.a(_w_5404),.q(_w_5405));
  bfr _b_11420(.a(_w_13322),.q(_w_13323));
  bfr _b_3500(.a(_w_5402),.q(_w_5403));
  bfr _b_9867(.a(_w_11769),.q(_w_11770));
  bfr _b_3496(.a(_w_5398),.q(_w_5399));
  bfr _b_7566(.a(_w_9468),.q(_w_9469));
  bfr _b_11063(.a(_w_12965),.q(_w_12966));
  spl4L N103_s_0(.a(_w_15525),.q0(N103_0),.q1(_w_6886),.q2(_w_6910),.q3(_w_6966));
  bfr _b_4625(.a(_w_6527),.q(_w_6528));
  and_bi g1204(.a(n1181_1),.b(n1202_1),.q(_w_13000));
  bfr _b_3491(.a(_w_5393),.q(_w_5394));
  bfr _b_3489(.a(_w_5391),.q(_w_5392));
  and_bi g580(.a(n530_1),.b(n578_1),.q(_w_13751));
  bfr _b_8815(.a(_w_10717),.q(_w_10718));
  bfr _b_3478(.a(_w_5380),.q(_w_5381));
  bfr _b_12795(.a(_w_14697),.q(_w_14698));
  bfr _b_3710(.a(_w_5612),.q(_w_5613));
  and_bi g499(.a(n498_0),.b(n442_0),.q(n499));
  bfr _b_6883(.a(_w_8785),.q(_w_8786));
  bfr _b_14300(.a(_w_16202),.q(_w_16203));
  bfr _b_10764(.a(_w_12666),.q(_w_12667));
  bfr _b_3476(.a(_w_5378),.q(_w_5379));
  bfr _b_7391(.a(_w_9293),.q(_w_9294));
  bfr _b_8398(.a(_w_10300),.q(_w_10301));
  bfr _b_8525(.a(_w_10427),.q(_w_10428));
  bfr _b_5355(.a(_w_7257),.q(_w_7258));
  bfr _b_10177(.a(_w_12079),.q(n1810));
  bfr _b_11446(.a(_w_13348),.q(_w_13349));
  bfr _b_3469(.a(_w_5371),.q(_w_5372));
  spl2 g570_s_0(.a(n570),.q0(n570_0),.q1(_w_13869));
  bfr _b_13046(.a(_w_14948),.q(_w_14949));
  bfr _b_3546(.a(_w_5448),.q(_w_5449));
  and_bi g1396(.a(n1381_1),.b(n1394_1),.q(_w_12216));
  bfr _b_3466(.a(_w_5368),.q(_w_5369));
  and_bb g1856(.a(N256_7),.b(N494_19),.q(_w_14674));
  bfr _b_13644(.a(_w_15546),.q(_w_15547));
  bfr _b_4259(.a(_w_6161),.q(_w_6162));
  bfr _b_3463(.a(_w_5365),.q(_w_5366));
  bfr _b_5427(.a(_w_7329),.q(_w_7330));
  bfr _b_3462(.a(_w_5364),.q(_w_5365));
  bfr _b_3453(.a(_w_5355),.q(_w_5356));
  bfr _b_9987(.a(_w_11889),.q(_w_11890));
  bfr _b_4561(.a(_w_6463),.q(N154_6));
  spl2 g1567_s_0(.a(n1567),.q0(n1567_0),.q1(n1567_1));
  bfr _b_5275(.a(_w_7177),.q(_w_7178));
  bfr _b_3446(.a(_w_5348),.q(_w_5349));
  and_bb g1471(.a(N256_14),.b(N375_19),.q(_w_9141));
  spl2 g735_s_0(.a(n735),.q0(n735_0),.q1(n735_1));
  bfr _b_4815(.a(_w_6717),.q(_w_6718));
  bfr _b_3444(.a(_w_5346),.q(N52_15));
  bfr _b_4456(.a(_w_6358),.q(_w_6359));
  bfr _b_9559(.a(_w_11461),.q(_w_11462));
  bfr _b_3443(.a(_w_5345),.q(_w_5346));
  spl2 g1053_s_0(.a(n1053),.q0(n1053_0),.q1(n1053_1));
  bfr _b_5581(.a(_w_7483),.q(_w_7484));
  bfr _b_3438(.a(_w_5340),.q(_w_5341));
  and_bi g1317(.a(n1315_0),.b(n1316),.q(n1317));
  bfr _b_7815(.a(_w_9717),.q(_w_9718));
  bfr _b_3437(.a(_w_5339),.q(_w_5340));
  bfr _b_3432(.a(_w_5334),.q(N52_14));
  bfr _b_10950(.a(_w_12852),.q(_w_12853));
  bfr _b_4377(.a(_w_6279),.q(n863_1));
  bfr _b_13960(.a(_w_15862),.q(_w_15863));
  and_bi g176(.a(n174_0),.b(n175),.q(n176));
  bfr _b_6343(.a(_w_8245),.q(_w_8246));
  bfr _b_3429(.a(_w_5331),.q(_w_5332));
  bfr _b_5926(.a(_w_7828),.q(_w_7829));
  bfr _b_9007(.a(_w_10909),.q(n266));
  bfr _b_4298(.a(_w_6200),.q(_w_6201));
  bfr _b_3424(.a(_w_5326),.q(_w_5327));
  bfr _b_11886(.a(_w_13788),.q(_w_13789));
  spl2 g1214_s_0(.a(n1214),.q0(n1214_0),.q1(n1214_1));
  bfr _b_3420(.a(_w_5322),.q(N52_13));
  spl2 g225_s_0(.a(n225),.q0(n225_0),.q1(n225_1));
  bfr _b_4792(.a(_w_6694),.q(_w_6695));
  bfr _b_13654(.a(_w_15556),.q(_w_15557));
  bfr _b_3417(.a(_w_5319),.q(_w_5320));
  and_bi g1674(.a(n1653_1),.b(n1656_1),.q(n1674));
  bfr _b_14370(.a(_w_16272),.q(_w_16273));
  bfr _b_8598(.a(_w_10500),.q(_w_10501));
  bfr _b_5052(.a(_w_6954),.q(_w_6955));
  bfr _b_4129(.a(_w_6031),.q(_w_6032));
  spl2 g1012_s_0(.a(n1012),.q0(n1012_0),.q1(n1012_1));
  and_bb g78(.a(n57_1),.b(n77_0),.q(n78));
  spl2 g857_s_0(.a(n857),.q0(n857_0),.q1(_w_5307));
  bfr _b_4096(.a(_w_5998),.q(_w_5999));
  spl2 g1083_s_0(.a(n1083),.q0(n1083_0),.q1(_w_5311));
  bfr _b_13043(.a(_w_14945),.q(_w_14946));
  bfr _b_4011(.a(_w_5913),.q(_w_5914));
  bfr _b_9875(.a(_w_11777),.q(_w_11778));
  bfr _b_12478(.a(_w_14380),.q(_w_14381));
  spl4L N52_s_3(.a(N52_2),.q0(N52_12),.q1(_w_5315),.q2(_w_5323),.q3(_w_5335));
  bfr _b_7911(.a(_w_9813),.q(_w_9814));
  bfr _b_10787(.a(_w_12689),.q(_w_12690));
  bfr _b_6076(.a(_w_7978),.q(_w_7979));
  bfr _b_7848(.a(_w_9750),.q(_w_9751));
  bfr _b_9063(.a(_w_10965),.q(_w_10966));
  spl4L N52_s_0(.a(_w_16197),.q0(N52_0),.q1(_w_5371),.q2(_w_5395),.q3(_w_5451));
  spl2 g1079_s_0(.a(n1079),.q0(n1079_0),.q1(n1079_1));
  bfr _b_5415(.a(_w_7317),.q(_w_7318));
  bfr _b_10495(.a(_w_12397),.q(_w_12398));
  spl2 g1740_s_0(.a(n1740),.q0(n1740_0),.q1(n1740_1));
  bfr _b_13484(.a(_w_15386),.q(_w_15387));
  and_bi g426(.a(n424_0),.b(n425),.q(n426));
  spl2 g1558_s_0(.a(n1558),.q0(n1558_0),.q1(_w_5543));
  bfr _b_3558(.a(_w_5460),.q(_w_5461));
  and_bi g527(.a(n496_1),.b(n499_1),.q(n527));
  bfr _b_5883(.a(_w_7785),.q(_w_7786));
  bfr _b_8477(.a(_w_10379),.q(_w_10380));
  bfr _b_13348(.a(_w_15250),.q(_w_15251));
  bfr _b_4408(.a(_w_6310),.q(_w_6311));
  bfr _b_11628(.a(_w_13530),.q(_w_13531));
  bfr _b_6816(.a(_w_8718),.q(_w_8719));
  bfr _b_13011(.a(_w_14913),.q(_w_14914));
  bfr _b_7540(.a(_w_9442),.q(_w_9443));
  spl2 g923_s_0(.a(n923),.q0(n923_0),.q1(_w_5551));
  bfr _b_4741(.a(_w_6643),.q(_w_6644));
  spl2 g187_s_0(.a(n187),.q0(n187_0),.q1(n187_1));
  bfr _b_13969(.a(_w_15871),.q(_w_15872));
  bfr _b_12942(.a(_w_14844),.q(_w_14845));
  bfr _b_10707(.a(_w_12609),.q(_w_12610));
  bfr _b_4302(.a(_w_6204),.q(_w_6205));
  spl2 g1051_s_0(.a(n1051),.q0(n1051_0),.q1(n1051_1));
  and_bi g1153(.a(n1050_1),.b(n1151_1),.q(_w_12858));
  spl2 g1050_s_0(.a(n1050),.q0(n1050_0),.q1(n1050_1));
  spl2 g1036_s_0(.a(n1036),.q0(n1036_0),.q1(n1036_1));
  bfr _b_10482(.a(_w_12384),.q(_w_12385));
  bfr _b_8556(.a(_w_10458),.q(n306));
  and_bi g164(.a(n162_0),.b(n163),.q(n164));
  spl2 g1007_s_0(.a(n1007),.q0(n1007_0),.q1(n1007_1));
  spl2 g1003_s_0(.a(n1003),.q0(n1003_0),.q1(n1003_1));
  spl2 g724_s_0(.a(n724),.q0(n724_0),.q1(n724_1));
  bfr _b_4064(.a(_w_5966),.q(_w_5967));
  bfr _b_6517(.a(_w_8419),.q(_w_8420));
  bfr _b_6903(.a(_w_8805),.q(_w_8806));
  bfr _b_6575(.a(_w_8477),.q(_w_8478));
  or_bb g979(.a(n977_0),.b(n978),.q(n979));
  and_bi g970(.a(n968_0),.b(n969),.q(n970));
  spl2 g455_s_0(.a(n455),.q0(n455_0),.q1(n455_1));
  spl4L N256_s_0(.a(_w_15534),.q0(_w_5699),.q1(_w_5749),.q2(_w_5815),.q3(N256_3));
  spl2 g1188_s_0(.a(n1188),.q0(n1188_0),.q1(_w_5820));
  bfr _b_5416(.a(_w_7318),.q(N86_1));
  bfr _b_3974(.a(_w_5876),.q(_w_5877));
  spl2 g985_s_0(.a(n985),.q0(n985_0),.q1(n985_1));
  spl2 g980_s_0(.a(n980),.q0(n980_0),.q1(_w_5827));
  and_bi g769(.a(n768_0),.b(n728_0),.q(n769));
  spl2 g979_s_0(.a(n979),.q0(n979_0),.q1(n979_1));
  spl2 g736_s_0(.a(n736),.q0(n736_0),.q1(n736_1));
  bfr _b_12902(.a(_w_14804),.q(_w_14805));
  spl2 g883_s_0(.a(n883),.q0(n883_0),.q1(n883_1));
  bfr _b_7571(.a(_w_9473),.q(_w_9474));
  spl2 g949_s_0(.a(n949),.q0(n949_0),.q1(n949_1));
  spl2 g974_s_0(.a(n974),.q0(n974_0),.q1(_w_5831));
  and_bi g800(.a(n718_1),.b(n798_1),.q(_w_12616));
  spl2 g833_s_0(.a(n833),.q0(n833_0),.q1(n833_1));
  bfr _b_11843(.a(_w_13745),.q(N1_3));
  spl2 g1596_s_0(.a(n1596),.q0(n1596_0),.q1(n1596_1));
  spl2 g739_s_0(.a(n739),.q0(n739_0),.q1(_w_5835));
  bfr _b_8745(.a(_w_10647),.q(_w_10648));
  spl2 g964_s_0(.a(n964),.q0(n964_0),.q1(n964_1));
  spl2 g937_s_0(.a(n937),.q0(n937_0),.q1(n937_1));
  bfr _b_4805(.a(_w_6707),.q(_w_6708));
  bfr _b_4596(.a(_w_6498),.q(_w_6499));
  bfr _b_12548(.a(_w_14450),.q(_w_14451));
  bfr _b_7765(.a(_w_9667),.q(_w_9668));
  bfr _b_4553(.a(_w_6455),.q(_w_6456));
  spl2 g932_s_0(.a(n932),.q0(n932_0),.q1(n932_1));
  bfr _b_4592(.a(_w_6494),.q(_w_6495));
  spl2 g1197_s_0(.a(n1197),.q0(n1197_0),.q1(n1197_1));
  spl3L g78_s_0(.a(n78),.q0(n78_0),.q1(_w_5837),.q2(_w_5839));
  spl2 g1466_s_0(.a(n1466),.q0(n1466_0),.q1(n1466_1));
  bfr _b_4765(.a(_w_6667),.q(_w_6668));
  bfr _b_8858(.a(_w_10760),.q(_w_10761));
  bfr _b_4143(.a(_w_6045),.q(_w_6046));
  and_bi g816(.a(n814_0),.b(n815),.q(n816));
  bfr _b_11438(.a(_w_13340),.q(_w_13341));
  spl2 g941_s_0(.a(n941),.q0(n941_0),.q1(n941_1));
  spl2 g1808_s_0(.a(n1808),.q0(n1808_0),.q1(n1808_1));
  spl2 g938_s_0(.a(n938),.q0(n938_0),.q1(n938_1));
  spl2 g1665_s_0(.a(n1665),.q0(n1665_0),.q1(_w_15002));
  spl2 g929_s_0(.a(n929),.q0(n929_0),.q1(_w_5841));
  spl2 g654_s_0(.a(n654),.q0(n654_0),.q1(n654_1));
  spl2 g1116_s_0(.a(n1116),.q0(n1116_0),.q1(n1116_1));
  and_bb g72(.a(N1_8),.b(N341_4),.q(n72));
  bfr _b_8069(.a(_w_9971),.q(_w_9972));
  bfr _b_4945(.a(_w_6847),.q(_w_6848));
  bfr _b_4153(.a(_w_6055),.q(_w_6056));
  bfr _b_6066(.a(_w_7968),.q(_w_7969));
  bfr _b_8042(.a(_w_9944),.q(_w_9945));
  spl2 g919_s_0(.a(n919),.q0(n919_0),.q1(n919_1));
  bfr _b_8087(.a(_w_9989),.q(_w_9990));
  bfr _b_3686(.a(_w_5588),.q(_w_5589));
  spl2 g460_s_0(.a(n460),.q0(n460_0),.q1(_w_13858));
  bfr _b_3712(.a(_w_5614),.q(_w_5615));
  spl2 g1635_s_0(.a(n1635),.q0(n1635_0),.q1(_w_5547));
  bfr _b_5420(.a(_w_7322),.q(_w_7323));
  spl2 g517_s_0(.a(n517),.q0(n517_0),.q1(n517_1));
  spl4L N239_s_2(.a(N239_1),.q0(N239_8),.q1(N239_9),.q2(N239_10),.q3(_w_5885));
  and_bi g1318(.a(n1317_0),.b(n1280_0),.q(n1318));
  spl4L N239_s_0(.a(_w_15533),.q0(N239_0),.q1(_w_5913),.q2(_w_5937),.q3(_w_5993));
  spl3L g1046_s_0(.a(n1046),.q0(n1046_0),.q1(n1046_1),.q2(n1046_2));
  bfr _b_9639(.a(_w_11541),.q(_w_11542));
  bfr _b_11998(.a(_w_13900),.q(n538));
  bfr _b_8015(.a(_w_9917),.q(_w_9918));
  bfr _b_3419(.a(_w_5321),.q(_w_5322));
  bfr _b_13460(.a(_w_15362),.q(_w_15363));
  bfr _b_5331(.a(_w_7233),.q(_w_7234));
  spl2 g1779_s_0(.a(n1779),.q0(n1779_0),.q1(n1779_1));
  bfr _b_5762(.a(_w_7664),.q(_w_7665));
  spl2 g884_s_0(.a(n884),.q0(n884_0),.q1(n884_1));
  bfr _b_4237(.a(_w_6139),.q(_w_6140));
  bfr _b_6300(.a(_w_8202),.q(n1084));
  spl2 g372_s_0(.a(n372),.q0(n372_0),.q1(n372_1));
  and_bb g716(.a(N35_16),.b(N477_6),.q(n716));
  spl2 g943_s_0(.a(n943),.q0(n943_0),.q1(n943_1));
  bfr _b_4891(.a(_w_6793),.q(_w_6794));
  bfr _b_12251(.a(_w_14153),.q(_w_14154));
  spl2 g258_s_0(.a(n258),.q0(n258_0),.q1(n258_1));
  spl2 g875_s_0(.a(n875),.q0(n875_0),.q1(_w_6081));
  bfr _b_7340(.a(_w_9242),.q(n1181));
  spl2 g1587_s_0(.a(n1587),.q0(n1587_0),.q1(n1587_1));
  bfr _b_13406(.a(_w_15308),.q(n496_1));
  bfr _b_5652(.a(_w_7554),.q(_w_7555));
  spl2 g862_s_0(.a(n862),.q0(n862_0),.q1(n862_1));
  bfr _b_7535(.a(_w_9437),.q(_w_9438));
  bfr _b_3785(.a(_w_5687),.q(_w_5688));
  bfr _b_4763(.a(_w_6665),.q(N1_15));
  spl2 g765_s_0(.a(n765),.q0(n765_0),.q1(n765_1));
  spl2 g844_s_0(.a(n844),.q0(n844_0),.q1(n844_1));
  and_bi g609(.a(n608_0),.b(n520_0),.q(n609));
  bfr _b_8135(.a(_w_10037),.q(_w_10038));
  spl2 g1054_s_0(.a(n1054),.q0(n1054_0),.q1(n1054_1));
  bfr _b_9038(.a(_w_10940),.q(_w_10941));
  bfr _b_4137(.a(_w_6039),.q(_w_6040));
  bfr _b_8116(.a(_w_10018),.q(_w_10019));
  bfr _b_3471(.a(_w_5373),.q(_w_5374));
  bfr _b_3445(.a(_w_5347),.q(_w_5348));
  spl2 g1250_s_0(.a(n1250),.q0(n1250_0),.q1(n1250_1));
  spl2 g702_s_0(.a(n702),.q0(n702_0),.q1(n702_1));
  bfr _b_7652(.a(_w_9554),.q(_w_9555));
  and_bi g464(.a(n454_1),.b(n462_1),.q(_w_12849));
  bfr _b_10331(.a(_w_12233),.q(_w_12234));
  bfr _b_9684(.a(_w_11586),.q(_w_11587));
  bfr _b_3911(.a(_w_5813),.q(_w_5814));
  bfr _b_13038(.a(_w_14940),.q(_w_14941));
  spl2 g828_s_0(.a(n828),.q0(n828_0),.q1(n828_1));
  and_bi g305(.a(n250_1),.b(n253_1),.q(n305));
  and_bb g1340(.a(n1273_1),.b(n1338_1),.q(_w_15019));
  bfr _b_8490(.a(_w_10392),.q(_w_10393));
  bfr _b_4009(.a(_w_5911),.q(_w_5912));
  bfr _b_11728(.a(_w_13630),.q(_w_13631));
  bfr _b_4816(.a(_w_6718),.q(_w_6719));
  bfr _b_12882(.a(_w_14784),.q(_w_14785));
  bfr _b_3952(.a(_w_5854),.q(_w_5855));
  spl2 g1735_s_0(.a(n1735),.q0(n1735_0),.q1(n1735_1));
  bfr _b_12611(.a(_w_14513),.q(_w_14514));
  bfr _b_4470(.a(_w_6372),.q(_w_6373));
  bfr _b_5650(.a(_w_7552),.q(_w_7553));
  spl2 g393_s_0(.a(n393),.q0(n393_0),.q1(n393_1));
  bfr _b_4576(.a(_w_6478),.q(_w_6479));
  bfr _b_3628(.a(_w_5530),.q(_w_5531));
  spl2 g1025_s_0(.a(n1025),.q0(n1025_0),.q1(n1025_1));
  bfr _b_4041(.a(_w_5943),.q(_w_5944));
  bfr _b_10516(.a(_w_12418),.q(_w_12419));
  bfr _b_7088(.a(_w_8990),.q(_w_8991));
  spl2 g995_s_0(.a(n995),.q0(n995_0),.q1(n995_1));
  bfr _b_10358(.a(_w_12260),.q(_w_12261));
  bfr _b_3981(.a(_w_5883),.q(_w_5884));
  bfr _b_7831(.a(_w_9733),.q(_w_9734));
  bfr _b_8165(.a(_w_10067),.q(_w_10068));
  bfr _b_12364(.a(_w_14266),.q(_w_14267));
  spl2 g217_s_0(.a(n217),.q0(n217_0),.q1(n217_1));
  bfr _b_3999(.a(_w_5901),.q(_w_5902));
  bfr _b_9488(.a(_w_11390),.q(_w_11391));
  spl2 g852_s_0(.a(n852),.q0(n852_0),.q1(_w_6085));
  bfr _b_4031(.a(_w_5933),.q(_w_5934));
  bfr _b_13919(.a(_w_15821),.q(_w_15822));
  bfr _b_4447(.a(_w_6349),.q(n1716_1));
  bfr _b_7258(.a(_w_9160),.q(n1471));
  bfr _b_4396(.a(_w_6298),.q(_w_6299));
  spl2 g440_s_0(.a(n440),.q0(n440_0),.q1(n440_1));
  bfr _b_14189(.a(_w_16091),.q(_w_16092));
  bfr _b_13235(.a(_w_15137),.q(_w_15138));
  spl2 g916_s_0(.a(n916),.q0(n916_0),.q1(n916_1));
  bfr _b_12591(.a(_w_14493),.q(_w_14494));
  bfr _b_7690(.a(_w_9592),.q(_w_9593));
  spl2 g802_s_0(.a(n802),.q0(n802_0),.q1(_w_6089));
  bfr _b_5226(.a(_w_7128),.q(_w_7129));
  bfr _b_5818(.a(_w_7720),.q(_w_7721));
  spl2 g1550_s_0(.a(n1550),.q0(n1550_0),.q1(n1550_1));
  and_bi g1816(.a(n1777_1),.b(n1814_1),.q(_w_13940));
  spl4L N171_s_3(.a(N171_2),.q0(N171_12),.q1(_w_6093),.q2(_w_6101),.q3(_w_6113));
  spl2 g1398_s_0(.a(n1398),.q0(n1398_0),.q1(_w_11396));
  spl4L N171_s_2(.a(N171_1),.q0(N171_8),.q1(N171_9),.q2(N171_10),.q3(_w_6125));
  spl2 g566_s_0(.a(n566),.q0(n566_0),.q1(n566_1));
  bfr _b_14219(.a(_w_16121),.q(_w_16122));
  bfr _b_9850(.a(_w_11752),.q(_w_11753));
  spl4L N171_s_1(.a(N171_0),.q0(N171_4),.q1(N171_5),.q2(_w_6149),.q3(_w_6151));
  spl2 g795_s_0(.a(n795),.q0(n795_0),.q1(n795_1));
  bfr _b_13347(.a(_w_15249),.q(_w_15250));
  bfr _b_12214(.a(_w_14116),.q(n1702));
  spl2 g1543_s_0(.a(n1543),.q0(n1543_0),.q1(n1543_1));
  spl2 g439_s_0(.a(n439),.q0(n439_0),.q1(n439_1));
  bfr _b_4965(.a(_w_6867),.q(_w_6868));
  bfr _b_11957(.a(_w_13859),.q(_w_13860));
  bfr _b_4135(.a(_w_6037),.q(_w_6038));
  bfr _b_8409(.a(_w_10311),.q(_w_10312));
  spl2 g792_s_0(.a(n792),.q0(n792_0),.q1(n792_1));
  bfr _b_4534(.a(_w_6436),.q(_w_6437));
  spl2 g1783_s_0(.a(n1783),.q0(n1783_0),.q1(n1783_1));
  bfr _b_6103(.a(_w_8005),.q(_w_8006));
  bfr _b_12668(.a(_w_14570),.q(n1760));
  bfr _b_10041(.a(_w_11943),.q(_w_11944));
  bfr _b_6768(.a(_w_8670),.q(_w_8671));
  bfr _b_3650(.a(_w_5552),.q(_w_5553));
  spl2 g780_s_0(.a(n780),.q0(n780_0),.q1(n780_1));
  bfr _b_11315(.a(_w_13217),.q(_w_13218));
  bfr _b_6445(.a(_w_8347),.q(_w_8348));
  spl2 g1324_s_0(.a(n1324),.q0(n1324_0),.q1(n1324_1));
  bfr _b_6025(.a(_w_7927),.q(N188_15));
  bfr _b_8445(.a(_w_10347),.q(_w_10348));
  and_bb g969(.a(n961_1),.b(n967_1),.q(_w_9208));
  bfr _b_11191(.a(_w_13093),.q(_w_13094));
  spl2 g756_s_0(.a(n756),.q0(n756_0),.q1(n756_1));
  spl2 g822_s_0(.a(n822),.q0(n822_0),.q1(n822_1));
  bfr _b_13797(.a(_w_15699),.q(_w_15700));
  or_bb g44(.a(n33_1),.b(n43_0),.q(_w_10622));
  bfr _b_4138(.a(_w_6040),.q(_w_6041));
  spl2 g824_s_0(.a(n824),.q0(n824_0),.q1(n824_1));
  spl2 g1010_s_0(.a(n1010),.q0(n1010_0),.q1(_w_6161));
  bfr _b_8075(.a(_w_9977),.q(_w_9978));
  spl2 g1348_s_0(.a(n1348),.q0(n1348_0),.q1(n1348_1));
  and_bi g642(.a(n640_0),.b(n641),.q(n642));
  spl2 g634_s_0(.a(n634),.q0(n634_0),.q1(n634_1));
  bfr _b_11414(.a(_w_13316),.q(_w_13317));
  bfr _b_10708(.a(_w_12610),.q(_w_12611));
  bfr _b_8456(.a(_w_10358),.q(_w_10359));
  bfr _b_7890(.a(_w_9792),.q(_w_9793));
  or_bb g1764(.a(n1762_0),.b(n1763),.q(n1764));
  bfr _b_5599(.a(_w_7501),.q(_w_7502));
  spl2 g731_s_0(.a(n731),.q0(n731_0),.q1(n731_1));
  bfr _b_9218(.a(_w_11120),.q(_w_11121));
  bfr _b_9832(.a(_w_11734),.q(_w_11735));
  bfr _b_4319(.a(_w_6221),.q(_w_6222));
  spl2 g1065_s_0(.a(n1065),.q0(n1065_0),.q1(n1065_1));
  bfr _b_7063(.a(_w_8965),.q(_w_8966));
  spl2 g726_s_0(.a(n726),.q0(n726_0),.q1(n726_1));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(_w_6173));
  bfr _b_11382(.a(_w_13284),.q(_w_13285));
  bfr _b_7525(.a(_w_9427),.q(_w_9428));
  spl2 g748_s_0(.a(n748),.q0(n748_0),.q1(_w_6177));
  bfr _b_3793(.a(_w_5695),.q(_w_5696));
  spl4L N86_s_2(.a(N86_1),.q0(N86_8),.q1(N86_9),.q2(N86_10),.q3(_w_7271));
  and_bi g1898(.a(n1895_0),.b(n1897),.q(n1898));
  bfr _b_7942(.a(_w_9844),.q(_w_9845));
  spl2 g718_s_0(.a(n718),.q0(n718_0),.q1(n718_1));
  bfr _b_10004(.a(_w_11906),.q(_w_11907));
  bfr _b_4606(.a(_w_6508),.q(_w_6509));
  bfr _b_7387(.a(_w_9289),.q(n1738));
  spl2 g713_s_0(.a(n713),.q0(n713_0),.q1(n713_1));
  bfr _b_6294(.a(_w_8196),.q(_w_8197));
  bfr _b_4086(.a(_w_5988),.q(_w_5989));
  bfr _b_7377(.a(_w_9279),.q(_w_9280));
  spl2 g706_s_0(.a(n706),.q0(n706_0),.q1(_w_6188));
  bfr _b_4918(.a(_w_6820),.q(_w_6821));
  spl4L N86_s_1(.a(N86_0),.q0(N86_4),.q1(N86_5),.q2(_w_12859),.q3(_w_12861));
  spl2 g590_s_0(.a(n590),.q0(n590_0),.q1(n590_1));
  bfr _b_13493(.a(_w_15395),.q(_w_15396));
  bfr _b_4560(.a(_w_6462),.q(_w_6463));
  bfr _b_3730(.a(_w_5632),.q(_w_5633));
  spl2 g1166_s_0(.a(n1166),.q0(n1166_0),.q1(n1166_1));
  bfr _b_12638(.a(_w_14540),.q(n1807));
  bfr _b_12470(.a(_w_14372),.q(_w_14373));
  bfr _b_7806(.a(_w_9708),.q(_w_9709));
  spl2 g688_s_0(.a(n688),.q0(n688_0),.q1(_w_6196));
  spl2 g60_s_0(.a(n60),.q0(n60_0),.q1(_w_14277));
  spl2 g59_s_0(.a(n59),.q0(n59_0),.q1(n59_1));
  spl2 g684_s_0(.a(n684),.q0(n684_0),.q1(n684_1));
  bfr _b_8439(.a(_w_10341),.q(_w_10342));
  spl2 g1675_s_0(.a(n1675),.q0(n1675_0),.q1(n1675_1));
  spl2 g1796_s_0(.a(n1796),.q0(n1796_0),.q1(n1796_1));
  spl2 g1668_s_0(.a(n1668),.q0(n1668_0),.q1(n1668_1));
  bfr _b_6655(.a(_w_8557),.q(_w_8558));
  bfr _b_13321(.a(_w_15223),.q(_w_15224));
  bfr _b_7694(.a(_w_9596),.q(_w_9597));
  bfr _b_12432(.a(_w_14334),.q(_w_14335));
  spl2 g681_s_0(.a(n681),.q0(n681_0),.q1(n681_1));
  spl2 g676_s_0(.a(n676),.q0(n676_0),.q1(_w_6200));
  bfr _b_3499(.a(_w_5401),.q(_w_5402));
  bfr _b_12894(.a(_w_14796),.q(_w_14797));
  or_bb g699(.a(n697_0),.b(n698),.q(n699));
  spl2 g675_s_0(.a(n675),.q0(n675_0),.q1(n675_1));
  spl4L N409_s_3(.a(N409_2),.q0(N409_12),.q1(N409_13),.q2(N409_14),.q3(N409_15));
  bfr _b_5909(.a(_w_7811),.q(_w_7812));
  bfr _b_7419(.a(_w_9321),.q(_w_9322));
  bfr _b_7924(.a(_w_9826),.q(_w_9827));
  bfr _b_3794(.a(_w_5696),.q(_w_5697));
  bfr _b_7846(.a(_w_9748),.q(_w_9749));
  or_bb g778(.a(n725_0),.b(n777_0),.q(n778));
  bfr _b_12143(.a(_w_14045),.q(_w_14046));
  spl2 g672_s_0(.a(n672),.q0(n672_0),.q1(n672_1));
  spl2 g144_s_0(.a(n144),.q0(n144_0),.q1(n144_1));
  spl2 g1377_s_0(.a(n1377),.q0(n1377_0),.q1(n1377_1));
  spl2 g1842_s_0(.a(n1842),.q0(n1842_0),.q1(n1842_1));
  bfr _b_4334(.a(_w_6236),.q(_w_6237));
  bfr _b_4708(.a(_w_6610),.q(_w_6611));
  spl4L N477_s_0(.a(_w_15930),.q0(N477_0),.q1(N477_1),.q2(N477_2),.q3(N477_3));
  bfr _b_4050(.a(_w_5952),.q(_w_5953));
  and_bi g1182(.a(n1089_1),.b(n1092_1),.q(n1182));
  and_bb g981(.a(n957_1),.b(n979_1),.q(_w_12396));
  bfr _b_5759(.a(_w_7661),.q(_w_7662));
  spl2 g670_s_0(.a(n670),.q0(n670_0),.q1(_w_6204));
  bfr _b_13700(.a(_w_15602),.q(_w_15603));
  spl2 g1895_s_0(.a(n1895),.q0(n1895_0),.q1(_w_14939));
  spl2 g669_s_0(.a(n669),.q0(n669_0),.q1(n669_1));
  bfr _b_13269(.a(_w_15171),.q(_w_15172));
  bfr _b_11299(.a(_w_13201),.q(_w_13202));
  bfr _b_10118(.a(_w_12020),.q(_w_12021));
  bfr _b_6923(.a(_w_8825),.q(_w_8826));
  bfr _b_8776(.a(_w_10678),.q(_w_10679));
  bfr _b_3642(.a(_w_5544),.q(_w_5545));
  spl2 g715_s_0(.a(n715),.q0(n715_0),.q1(n715_1));
  spl2 g667_s_0(.a(n667),.q0(n667_0),.q1(n667_1));
  bfr _b_9508(.a(_w_11410),.q(_w_11411));
  bfr _b_12555(.a(_w_14457),.q(_w_14458));
  bfr _b_12223(.a(_w_14125),.q(_w_14126));
  bfr _b_4747(.a(_w_6649),.q(_w_6650));
  bfr _b_10648(.a(_w_12550),.q(_w_12551));
  bfr _b_6155(.a(_w_8057),.q(_w_8058));
  bfr _b_13958(.a(_w_15860),.q(_w_15792));
  bfr _b_12197(.a(_w_14099),.q(_w_14100));
  spl2 g664_s_0(.a(n664),.q0(n664_0),.q1(_w_6208));
  spl2 g1535_s_0(.a(n1535),.q0(n1535_0),.q1(n1535_1));
  spl4L N120_s_4(.a(N120_3),.q0(N120_16),.q1(N120_17),.q2(N120_18),.q3(N120_19));
  and_bb g1322(.a(n1279_1),.b(n1320_1),.q(_w_8950));
  bfr _b_11625(.a(_w_13527),.q(_w_13528));
  and_bi g1700(.a(n1698_0),.b(n1699),.q(n1700));
  spl4L N120_s_3(.a(N120_2),.q0(N120_12),.q1(_w_6212),.q2(_w_6220),.q3(_w_6232));
  bfr _b_5572(.a(_w_7474),.q(n1800_1));
  bfr _b_8777(.a(_w_10679),.q(_w_10680));
  bfr _b_3673(.a(_w_5575),.q(_w_5576));
  bfr _b_10577(.a(_w_12479),.q(_w_12480));
  spl4L N120_s_1(.a(N120_0),.q0(N120_4),.q1(N120_5),.q2(_w_6268),.q3(_w_6270));
  spl2 g655_s_0(.a(n655),.q0(n655_0),.q1(n655_1));
  bfr _b_9546(.a(_w_11448),.q(_w_11449));
  spl2 g1470_s_0(.a(n1470),.q0(n1470_0),.q1(n1470_1));
  bfr _b_11186(.a(_w_13088),.q(_w_13089));
  bfr _b_4598(.a(_w_6500),.q(_w_6501));
  or_bb g286(.a(n233_0),.b(n285_0),.q(n286));
  bfr _b_3423(.a(_w_5325),.q(_w_5326));
  spl2 g640_s_0(.a(n640),.q0(n640_0),.q1(_w_6272));
  spl2 g639_s_0(.a(n639),.q0(n639_0),.q1(n639_1));
  bfr _b_8073(.a(_w_9975),.q(_w_9976));
  bfr _b_11356(.a(_w_13258),.q(_w_13259));
  spl2 g1027_s_0(.a(n1027),.q0(n1027_0),.q1(n1027_1));
  spl2 g957_s_0(.a(n957),.q0(n957_0),.q1(n957_1));
  spl2 g633_s_0(.a(n633),.q0(n633_0),.q1(n633_1));
  spl2 g651_s_0(.a(n651),.q0(n651_0),.q1(n651_1));
  and_bi g228(.a(n226_0),.b(n227),.q(n228));
  bfr _b_5555(.a(_w_7457),.q(_w_7458));
  spl2 g632_s_0(.a(n632),.q0(n632_0),.q1(n632_1));
  spl2 g532_s_0(.a(n532),.q0(n532_0),.q1(n532_1));
  spl2 g630_s_0(.a(n630),.q0(n630_0),.q1(n630_1));
  bfr _b_8806(.a(_w_10708),.q(_w_10709));
  and_bi g1376(.a(n1315_1),.b(n1318_1),.q(n1376));
  bfr _b_10352(.a(_w_12254),.q(_w_12255));
  bfr _b_5752(.a(_w_7654),.q(_w_7655));
  spl2 g620_s_0(.a(n620),.q0(n620_0),.q1(n620_1));
  bfr _b_4352(.a(_w_6254),.q(_w_6255));
  bfr _b_5655(.a(_w_7557),.q(_w_7558));
  spl2 g617_s_0(.a(n617),.q0(n617_0),.q1(n617_1));
  bfr _b_13301(.a(_w_15203),.q(_w_15204));
  spl2 g616_s_0(.a(n616),.q0(n616_0),.q1(n616_1));
  bfr _b_7684(.a(_w_9586),.q(_w_9587));
  spl2 g615_s_0(.a(n615),.q0(n615_0),.q1(n615_1));
  bfr _b_4067(.a(_w_5969),.q(_w_5970));
  bfr _b_12730(.a(_w_14632),.q(_w_14633));
  and_bi g314(.a(n312_0),.b(n313),.q(n314));
  bfr _b_4364(.a(_w_6266),.q(_w_6267));
  bfr _b_7800(.a(_w_9702),.q(_w_9703));
  spl2 g1202_s_0(.a(n1202),.q0(n1202_0),.q1(n1202_1));
  bfr _b_5130(.a(_w_7032),.q(_w_7033));
  spl2 g608_s_0(.a(n608),.q0(n608_0),.q1(n608_1));
  bfr _b_9762(.a(_w_11664),.q(_w_11665));
  or_bb g849(.a(n737_1),.b(n848_0),.q(n849));
  spl2 g237_s_0(.a(n237),.q0(n237_0),.q1(n237_1));
  bfr _b_5062(.a(_w_6964),.q(_w_6965));
  bfr _b_8753(.a(_w_10655),.q(_w_10656));
  spl2 g1563_s_0(.a(n1563),.q0(n1563_0),.q1(n1563_1));
  spl2 g588_s_0(.a(n588),.q0(n588_0),.q1(_w_6288));
  bfr _b_11400(.a(_w_13302),.q(_w_13303));
  spl2 g587_s_0(.a(n587),.q0(n587_0),.q1(n587_1));
  bfr _b_5237(.a(_w_7139),.q(_w_7140));
  spl2 g931_s_0(.a(n931),.q0(n931_0),.q1(n931_1));
  bfr _b_11796(.a(_w_13698),.q(_w_13699));
  bfr _b_4467(.a(_w_6369),.q(n118_1));
  bfr _b_6041(.a(_w_7943),.q(_w_7944));
  bfr _b_6990(.a(_w_8892),.q(_w_8893));
  bfr _b_6838(.a(_w_8740),.q(_w_8741));
  bfr _b_7189(.a(_w_9091),.q(_w_9092));
  bfr _b_8656(.a(_w_10558),.q(N4591));
  bfr _b_3717(.a(_w_5619),.q(_w_5620));
  spl2 g1076_s_0(.a(n1076),.q0(n1076_0),.q1(n1076_1));
  bfr _b_8682(.a(_w_10584),.q(_w_10585));
  spl2 g72_s_0(.a(n72),.q0(n72_0),.q1(n72_1));
  bfr _b_13314(.a(_w_15216),.q(_w_15217));
  spl2 g1573_s_0(.a(n1573),.q0(n1573_0),.q1(n1573_1));
  bfr _b_4454(.a(_w_6356),.q(_w_6357));
  spl2 g759_s_0(.a(n759),.q0(n759_0),.q1(n759_1));
  bfr _b_4750(.a(_w_6652),.q(_w_6653));
  spl2 g823_s_0(.a(n823),.q0(n823_0),.q1(n823_1));
  bfr _b_10081(.a(_w_11983),.q(_w_11984));
  bfr _b_9349(.a(_w_11251),.q(N35_1));
  or_bb g928(.a(n926_0),.b(n927),.q(n928));
  spl2 g306_s_0(.a(n306),.q0(n306_0),.q1(n306_1));
  spl2 g835_s_0(.a(n835),.q0(n835_0),.q1(n835_1));
  bfr _b_8457(.a(_w_10359),.q(_w_10360));
  bfr _b_11059(.a(_w_12961),.q(_w_12962));
  bfr _b_3938(.a(_w_5840),.q(n78_2));
  bfr _b_7551(.a(_w_9453),.q(_w_9454));
  spl2 g564_s_0(.a(n564),.q0(n564_0),.q1(_w_6300));
  bfr _b_10066(.a(_w_11968),.q(_w_11969));
  spl2 g554_s_0(.a(n554),.q0(n554_0),.q1(n554_1));
  bfr _b_10481(.a(_w_12383),.q(_w_12384));
  spl2 g877_s_0(.a(n877),.q0(n877_0),.q1(n877_1));
  spl2 g629_s_0(.a(n629),.q0(n629_0),.q1(n629_1));
  bfr _b_7423(.a(_w_9325),.q(_w_9326));
  spl2 g708_s_0(.a(n708),.q0(n708_0),.q1(n708_1));
  bfr _b_4241(.a(_w_6143),.q(_w_6144));
  bfr _b_4220(.a(_w_6122),.q(_w_6123));
  bfr _b_13742(.a(_w_15644),.q(_w_15645));
  bfr _b_6929(.a(_w_8831),.q(_w_8832));
  bfr _b_4843(.a(_w_6745),.q(_w_6746));
  spl2 g541_s_0(.a(n541),.q0(n541_0),.q1(n541_1));
  bfr _b_12410(.a(_w_14312),.q(_w_14313));
  spl2 g1662_s_0(.a(n1662),.q0(n1662_0),.q1(n1662_1));
  bfr _b_13649(.a(_w_15551),.q(_w_15552));
  bfr _b_9563(.a(_w_11465),.q(_w_11466));
  bfr _b_5082(.a(_w_6984),.q(_w_6985));
  bfr _b_5500(.a(_w_7402),.q(_w_7403));
  bfr _b_12369(.a(_w_14271),.q(_w_14272));
  spl2 g911_s_0(.a(n911),.q0(n911_0),.q1(_w_6169));
  bfr _b_4325(.a(_w_6227),.q(_w_6228));
  bfr _b_13609(.a(_w_15511),.q(_w_15512));
  spl2 g826_s_0(.a(n826),.q0(n826_0),.q1(n826_1));
  bfr _b_9030(.a(_w_10932),.q(_w_10933));
  spl2 g1777_s_0(.a(n1777),.q0(n1777_0),.q1(n1777_1));
  bfr _b_6813(.a(_w_8715),.q(_w_8716));
  spl2 g367_s_0(.a(n367),.q0(n367_0),.q1(n367_1));
  bfr _b_12969(.a(_w_14871),.q(_w_14872));
  bfr _b_5853(.a(_w_7755),.q(_w_7756));
  spl2 g533_s_0(.a(n533),.q0(n533_0),.q1(n533_1));
  bfr _b_9819(.a(_w_11721),.q(_w_11722));
  spl2 g1403_s_0(.a(n1403),.q0(n1403_0),.q1(n1403_1));
  bfr _b_4809(.a(_w_6711),.q(_w_6712));
  and_bi g363(.a(n348_1),.b(n351_1),.q(n363));
  bfr _b_9130(.a(_w_11032),.q(_w_11033));
  bfr _b_4192(.a(_w_6094),.q(_w_6095));
  or_bb g1434(.a(n1368_0),.b(n1433_0),.q(n1434));
  bfr _b_9513(.a(_w_11415),.q(_w_11416));
  spl2 g530_s_0(.a(n530),.q0(n530_0),.q1(n530_1));
  bfr _b_4919(.a(_w_6821),.q(_w_6822));
  bfr _b_3872(.a(_w_5774),.q(_w_5775));
  bfr _b_10867(.a(_w_12769),.q(_w_12770));
  bfr _b_4986(.a(_w_6888),.q(_w_6889));
  spl2 g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1));
  bfr _b_13674(.a(_w_15576),.q(_w_15577));
  bfr _b_8603(.a(_w_10505),.q(_w_10506));
  bfr _b_9102(.a(_w_11004),.q(_w_11005));
  spl2 g1681_s_0(.a(n1681),.q0(n1681_0),.q1(n1681_1));
  spl2 g1725_s_0(.a(n1725),.q0(n1725_0),.q1(n1725_1));
  spl2 g1613_s_0(.a(n1613),.q0(n1613_0),.q1(n1613_1));
  bfr _b_14003(.a(_w_15905),.q(_w_15906));
  spl2 g902_s_0(.a(n902),.q0(n902_0),.q1(n902_1));
  bfr _b_10685(.a(_w_12587),.q(_w_12588));
  bfr _b_8657(.a(_w_10559),.q(n209));
  spl2 g1075_s_0(.a(n1075),.q0(n1075_0),.q1(n1075_1));
  bfr _b_4788(.a(_w_6690),.q(_w_6691));
  bfr _b_13291(.a(_w_15193),.q(_w_15194));
  spl2 g1306_s_0(.a(n1306),.q0(n1306_0),.q1(n1306_1));
  bfr _b_3431(.a(_w_5333),.q(_w_5334));
  spl2 g635_s_0(.a(n635),.q0(n635_0),.q1(_w_6304));
  spl2 g174_s_0(.a(n174),.q0(n174_0),.q1(_w_6309));
  bfr _b_7778(.a(_w_9680),.q(_w_9681));
  spl2 g535_s_0(.a(n535),.q0(n535_0),.q1(n535_1));
  bfr _b_4994(.a(_w_6896),.q(_w_6897));
  spl2 g1031_s_0(.a(n1031),.q0(n1031_0),.q1(n1031_1));
  bfr _b_7761(.a(_w_9663),.q(_w_9664));
  spl2 g1039_s_0(.a(n1039),.q0(n1039_0),.q1(n1039_1));
  and_bi g128(.a(n102_1),.b(n126_1),.q(_w_11061));
  bfr _b_6099(.a(_w_8001),.q(_w_8002));
  spl2 g741_s_0(.a(n741),.q0(n741_0),.q1(n741_1));
  bfr _b_4368(.a(_w_6270),.q(_w_6271));
  spl2 g477_s_0(.a(n477),.q0(n477_0),.q1(n477_1));
  bfr _b_10383(.a(_w_12285),.q(_w_12286));
  or_bb g1776(.a(n1774_0),.b(n1775),.q(_w_14058));
  bfr _b_13367(.a(_w_15269),.q(_w_15270));
  bfr _b_12458(.a(_w_14360),.q(_w_14361));
  spl2 g1149_s_0(.a(n1149),.q0(n1149_0),.q1(_w_6317));
  bfr _b_8831(.a(_w_10733),.q(_w_10734));
  bfr _b_4804(.a(_w_6706),.q(_w_6707));
  spl3L g108_s_0(.a(n108),.q0(n108_0),.q1(_w_6321),.q2(_w_6323));
  bfr _b_11252(.a(_w_13154),.q(_w_13155));
  or_bb g1794(.a(n1784_0),.b(n1793_0),.q(n1794));
  spl2 g600_s_0(.a(n600),.q0(n600_0),.q1(_w_6325));
  bfr _b_10471(.a(_w_12373),.q(_w_12374));
  spl2 g201_s_0(.a(n201),.q0(n201_0),.q1(n201_1));
  spl2 g195_s_0(.a(n195),.q0(n195_0),.q1(n195_1));
  bfr _b_14159(.a(_w_16061),.q(_w_16062));
  bfr _b_8041(.a(_w_9943),.q(_w_9944));
  spl2 g373_s_0(.a(n373),.q0(n373_0),.q1(n373_1));
  bfr _b_6970(.a(_w_8872),.q(_w_8873));
  and_bb g57(.a(N273_7),.b(N52_5),.q(n57));
  or_bb g1154(.a(n1152_0),.b(n1153),.q(n1154));
  bfr _b_10141(.a(_w_12043),.q(_w_12044));
  bfr _b_13971(.a(_w_15873),.q(_w_15874));
  spl2 g36_s_0(.a(n36),.q0(_w_6329),.q1(n36_1));
  spl2 g1028_s_0(.a(n1028),.q0(n1028_0),.q1(_w_6330));
  bfr _b_4586(.a(_w_6488),.q(_w_6489));
  and_bi g1645(.a(n1614_1),.b(n1643_1),.q(_w_11227));
  bfr _b_8707(.a(_w_10609),.q(_w_10610));
  bfr _b_10701(.a(_w_12603),.q(_w_12604));
  bfr _b_6174(.a(_w_8076),.q(_w_8077));
  spl2 g1158_s_0(.a(n1158),.q0(n1158_0),.q1(n1158_1));
  spl2 g1412_s_0(.a(n1412),.q0(n1412_0),.q1(n1412_1));
  bfr _b_10120(.a(_w_12022),.q(_w_12023));
  spl2 g854_s_0(.a(n854),.q0(n854_0),.q1(n854_1));
  spl2 g723_s_0(.a(n723),.q0(n723_0),.q1(n723_1));
  bfr _b_13863(.a(_w_15765),.q(_w_15766));
  spl2 g524_s_0(.a(n524),.q0(n524_0),.q1(n524_1));
  bfr _b_8142(.a(_w_10044),.q(_w_10045));
  bfr _b_14368(.a(_w_16270),.q(_w_16271));
  spl2 g171_s_0(.a(n171),.q0(n171_0),.q1(n171_1));
  bfr _b_13403(.a(_w_15305),.q(_w_15306));
  spl4L N52_s_4(.a(N52_3),.q0(N52_16),.q1(N52_17),.q2(N52_18),.q3(N52_19));
  spl2 g625_s_0(.a(n625),.q0(n625_0),.q1(n625_1));
  spl2 g162_s_0(.a(n162),.q0(n162_0),.q1(_w_6334));
  spl2 g613_s_0(.a(n613),.q0(n613_0),.q1(n613_1));
  spl2 g1113_s_0(.a(n1113),.q0(n1113_0),.q1(_w_6338));
  bfr _b_12932(.a(_w_14834),.q(_w_14835));
  bfr _b_12529(.a(_w_14431),.q(_w_14432));
  bfr _b_11061(.a(_w_12963),.q(n1183));
  and_bi g1226(.a(n1224_0),.b(n1225),.q(n1226));
  and_bb g940(.a(N494_7),.b(N52_17),.q(_w_14281));
  and_bb g1029(.a(n1027_1),.b(n941_1),.q(_w_8360));
  spl2 g1376_s_0(.a(n1376),.q0(n1376_0),.q1(n1376_1));
  bfr _b_12495(.a(_w_14397),.q(_w_14398));
  bfr _b_12108(.a(_w_14010),.q(_w_14011));
  bfr _b_6772(.a(_w_8674),.q(_w_8675));
  and_bi g1782(.a(n1753_1),.b(n1756_1),.q(n1782));
  spl2 g214_s_0(.a(n214),.q0(n214_0),.q1(_w_6342));
  bfr _b_7987(.a(_w_9889),.q(_w_9890));
  bfr _b_4451(.a(_w_6353),.q(n658_1));
  bfr _b_8555(.a(_w_10457),.q(_w_10458));
  bfr _b_7752(.a(_w_9654),.q(n632));
  spl2 g1332_s_0(.a(n1332),.q0(n1332_0),.q1(n1332_1));
  bfr _b_3885(.a(_w_5787),.q(_w_5788));
  bfr _b_13175(.a(_w_15077),.q(_w_15078));
  bfr _b_12798(.a(_w_14700),.q(_w_14701));
  spl2 g727_s_0(.a(n727),.q0(n727_0),.q1(n727_1));
  spl2 g697_s_0(.a(n697),.q0(n697_0),.q1(n697_1));
  spl2 g415_s_0(.a(n415),.q0(n415_0),.q1(n415_1));
  bfr _b_7699(.a(_w_9601),.q(_w_9602));
  bfr _b_14357(.a(_w_16259),.q(_w_16260));
  bfr _b_12505(.a(_w_14407),.q(_w_14408));
  spl2 g1259_s_0(.a(n1259),.q0(n1259_0),.q1(n1259_1));
  spl2 g658_s_0(.a(n658),.q0(n658_0),.q1(_w_6350));
  bfr _b_14134(.a(_w_16036),.q(_w_16037));
  and_bi g1518(.a(n1517_0),.b(n1456_0),.q(n1518));
  bfr _b_3924(.a(_w_5826),.q(n1188_1));
  bfr _b_7315(.a(_w_9217),.q(n707));
  spl2 g663_s_0(.a(n663),.q0(n663_0),.q1(n663_1));
  bfr _b_4580(.a(_w_6482),.q(_w_6483));
  spl2 g1127_s_0(.a(n1127),.q0(n1127_0),.q1(n1127_1));
  spl4L N52_s_2(.a(N52_1),.q0(N52_8),.q1(N52_9),.q2(N52_10),.q3(_w_5347));
  or_bb g1410(.a(n1376_0),.b(n1409_0),.q(n1410));
  spl2 g1594_s_0(.a(n1594),.q0(n1594_0),.q1(_w_6354));
  bfr _b_5510(.a(_w_7412),.q(_w_7413));
  bfr _b_8288(.a(_w_10190),.q(_w_10191));
  spl2 g150_s_0(.a(n150),.q0(n150_0),.q1(_w_6358));
  spl2 g1610_s_0(.a(n1610),.q0(n1610_0),.q1(n1610_1));
  bfr _b_5721(.a(_w_7623),.q(_w_7624));
  bfr _b_13147(.a(_w_15049),.q(_w_15050));
  bfr _b_3439(.a(_w_5341),.q(_w_5342));
  bfr _b_10309(.a(_w_12211),.q(n272));
  spl2 g1221_s_0(.a(n1221),.q0(n1221_0),.q1(n1221_1));
  bfr _b_4828(.a(_w_6730),.q(_w_6731));
  spl4L N358_s_2(.a(N358_1),.q0(N358_8),.q1(N358_9),.q2(N358_10),.q3(N358_11));
  bfr _b_3501(.a(_w_5403),.q(_w_5404));
  spl2 g350_s_0(.a(n350),.q0(n350_0),.q1(n350_1));
  or_bb g1229(.a(n1227_0),.b(n1228),.q(n1229));
  and_bi g1307(.a(n1284_1),.b(n1305_1),.q(_w_13205));
  bfr _b_6664(.a(_w_8566),.q(_w_8567));
  bfr _b_5132(.a(_w_7034),.q(_w_7035));
  bfr _b_3531(.a(_w_5433),.q(_w_5434));
  bfr _b_5535(.a(_w_7437),.q(_w_7438));
  spl2 g198_s_0(.a(n198),.q0(n198_0),.q1(n198_1));
  bfr _b_3809(.a(_w_5711),.q(_w_5712));
  spl2 g1013_s_0(.a(n1013),.q0(n1013_0),.q1(n1013_1));
  bfr _b_3772(.a(_w_5674),.q(_w_5675));
  spl2 g454_s_0(.a(n454),.q0(n454_0),.q1(n454_1));
  spl2 g326_s_0(.a(n326),.q0(n326_0),.q1(n326_1));
  bfr _b_5770(.a(_w_7672),.q(_w_7673));
  bfr _b_8679(.a(_w_10581),.q(_w_10582));
  bfr _b_4682(.a(_w_6584),.q(_w_6585));
  spl2 g168_s_0(.a(n168),.q0(n168_0),.q1(_w_6362));
  and_bi g792(.a(n790_0),.b(n791),.q(n792));
  bfr _b_4093(.a(_w_5995),.q(_w_5996));
  spl2 g136_s_0(.a(n136),.q0(n136_0),.q1(n136_1));
  bfr _b_13998(.a(_w_15900),.q(_w_15901));
  spl2 g406_s_0(.a(n406),.q0(n406_0),.q1(_w_13492));
  bfr _b_8938(.a(_w_10840),.q(_w_10841));
  bfr _b_4836(.a(_w_6738),.q(_w_6739));
  bfr _b_10733(.a(_w_12635),.q(_w_12636));
  bfr _b_4593(.a(_w_6495),.q(_w_6496));
  and_bi g1187(.a(n1077_1),.b(n1080_1),.q(n1187));
  bfr _b_4346(.a(_w_6248),.q(_w_6249));
  spl2 g118_s_0(.a(n118),.q0(n118_0),.q1(_w_6366));
  or_bb g336(.a(n299_0),.b(n335_0),.q(n336));
  spl2 g1579_s_0(.a(n1579),.q0(n1579_0),.q1(n1579_1));
  bfr _b_14263(.a(_w_16165),.q(_w_16166));
  bfr _b_3646(.a(_w_5548),.q(_w_5549));
  bfr _b_12919(.a(_w_14821),.q(_w_14822));
  bfr _b_5740(.a(_w_7642),.q(_w_7643));
  spl2 g1782_s_0(.a(n1782),.q0(n1782_0),.q1(n1782_1));
  bfr _b_14284(.a(_w_16186),.q(_w_16187));
  bfr _b_8651(.a(_w_10553),.q(_w_10554));
  bfr _b_3921(.a(_w_5823),.q(_w_5824));
  spl2 g271_s_0(.a(n271),.q0(n271_0),.q1(n271_1));
  bfr _b_5042(.a(_w_6944),.q(_w_6945));
  bfr _b_7950(.a(_w_9852),.q(_w_9853));
  spl2 g685_s_0(.a(n685),.q0(n685_0),.q1(n685_1));
  spl2 g126_s_0(.a(n126),.q0(n126_0),.q1(n126_1));
  spl2 g1176_s_0(.a(n1176),.q0(n1176_0),.q1(n1176_1));
  bfr _b_4119(.a(_w_6021),.q(_w_6022));
  bfr _b_5301(.a(_w_7203),.q(_w_7204));
  spl2 g1070_s_0(.a(n1070),.q0(n1070_0),.q1(n1070_1));
  bfr _b_5547(.a(_w_7449),.q(_w_7450));
  bfr _b_11727(.a(_w_13629),.q(_w_13630));
  spl2 g784_s_0(.a(n784),.q0(n784_0),.q1(_w_6370));
  spl2 g107_s_0(.a(n107),.q0(n107_0),.q1(n107_1));
  bfr _b_13140(.a(_w_15042),.q(_w_15043));
  spl2 g757_s_0(.a(n757),.q0(n757_0),.q1(n757_1));
  spl2 g124_s_0(.a(n124),.q0(n124_0),.q1(_w_6374));
  spl2 g117_s_0(.a(n117),.q0(n117_0),.q1(n117_1));
  bfr _b_4004(.a(_w_5906),.q(_w_5907));
  spl2 g111_s_0(.a(n111),.q0(n111_0),.q1(n111_1));
  spl2 g1848_s_0(.a(n1848),.q0(n1848_0),.q1(n1848_1));
  bfr _b_13987(.a(_w_15889),.q(_w_15890));
  spl3L g42_s_0(.a(n42),.q0(n42_0),.q1(_w_6378),.q2(_w_6380));
  spl4L N205_s_4(.a(N205_3),.q0(N205_16),.q1(N205_17),.q2(N205_18),.q3(N205_19));
  spl2 g742_s_0(.a(n742),.q0(n742_0),.q1(_w_6165));
  bfr _b_3487(.a(_w_5389),.q(_w_5390));
  bfr _b_5446(.a(_w_7348),.q(_w_7349));
  bfr _b_10402(.a(_w_12304),.q(_w_12305));
  spl2 g390_s_0(.a(n390),.q0(n390_0),.q1(n390_1));
  bfr _b_10264(.a(_w_12166),.q(_w_12167));
  spl2 g447_s_0(.a(n447),.q0(n447_0),.q1(n447_1));
  bfr _b_6200(.a(_w_8102),.q(_w_8103));
  bfr _b_11946(.a(_w_13848),.q(_w_13849));
  bfr _b_9305(.a(_w_11207),.q(_w_11208));
  and_bi g303(.a(n256_1),.b(n259_1),.q(n303));
  bfr _b_3789(.a(_w_5691),.q(_w_5692));
  or_bb g1886(.a(n1884_0),.b(n1885),.q(_w_14771));
  spl2 g968_s_0(.a(n968),.q0(n968_0),.q1(_w_6382));
  bfr _b_14202(.a(_w_16104),.q(_w_16105));
  and_bi g1867(.a(n1866_0),.b(n1853_0),.q(n1867));
  and_bi g996(.a(n952_1),.b(n994_1),.q(_w_12513));
  spl2 g1080_s_0(.a(n1080),.q0(n1080_0),.q1(n1080_1));
  spl2 g242_s_0(.a(n242),.q0(n242_0),.q1(n242_1));
  spl2 g1137_s_0(.a(n1137),.q0(n1137_0),.q1(_w_6386));
  or_bb g863(.a(n843_0),.b(n862_0),.q(n863));
  spl4L N528_s_3(.a(N528_2),.q0(N528_12),.q1(N528_13),.q2(N528_14),.q3(N528_15));
  bfr _b_10470(.a(_w_12372),.q(_w_12373));
  bfr _b_8609(.a(_w_10511),.q(_w_10512));
  spl4L N256_s_4(.a(N256_3),.q0(_w_5569),.q1(N256_17),.q2(N256_18),.q3(N256_19));
  bfr _b_9308(.a(_w_11210),.q(_w_11211));
  bfr _b_13734(.a(_w_15636),.q(_w_15637));
  spl4L N528_s_0(.a(_w_16198),.q0(N528_0),.q1(N528_1),.q2(N528_2),.q3(N528_3));
  bfr _b_7777(.a(_w_9679),.q(_w_9680));
  bfr _b_7843(.a(_w_9745),.q(_w_9746));
  spl2 g827_s_0(.a(n827),.q0(n827_0),.q1(n827_1));
  bfr _b_9072(.a(_w_10974),.q(_w_10975));
  spl2 g222_s_0(.a(n222),.q0(n222_0),.q1(n222_1));
  bfr _b_3771(.a(_w_5673),.q(_w_5674));
  bfr _b_10629(.a(_w_12531),.q(_w_12532));
  spl2 g825_s_0(.a(n825),.q0(n825_0),.q1(n825_1));
  bfr _b_3875(.a(_w_5777),.q(_w_5778));
  bfr _b_7510(.a(_w_9412),.q(_w_9413));
  spl4L N137_s_4(.a(N137_3),.q0(N137_16),.q1(N137_17),.q2(N137_18),.q3(N137_19));
  bfr _b_14039(.a(_w_15941),.q(_w_15942));
  bfr _b_8393(.a(_w_10295),.q(_w_10296));
  spl4L N137_s_3(.a(N137_2),.q0(N137_12),.q1(_w_6394),.q2(_w_6402),.q3(_w_6414));
  spl4L N137_s_1(.a(N137_0),.q0(N137_4),.q1(N137_5),.q2(_w_6426),.q3(_w_6428));
  bfr _b_7106(.a(_w_9008),.q(_w_9009));
  bfr _b_3818(.a(_w_5720),.q(_w_5721));
  bfr _b_11096(.a(_w_12998),.q(_w_12999));
  bfr _b_5928(.a(_w_7830),.q(_w_7831));
  bfr _b_5077(.a(_w_6979),.q(_w_6980));
  spl2 g717_s_0(.a(n717),.q0(n717_0),.q1(n717_1));
  spl2 g289_s_0(.a(n289),.q0(n289_0),.q1(n289_1));
  and_bi g439(.a(n424_1),.b(n427_1),.q(n439));
  bfr _b_6405(.a(_w_8307),.q(_w_8308));
  bfr _b_13112(.a(_w_15014),.q(n226_1));
  spl2 g102_s_0(.a(n102),.q0(n102_0),.q1(n102_1));
  spl4L N154_s_0(.a(_w_15528),.q0(N154_0),.q1(_w_6466),.q2(_w_6490),.q3(_w_6546));
  bfr _b_12272(.a(_w_14174),.q(_w_14175));
  bfr _b_9948(.a(_w_11850),.q(_w_11851));
  spl2 g471_s_0(.a(n471),.q0(n471_0),.q1(n471_1));
  or_bb g869(.a(n841_0),.b(n868_0),.q(n869));
  and_bi g983(.a(n982_0),.b(n956_0),.q(n983));
  bfr _b_10478(.a(_w_12380),.q(_w_12381));
  and_bb g809(.a(n715_1),.b(n807_1),.q(_w_12078));
  spl4L N1_s_3(.a(N1_2),.q0(N1_12),.q1(_w_6634),.q2(_w_6642),.q3(_w_6654));
  bfr _b_12360(.a(_w_14262),.q(_w_14263));
  spl4L N1_s_2(.a(N1_1),.q0(N1_8),.q1(N1_9),.q2(N1_10),.q3(_w_6666));
  spl2 g156_s_0(.a(n156),.q0(n156_0),.q1(_w_6690));
  or_bb g1770(.a(n1768_0),.b(n1769),.q(_w_14308));
  spl2 g293_s_0(.a(n293),.q0(n293_0),.q1(n293_1));
  bfr _b_4226(.a(_w_6128),.q(_w_6129));
  bfr _b_12157(.a(_w_14059),.q(_w_14060));
  or_bb g1473(.a(n1471_0),.b(n1472_0),.q(n1473));
  bfr _b_5470(.a(_w_7372),.q(_w_7373));
  spl2 g240_s_0(.a(n240),.q0(n240_0),.q1(n240_1));
  spl2 g945_s_0(.a(n945),.q0(n945_0),.q1(n945_1));
  bfr _b_9998(.a(_w_11900),.q(_w_11901));
  bfr _b_10164(.a(_w_12066),.q(n1304));
  bfr _b_10249(.a(_w_12151),.q(_w_12152));
  spl2 g219_s_0(.a(n219),.q0(n219_0),.q1(n219_1));
  bfr _b_9033(.a(_w_10935),.q(_w_10936));
  spl2 g1803_s_0(.a(n1803),.q0(n1803_0),.q1(n1803_1));
  spl2 g631_s_0(.a(n631),.q0(n631_0),.q1(n631_1));
  spl2 g495_s_0(.a(n495),.q0(n495_0),.q1(n495_1));
  bfr _b_6722(.a(_w_8624),.q(_w_8625));
  spl2 g1037_s_0(.a(n1037),.q0(n1037_0),.q1(n1037_1));
  bfr _b_12704(.a(_w_14606),.q(_w_14607));
  bfr _b_9940(.a(_w_11842),.q(_w_11843));
  bfr _b_9437(.a(_w_11339),.q(_w_11340));
  bfr _b_14349(.a(_w_16251),.q(_w_16252));
  spl2 g1512_s_0(.a(n1512),.q0(n1512_0),.q1(n1512_1));
  spl2 g958_s_0(.a(n958),.q0(n958_0),.q1(n958_1));
  bfr _b_11689(.a(_w_13591),.q(_w_13592));
  bfr _b_4218(.a(_w_6120),.q(_w_6121));
  bfr _b_7946(.a(_w_9848),.q(_w_9849));
  bfr _b_11993(.a(_w_13895),.q(_w_13896));
  spl2 g1016_s_0(.a(n1016),.q0(n1016_0),.q1(_w_7571));
  and_bb g448(.a(N103_9),.b(N358_10),.q(_w_12434));
  spl2 g1033_s_0(.a(n1033),.q0(n1033_0),.q1(n1033_1));
  bfr _b_13188(.a(_w_15090),.q(_w_15091));
  bfr _b_9980(.a(_w_11882),.q(_w_11883));
  spl2 g1678_s_0(.a(n1678),.q0(n1678_0),.q1(n1678_1));
  bfr _b_5489(.a(_w_7391),.q(_w_7392));
  spl2 g498_s_0(.a(n498),.q0(n498_0),.q1(n498_1));
  bfr _b_4116(.a(_w_6018),.q(_w_6019));
  bfr _b_12013(.a(_w_13915),.q(_w_13916));
  bfr _b_11436(.a(_w_13338),.q(_w_13339));
  bfr _b_8432(.a(_w_10334),.q(_w_10335));
  bfr _b_10606(.a(_w_12508),.q(_w_12509));
  spl2 g1883_s_0(.a(n1883),.q0(n1883_0),.q1(n1883_1));
  spl2 g76_s_0(.a(n76),.q0(n76_0),.q1(n76_1));
  bfr _b_4410(.a(_w_6312),.q(n174_1));
  bfr _b_6605(.a(_w_8507),.q(_w_8508));
  bfr _b_7758(.a(_w_9660),.q(_w_9661));
  spl2 g54_s_0(.a(n54),.q0(n54_0),.q1(n54_1));
  spl4L N273_s_3(.a(N273_2),.q0(N273_12),.q1(N273_13),.q2(N273_14),.q3(N273_15));
  spl2 g48_s_0(.a(n48),.q0(n48_0),.q1(n48_1));
  spl4L N324_s_4(.a(N324_3),.q0(N324_16),.q1(N324_17),.q2(N324_18),.q3(N324_19));
  bfr _b_4859(.a(_w_6761),.q(_w_6762));
  bfr _b_13501(.a(_w_15403),.q(_w_15404));
  bfr _b_9388(.a(_w_11290),.q(_w_11291));
  spl4L N324_s_3(.a(N324_2),.q0(N324_12),.q1(N324_13),.q2(N324_14),.q3(N324_15));
  spl4L N426_s_3(.a(N426_2),.q0(N426_12),.q1(N426_13),.q2(N426_14),.q3(N426_15));
  bfr _b_5692(.a(_w_7594),.q(_w_7595));
  bfr _b_4591(.a(_w_6493),.q(_w_6494));
  bfr _b_4516(.a(_w_6418),.q(_w_6419));
  bfr _b_4167(.a(_w_6069),.q(_w_6070));
  bfr _b_4232(.a(_w_6134),.q(_w_6135));
  bfr _b_10204(.a(_w_12106),.q(_w_12107));
  bfr _b_3787(.a(_w_5689),.q(_w_5690));
  spl2 g928_s_0(.a(n928),.q0(n928_0),.q1(n928_1));
  bfr _b_4062(.a(_w_5964),.q(_w_5965));
  bfr _b_9343(.a(_w_11245),.q(_w_11246));
  spl2 g1694_s_0(.a(n1694),.q0(n1694_0),.q1(n1694_1));
  bfr _b_7986(.a(_w_9888),.q(_w_9889));
  spl2 g180_s_0(.a(n180),.q0(n180_0),.q1(n180_1));
  and_bi g332(.a(n330_0),.b(n331),.q(n332));
  bfr _b_10856(.a(_w_12758),.q(_w_12759));
  bfr _b_3557(.a(_w_5459),.q(_w_5460));
  spl4L N341_s_0(.a(_w_15545),.q0(N341_0),.q1(N341_1),.q2(N341_2),.q3(N341_3));
  spl2 g1235_s_0(.a(n1235),.q0(n1235_0),.q1(n1235_1));
  bfr _b_10344(.a(_w_12246),.q(_w_12247));
  and_bb g1687(.a(n1684_1),.b(n1685_1),.q(_w_12097));
  spl2 g145_s_0(.a(n145),.q0(n145_0),.q1(n145_1));
  bfr _b_8606(.a(_w_10508),.q(_w_10509));
  bfr _b_4178(.a(_w_6080),.q(N239_3));
  bfr _b_8175(.a(_w_10077),.q(_w_10078));
  spl4L N358_s_0(.a(_w_15571),.q0(N358_0),.q1(N358_1),.q2(N358_2),.q3(N358_3));
  bfr _b_4318(.a(_w_6220),.q(_w_6221));
  bfr _b_6116(.a(_w_8018),.q(_w_8019));
  spl4L N409_s_1(.a(N409_0),.q0(N409_4),.q1(N409_5),.q2(N409_6),.q3(N409_7));
  bfr _b_4370(.a(_w_6272),.q(_w_6273));
  spl4L N409_s_0(.a(_w_15670),.q0(N409_0),.q1(N409_1),.q2(N409_2),.q3(N409_3));
  bfr _b_8899(.a(_w_10801),.q(n1096));
  bfr _b_4699(.a(_w_6601),.q(_w_6602));
  bfr _b_9719(.a(_w_11621),.q(_w_11622));
  spl2 g77_s_0(.a(n77),.q0(n77_0),.q1(n77_1));
  spl2 g1650_s_0(.a(n1650),.q0(n1650_0),.q1(n1650_1));
  spl3L g192_s_0(.a(n192),.q0(n192_0),.q1(_w_6694),.q2(_w_6696));
  bfr _b_13092(.a(_w_14994),.q(_w_14995));
  bfr _b_4187(.a(_w_6089),.q(_w_6090));
  and_bi g990(.a(n954_1),.b(n988_1),.q(_w_8368));
  bfr _b_6022(.a(_w_7924),.q(_w_7925));
  spl4L N426_s_4(.a(N426_3),.q0(N426_16),.q1(N426_17),.q2(N426_18),.q3(_w_6702));
  and_bi g710(.a(n612_1),.b(n708_1),.q(_w_9210));
  bfr _b_8503(.a(_w_10405),.q(_w_10406));
  bfr _b_13488(.a(_w_15390),.q(_w_15391));
  spl2 g789_s_0(.a(n789),.q0(n789_0),.q1(n789_1));
  and_bi g1857(.a(n1827_1),.b(n1830_1),.q(n1857));
  spl4L N460_s_4(.a(N460_3),.q0(N460_16),.q1(N460_17),.q2(N460_18),.q3(N460_19));
  bfr _b_7128(.a(_w_9030),.q(_w_9031));
  bfr _b_11768(.a(_w_13670),.q(_w_13671));
  spl4L N460_s_3(.a(N460_2),.q0(N460_12),.q1(N460_13),.q2(N460_14),.q3(N460_15));
  bfr _b_4951(.a(_w_6853),.q(_w_6854));
  bfr _b_11972(.a(_w_13874),.q(_w_13875));
  bfr _b_8294(.a(_w_10196),.q(_w_10197));
  spl2 g1226_s_0(.a(n1226),.q0(n1226_0),.q1(n1226_1));
  spl4L N477_s_3(.a(N477_2),.q0(N477_12),.q1(N477_13),.q2(N477_14),.q3(N477_15));
  bfr _b_13172(.a(_w_15074),.q(_w_15075));
  bfr _b_5208(.a(_w_7110),.q(_w_7111));
  bfr _b_4203(.a(_w_6105),.q(_w_6106));
  spl2 g216_s_0(.a(n216),.q0(n216_0),.q1(n216_1));
  spl2 g1279_s_0(.a(n1279),.q0(n1279_0),.q1(n1279_1));
  bfr _b_6790(.a(_w_8692),.q(_w_8693));
  spl4L N477_s_2(.a(N477_1),.q0(N477_8),.q1(N477_9),.q2(N477_10),.q3(N477_11));
  bfr _b_4418(.a(_w_6320),.q(n1149_1));
  bfr _b_11203(.a(_w_13105),.q(_w_13106));
  bfr _b_6580(.a(_w_8482),.q(_w_8483));
  spl2 g971_s_0(.a(n971),.q0(n971_0),.q1(n971_1));
  spl2 g277_s_0(.a(n277),.q0(n277_0),.q1(n277_1));
  bfr _b_14151(.a(_w_16053),.q(_w_16054));
  bfr _b_11270(.a(_w_13172),.q(_w_13173));
  or_bb g330(.a(n301_0),.b(n329_0),.q(n330));
  spl4L N477_s_1(.a(N477_0),.q0(N477_4),.q1(N477_5),.q2(N477_6),.q3(N477_7));
  bfr _b_4322(.a(_w_6224),.q(_w_6225));
  spl4L N511_s_4(.a(N511_3),.q0(N511_16),.q1(N511_17),.q2(N511_18),.q3(N511_19));
  bfr _b_4980(.a(_w_6882),.q(_w_6883));
  bfr _b_6178(.a(_w_8080),.q(_w_8081));
  spl4L N511_s_2(.a(N511_1),.q0(N511_8),.q1(N511_9),.q2(N511_10),.q3(N511_11));
  bfr _b_7528(.a(_w_9430),.q(_w_9431));
  bfr _b_14205(.a(_w_16107),.q(_w_16019));
  spl4L N511_s_0(.a(_w_16108),.q0(N511_0),.q1(N511_1),.q2(N511_2),.q3(N511_3));
  bfr _b_6696(.a(_w_8598),.q(_w_8599));
  bfr _b_8252(.a(_w_10154),.q(_w_10155));
  bfr _b_3461(.a(_w_5363),.q(_w_5364));
  bfr _b_12137(.a(_w_14039),.q(_w_14040));
  spl2 g1887_s_0(.a(n1887),.q0(n1887_0),.q1(_w_14943));
  bfr _b_5704(.a(_w_7606),.q(_w_7607));
  spl2 g1162_s_0(.a(n1162),.q0(n1162_0),.q1(n1162_1));
  spl4L N137_s_0(.a(_w_15527),.q0(N137_0),.q1(_w_6710),.q2(_w_6734),.q3(_w_6790));
  spl2 g1433_s_0(.a(n1433),.q0(n1433_0),.q1(n1433_1));
  spl2 g115_s_0(.a(n115),.q0(n115_0),.q1(n115_1));
  spl2 g480_s_0(.a(n480),.q0(n480_0),.q1(n480_1));
  bfr _b_9811(.a(_w_11713),.q(_w_11714));
  bfr _b_4844(.a(_w_6746),.q(_w_6747));
  spl2 g1815_s_0(.a(n1815),.q0(n1815_0),.q1(n1815_1));
  spl2 g1653_s_0(.a(n1653),.q0(n1653_0),.q1(_w_6878));
  spl4L N103_s_4(.a(N103_3),.q0(N103_16),.q1(N103_17),.q2(N103_18),.q3(N103_19));
  spl2 g205_s_0(.a(n205),.q0(n205_0),.q1(n205_1));
  bfr _b_13659(.a(_w_15561),.q(_w_15562));
  bfr _b_8901(.a(_w_10803),.q(_w_10804));
  bfr _b_3408(.a(_w_5310),.q(n857_1));
  spl2 g1430_s_0(.a(n1430),.q0(n1430_0),.q1(n1430_1));
  bfr _b_10414(.a(_w_12316),.q(_w_12317));
  spl2 g720_s_0(.a(n720),.q0(n720_0),.q1(n720_1));
  bfr _b_3601(.a(_w_5503),.q(_w_5504));
  bfr _b_8595(.a(_w_10497),.q(_w_10498));
  bfr _b_8221(.a(_w_10123),.q(_w_10124));
  bfr _b_8880(.a(_w_10782),.q(N52_6));
  spl2 g208_s_0(.a(n208),.q0(n208_0),.q1(_w_7054));
  spl2 g1030_s_0(.a(n1030),.q0(n1030_0),.q1(n1030_1));
  spl2 g259_s_0(.a(n259),.q0(n259_0),.q1(n259_1));
  bfr _b_10865(.a(_w_12767),.q(_w_12768));
  bfr _b_5479(.a(_w_7381),.q(_w_7382));
  bfr _b_3790(.a(_w_5692),.q(_w_5693));
  bfr _b_3495(.a(_w_5397),.q(_w_5398));
  spl2 g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1));
  spl2 g1223_s_0(.a(n1223),.q0(n1223_0),.q1(n1223_1));
  spl2 g948_s_0(.a(n948),.q0(n948_0),.q1(n948_1));
  or_bb g670(.a(n625_0),.b(n669_0),.q(n670));
  bfr _b_11676(.a(_w_13578),.q(n577));
  bfr _b_3610(.a(_w_5512),.q(_w_5513));
  bfr _b_10149(.a(_w_12051),.q(_w_12052));
  bfr _b_7360(.a(_w_9262),.q(_w_9263));
  bfr _b_4348(.a(_w_6250),.q(_w_6251));
  bfr _b_5858(.a(_w_7760),.q(_w_7761));
  spl2 g1697_s_0(.a(n1697),.q0(n1697_0),.q1(n1697_1));
  spl2 g236_s_0(.a(n236),.q0(n236_0),.q1(n236_1));
  spl2 g34_s_0(.a(N545_0),.q0(_w_7062),.q1(N545_1));
  bfr _b_4652(.a(_w_6554),.q(_w_6555));
  or_bb g1327(.a(n1277_0),.b(n1326_0),.q(n1327));
  spl4L N35_s_4(.a(N35_3),.q0(N35_16),.q1(N35_17),.q2(N35_18),.q3(N35_19));
  spl4L N35_s_2(.a(N35_1),.q0(N35_8),.q1(N35_9),.q2(N35_10),.q3(_w_7235));
  bfr _b_4662(.a(_w_6564),.q(_w_6565));
  bfr _b_6625(.a(_w_8527),.q(_w_8528));
  bfr _b_8256(.a(_w_10158),.q(_w_10159));
  bfr _b_8926(.a(_w_10828),.q(_w_10829));
  spl2 g569_s_0(.a(n569),.q0(n569_0),.q1(n569_1));
  spl2 g1759_s_0(.a(n1759),.q0(n1759_0),.q1(_w_7263));
  bfr _b_10523(.a(_w_12425),.q(n482));
  spl2 g315_s_0(.a(n315),.q0(n315_0),.q1(n315_1));
  bfr _b_8983(.a(_w_10885),.q(_w_10886));
  spl2 g417_s_0(.a(n417),.q0(n417_0),.q1(n417_1));
  bfr _b_7139(.a(_w_9041),.q(_w_9042));
  bfr _b_9226(.a(_w_11128),.q(_w_11129));
  bfr _b_6751(.a(_w_8653),.q(_w_8654));
  spl2 g1064_s_0(.a(n1064),.q0(n1064_0),.q1(n1064_1));
  bfr _b_7664(.a(_w_9566),.q(n604));
  spl2 g1379_s_0(.a(n1379),.q0(n1379_0),.q1(n1379_1));
  spl4L N307_s_2(.a(N307_1),.q0(N307_8),.q1(N307_9),.q2(N307_10),.q3(N307_11));
  bfr _b_4902(.a(_w_6804),.q(_w_6805));
  bfr _b_4151(.a(_w_6053),.q(_w_6054));
  spl2 g465_s_0(.a(n465),.q0(n465_0),.q1(n465_1));
  spl2 g1049_s_0(.a(n1049),.q0(n1049_0),.q1(n1049_1));
  spl2 g335_s_0(.a(n335),.q0(n335_0),.q1(n335_1));
  spl2 g649_s_0(.a(n649),.q0(n649_0),.q1(n649_1));
  or_bb g1892(.a(n1890_0),.b(n1891),.q(_w_14825));
  spl2 g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1));
  bfr _b_3897(.a(_w_5799),.q(_w_5800));
  bfr _b_13400(.a(_w_15302),.q(_w_15303));
  bfr _b_6375(.a(_w_8277),.q(_w_8278));
  bfr _b_5072(.a(_w_6974),.q(_w_6975));
  bfr _b_12801(.a(_w_14703),.q(_w_14704));
  spl2 g353_s_0(.a(n353),.q0(n353_0),.q1(n353_1));
  bfr _b_11905(.a(_w_13807),.q(_w_13808));
  spl2 g1746_s_0(.a(n1746),.q0(n1746_0),.q1(n1746_1));
  spl2 g1338_s_0(.a(n1338),.q0(n1338_0),.q1(n1338_1));
  bfr _b_9918(.a(_w_11820),.q(_w_11821));
  spl2 g427_s_0(.a(n427),.q0(n427_0),.q1(n427_1));
  bfr _b_9688(.a(_w_11590),.q(_w_11591));
  spl2 g333_s_0(.a(n333),.q0(n333_0),.q1(n333_1));
  spl2 g1272_s_0(.a(n1272),.q0(n1272_0),.q1(n1272_1));
  spl2 g1040_s_0(.a(n1040),.q0(n1040_0),.q1(_w_5561));
  and_bb g924(.a(n823_1),.b(n922_1),.q(_w_11068));
  bfr _b_7228(.a(_w_9130),.q(n1504));
  and_bi g1469(.a(n1392_1),.b(n1395_1),.q(n1469));
  bfr _b_9022(.a(_w_10924),.q(_w_10925));
  bfr _b_10381(.a(_w_12283),.q(_w_12284));
  bfr _b_5694(.a(_w_7596),.q(_w_7597));
  spl2 g961_s_0(.a(n961),.q0(n961_0),.q1(n961_1));
  spl2 g91_s_0(.a(n91),.q0(n91_0),.q1(n91_1));
  spl2 g839_s_0(.a(n839),.q0(n839_0),.q1(n839_1));
  bfr _b_5679(.a(_w_7581),.q(_w_7582));
  bfr _b_9076(.a(_w_10978),.q(_w_10979));
  spl2 g1800_s_0(.a(n1800),.q0(n1800_0),.q1(_w_7471));
  bfr _b_7759(.a(_w_9661),.q(_w_9662));
  bfr _b_12327(.a(_w_14229),.q(n1410_1));
  bfr _b_11834(.a(_w_13736),.q(_w_13737));
  bfr _b_5941(.a(_w_7843),.q(_w_7844));
  spl2 g527_s_0(.a(n527),.q0(n527_0),.q1(n527_1));
  spl2 g1042_s_0(.a(n1042),.q0(n1042_0),.q1(n1042_1));
  spl2 g270_s_0(.a(n270),.q0(n270_0),.q1(n270_1));
  bfr _b_9803(.a(_w_11705),.q(_w_11706));
  spl2 g41_s_0(.a(n41),.q0(n41_0),.q1(n41_1));
  bfr _b_12949(.a(_w_14851),.q(_w_14852));
  spl2 g1619_s_0(.a(n1619),.q0(n1619_0),.q1(n1619_1));
  spl2 g82_s_0(.a(n82),.q0(n82_0),.q1(_w_7475));
  bfr _b_9109(.a(_w_11011),.q(_w_11012));
  bfr _b_5051(.a(_w_6953),.q(_w_6954));
  bfr _b_7578(.a(_w_9480),.q(_w_9481));
  spl4L N69_s_2(.a(N69_1),.q0(N69_8),.q1(N69_9),.q2(N69_10),.q3(_w_7511));
  bfr _b_14304(.a(_w_16206),.q(_w_16207));
  bfr _b_7369(.a(_w_9271),.q(_w_9272));
  spl2 g489_s_0(.a(n489),.q0(n489_0),.q1(n489_1));
  and_bi g195(.a(n194),.b(n192_0),.q(n195));
  bfr _b_11859(.a(_w_13761),.q(_w_13762));
  bfr _b_3950(.a(_w_5852),.q(n905_1));
  bfr _b_8596(.a(_w_10498),.q(_w_10499));
  spl2 g312_s_0(.a(n312),.q0(n312_0),.q1(_w_7539));
  bfr _b_7083(.a(_w_8985),.q(_w_8986));
  spl2 g52_s_0(.a(n52),.q0(n52_0),.q1(n52_1));
  bfr _b_3782(.a(_w_5684),.q(_w_5685));
  bfr _b_11086(.a(_w_12988),.q(_w_12989));
  and_bi g574(.a(n532_1),.b(n572_1),.q(_w_11022));
  spl2 g264_s_0(.a(n264),.q0(n264_0),.q1(n264_1));
  bfr _b_11960(.a(_w_13862),.q(n1498));
  bfr _b_4903(.a(_w_6805),.q(_w_6806));
  spl2 g234_s_0(.a(n234),.q0(n234_0),.q1(n234_1));
  spl2 g526_s_0(.a(n526),.q0(n526_0),.q1(n526_1));
  bfr _b_12520(.a(_w_14422),.q(_w_14423));
  bfr _b_10755(.a(_w_12657),.q(_w_12658));
  bfr _b_4539(.a(_w_6441),.q(_w_6442));
  bfr _b_6420(.a(_w_8322),.q(_w_8323));
  or_bb g514(.a(n437_0),.b(n513_0),.q(n514));
  bfr _b_4510(.a(_w_6412),.q(_w_6413));
  spl2 g1452_s_0(.a(n1452),.q0(n1452_0),.q1(n1452_1));
  bfr _b_5586(.a(_w_7488),.q(_w_7489));
  bfr _b_8557(.a(_w_10459),.q(_w_10460));
  bfr _b_4698(.a(_w_6600),.q(_w_6601));
  bfr _b_12102(.a(_w_14004),.q(_w_14005));
  bfr _b_8653(.a(_w_10555),.q(_w_10556));
  spl2 g65_s_0(.a(n65),.q0(n65_0),.q1(n65_1));
  and_bi g1271(.a(n1242_1),.b(n1245_1),.q(n1271));
  bfr _b_11196(.a(_w_13098),.q(_w_13099));
  bfr _b_9164(.a(_w_11066),.q(n887_1));
  spl4L N494_s_4(.a(N494_3),.q0(N494_16),.q1(N494_17),.q2(N494_18),.q3(N494_19));
  spl4L N494_s_2(.a(N494_1),.q0(N494_8),.q1(N494_9),.q2(N494_10),.q3(N494_11));
  bfr _b_7014(.a(_w_8916),.q(_w_8917));
  spl4L N494_s_1(.a(N494_0),.q0(N494_4),.q1(N494_5),.q2(N494_6),.q3(N494_7));
  bfr _b_3465(.a(_w_5367),.q(_w_5368));
  bfr _b_13808(.a(_w_15710),.q(_w_15711));
  spl4L N494_s_0(.a(_w_16019),.q0(N494_0),.q1(N494_1),.q2(N494_2),.q3(N494_3));
  spl2 g520_s_0(.a(n520),.q0(n520_0),.q1(n520_1));
  bfr _b_9793(.a(_w_11695),.q(_w_11696));
  spl2 g1185_s_0(.a(n1185),.q0(n1185_0),.q1(n1185_1));
  spl2 g1244_s_0(.a(n1244),.q0(n1244_0),.q1(n1244_1));
  bfr _b_5028(.a(_w_6930),.q(_w_6931));
  bfr _b_13212(.a(_w_15114),.q(n313));
  bfr _b_10404(.a(_w_12306),.q(_w_12307));
  bfr _b_3806(.a(_w_5708),.q(_w_5709));
  spl2 g1073_s_0(.a(n1073),.q0(n1073_0),.q1(n1073_1));
  bfr _b_8298(.a(_w_10200),.q(n888));
  spl4L N222_s_4(.a(N222_3),.q0(_w_7577),.q1(_w_7602),.q2(_w_7605),.q3(N222_19));
  bfr _b_4475(.a(_w_6377),.q(n124_1));
  spl4L N222_s_2(.a(N222_1),.q0(_w_7608),.q1(_w_7632),.q2(_w_7636),.q3(N222_11));
  bfr _b_7337(.a(_w_9239),.q(_w_9240));
  bfr _b_13087(.a(_w_14989),.q(_w_14990));
  bfr _b_11939(.a(_w_13841),.q(_w_13842));
  bfr _b_8769(.a(_w_10671),.q(_w_10672));
  bfr _b_12160(.a(_w_14062),.q(_w_14063));
  spl4L N222_s_1(.a(N222_0),.q0(N222_4),.q1(_w_7640),.q2(_w_7680),.q3(_w_7720));
  spl4L N273_s_2(.a(N273_1),.q0(N273_8),.q1(N273_9),.q2(N273_10),.q3(N273_11));
  bfr _b_8961(.a(_w_10863),.q(n1125_1));
  spl4L N273_s_1(.a(N273_0),.q0(_w_7875),.q1(N273_5),.q2(N273_6),.q3(N273_7));
  bfr _b_3644(.a(_w_5546),.q(n1558_1));
  bfr _b_8071(.a(_w_9973),.q(n595));
  spl2 g1485_s_0(.a(n1485),.q0(n1485_0),.q1(_w_7877));
  or_bb g594(.a(n525_0),.b(n593_0),.q(n594));
  bfr _b_5934(.a(_w_7836),.q(_w_7837));
  spl2 g1756_s_0(.a(n1756),.q0(n1756_0),.q1(n1756_1));
  bfr _b_6453(.a(_w_8355),.q(n1045));
  spl2 g1063_s_0(.a(n1063),.q0(n1063_0),.q1(n1063_1));
  bfr _b_11219(.a(_w_13121),.q(_w_13122));
  bfr _b_4469(.a(_w_6371),.q(_w_6372));
  spl2 g106_s_0(.a(n106),.q0(n106_0),.q1(n106_1));
  bfr _b_10620(.a(_w_12522),.q(n1833_1));
  bfr _b_4579(.a(_w_6481),.q(_w_6482));
  bfr _b_4460(.a(_w_6362),.q(_w_6363));
  spl4L N290_s_0(.a(_w_15538),.q0(N290_0),.q1(N290_1),.q2(N290_2),.q3(N290_3));
  spl2 g1600_s_0(.a(n1600),.q0(n1600_0),.q1(_w_9655));
  bfr _b_3550(.a(_w_5452),.q(_w_5453));
  spl2 g1802_s_0(.a(n1802),.q0(n1802_0),.q1(n1802_1));
  spl2 g1089_s_0(.a(n1089),.q0(n1089_0),.q1(_w_10561));
  spl2 g1366_s_0(.a(n1366),.q0(n1366_0),.q1(n1366_1));
  spl2 g843_s_0(.a(n843),.q0(n843_0),.q1(n843_1));
  bfr _b_7503(.a(_w_9405),.q(_w_9406));
  bfr _b_13284(.a(_w_15186),.q(_w_15187));
  bfr _b_12393(.a(_w_14295),.q(_w_14296));
  bfr _b_12348(.a(_w_14250),.q(_w_14251));
  spl2 g238_s_0(.a(n238),.q0(n238_0),.q1(n238_1));
  bfr _b_4970(.a(_w_6872),.q(_w_6873));
  spl2 g245_s_0(.a(n245),.q0(n245_0),.q1(n245_1));
  bfr _b_5056(.a(_w_6958),.q(_w_6959));
  spl2 g1062_s_0(.a(n1062),.q0(n1062_0),.q1(n1062_1));
  spl3L g378_s_0(.a(n378),.q0(n378_0),.q1(_w_7892),.q2(_w_7894));
  spl2 g714_s_0(.a(n714),.q0(n714_0),.q1(n714_1));
  spl4L N460_s_0(.a(_w_15861),.q0(N460_0),.q1(N460_1),.q2(N460_2),.q3(N460_3));
  bfr _b_7156(.a(_w_9058),.q(_w_9059));
  spl4L N188_s_3(.a(N188_2),.q0(N188_12),.q1(_w_7896),.q2(_w_7904),.q3(_w_7916));
  bfr _b_5279(.a(_w_7181),.q(_w_7182));
  bfr _b_4118(.a(_w_6020),.q(_w_6021));
  spl2 g1566_s_0(.a(n1566),.q0(n1566_0),.q1(n1566_1));
  bfr _b_9028(.a(_w_10930),.q(_w_10931));
  bfr _b_3744(.a(_w_5646),.q(_w_5647));
  bfr _b_4436(.a(_w_6338),.q(_w_6339));
  spl3L g35_s_0(.a(n35),.q0(n35_0),.q1(n35_1),.q2(n35_2));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(_w_7956));
  bfr _b_11603(.a(_w_13505),.q(_w_13506));
  bfr _b_8545(.a(_w_10447),.q(_w_10448));
  spl2 g834_s_0(.a(n834),.q0(n834_0),.q1(n834_1));
  spl3L g246_s_0(.a(n246),.q0(n246_0),.q1(_w_7960),.q2(_w_7962));
  spl2 g403_s_0(.a(n403),.q0(n403_0),.q1(n403_1));
  or_bb g1206(.a(n1180_0),.b(n1205_0),.q(n1206));
  bfr _b_5520(.a(_w_7422),.q(_w_7423));
  bfr _b_4441(.a(_w_6343),.q(_w_6344));
  bfr _b_9344(.a(_w_11246),.q(_w_11247));
  bfr _b_8368(.a(_w_10270),.q(_w_10271));
  spl2 g563_s_0(.a(n563),.q0(n563_0),.q1(n563_1));
  bfr _b_11181(.a(_w_13083),.q(_w_13084));
  bfr _b_7314(.a(_w_9216),.q(n106));
  bfr _b_5631(.a(_w_7533),.q(_w_7534));
  spl2 g1056_s_0(.a(n1056),.q0(n1056_0),.q1(n1056_1));
  bfr _b_9622(.a(_w_11524),.q(_w_11525));
  spl2 g1022_s_0(.a(n1022),.q0(n1022_0),.q1(_w_8028));
  bfr _b_11180(.a(_w_13082),.q(_w_13083));
  spl2 g1019_s_0(.a(n1019),.q0(n1019_0),.q1(n1019_1));
  bfr _b_3908(.a(_w_5810),.q(_w_5811));
  and_bi g344(.a(n342_0),.b(n343),.q(n344));
  bfr _b_11700(.a(_w_13602),.q(_w_13603));
  bfr _b_4240(.a(_w_6142),.q(_w_6143));
  and_bb g374(.a(N120_7),.b(N324_11),.q(_w_8565));
  spl2 g729_s_0(.a(n729),.q0(n729_0),.q1(n729_1));
  bfr _b_5816(.a(_w_7718),.q(_w_7719));
  bfr _b_11743(.a(_w_13645),.q(_w_13646));
  bfr _b_10906(.a(_w_12808),.q(_w_12809));
  bfr _b_10540(.a(_w_12442),.q(_w_12443));
  and_bi g1127(.a(n1125_0),.b(n1126),.q(n1127));
  bfr _b_8129(.a(_w_10031),.q(_w_10032));
  spl2 g609_s_0(.a(n609),.q0(n609_0),.q1(n609_1));
  bfr _b_6057(.a(_w_7959),.q(n250_1));
  spl2 g279_s_0(.a(n279),.q0(n279_0),.q1(n279_1));
  bfr _b_11392(.a(_w_13294),.q(_w_13295));
  bfr _b_9970(.a(_w_11872),.q(_w_11873));
  spl2 g282_s_0(.a(n282),.q0(n282_0),.q1(n282_1));
  spl2 g446_s_0(.a(n446),.q0(n446_0),.q1(n446_1));
  or_bb g117(.a(n115_0),.b(n116),.q(n117));
  bfr _b_13498(.a(_w_15400),.q(_w_15401));
  bfr _b_11811(.a(_w_13713),.q(_w_13714));
  bfr _b_5954(.a(_w_7856),.q(_w_7857));
  bfr _b_6010(.a(_w_7912),.q(_w_7913));
  bfr _b_13595(.a(_w_15497),.q(_w_15498));
  bfr _b_9611(.a(_w_11513),.q(_w_11514));
  bfr _b_6956(.a(_w_8858),.q(_w_8859));
  spl2 g283_s_0(.a(n283),.q0(n283_0),.q1(n283_1));
  bfr _b_3627(.a(_w_5529),.q(_w_5530));
  or_bb g1439(.a(n1437_0),.b(n1438),.q(n1439));
  bfr _b_4884(.a(_w_6786),.q(_w_6787));
  bfr _b_14279(.a(_w_16181),.q(_w_16182));
  bfr _b_12506(.a(_w_14408),.q(_w_14409));
  bfr _b_3991(.a(_w_5893),.q(_w_5894));
  bfr _b_13545(.a(_w_15447),.q(_w_15448));
  bfr _b_9854(.a(_w_11756),.q(_w_11757));
  spl2 g1869_s_0(.a(n1869),.q0(n1869_0),.q1(n1869_1));
  spl2 g244_s_0(.a(n244),.q0(n244_0),.q1(n244_1));
  spl2 g285_s_0(.a(n285),.q0(n285_0),.q1(n285_1));
  bfr _b_5563(.a(_w_7465),.q(_w_7466));
  bfr _b_7206(.a(_w_9108),.q(_w_9109));
  bfr _b_3960(.a(_w_5862),.q(_w_5863));
  bfr _b_7683(.a(_w_9585),.q(_w_9586));
  spl2 g371_s_0(.a(n371),.q0(n371_0),.q1(n371_1));
  spl2 g1832_s_0(.a(n1832),.q0(n1832_0),.q1(n1832_1));
  and_bi g578(.a(n576_0),.b(n577),.q(n578));
  spl2 g233_s_0(.a(n233),.q0(n233_0),.q1(n233_1));
  spl2 g338_s_0(.a(n338),.q0(n338_0),.q1(n338_1));
  bfr _b_7505(.a(_w_9407),.q(_w_9408));
  spl2 g196_s_0(.a(n196),.q0(n196_0),.q1(_w_8032));
  spl2 g614_s_0(.a(n614),.q0(n614_0),.q1(n614_1));
  spl2 g414_s_0(.a(n414),.q0(n414_0),.q1(n414_1));
  bfr _b_8930(.a(_w_10832),.q(_w_10833));
  bfr _b_9438(.a(_w_11340),.q(_w_11341));
  bfr _b_12585(.a(_w_14487),.q(_w_14488));
  bfr _b_11537(.a(_w_13439),.q(_w_13440));
  bfr _b_4056(.a(_w_5958),.q(_w_5959));
  bfr _b_3780(.a(_w_5682),.q(_w_5683));
  spl2 g950_s_0(.a(n950),.q0(n950_0),.q1(n950_1));
  and_bb g1679(.a(N205_16),.b(N477_16),.q(n1679));
  bfr _b_9915(.a(_w_11817),.q(_w_11818));
  bfr _b_8394(.a(_w_10296),.q(_w_10297));
  bfr _b_12482(.a(_w_14384),.q(_w_14385));
  spl2 g341_s_0(.a(n341),.q0(n341_0),.q1(n341_1));
  spl2 g627_s_0(.a(n627),.q0(n627_0),.q1(n627_1));
  spl2 g317_s_0(.a(n317),.q0(n317_0),.q1(n317_1));
  bfr _b_7282(.a(_w_9184),.q(n730));
  bfr _b_12551(.a(_w_14453),.q(_w_14454));
  bfr _b_8451(.a(_w_10353),.q(_w_10354));
  bfr _b_9373(.a(_w_11275),.q(_w_11276));
  bfr _b_12220(.a(_w_14122),.q(n1720));
  spl2 g1281_s_0(.a(n1281),.q0(n1281_0),.q1(n1281_1));
  spl2 g1350_s_0(.a(n1350),.q0(n1350_0),.q1(n1350_1));
  bfr _b_6012(.a(_w_7914),.q(_w_7915));
  spl2 g801_s_0(.a(n801),.q0(n801_0),.q1(n801_1));
  bfr _b_5084(.a(_w_6986),.q(_w_6987));
  bfr _b_9298(.a(_w_11200),.q(_w_11201));
  bfr _b_11342(.a(_w_13244),.q(_w_13245));
  bfr _b_3816(.a(_w_5718),.q(_w_5719));
  spl4L N392_s_0(.a(_w_15621),.q0(N392_0),.q1(N392_1),.q2(N392_2),.q3(N392_3));
  spl2 g1344_s_0(.a(n1344),.q0(n1344_0),.q1(n1344_1));
  bfr _b_13946(.a(_w_15848),.q(_w_15849));
  bfr _b_7445(.a(_w_9347),.q(_w_9348));
  spl2 g239_s_0(.a(n239),.q0(n239_0),.q1(n239_1));
  bfr _b_11952(.a(_w_13854),.q(n224));
  bfr _b_9273(.a(_w_11175),.q(_w_11176));
  bfr _b_6333(.a(_w_8235),.q(_w_8236));
  spl2 g164_s_0(.a(n164),.q0(n164_0),.q1(n164_1));
  bfr _b_9178(.a(_w_11080),.q(n1171));
  spl2 g478_s_0(.a(n478),.q0(n478_0),.q1(_w_8123));
  and_bi g1573(.a(n1572_0),.b(n1543_0),.q(n1573));
  bfr _b_7912(.a(_w_9814),.q(_w_9815));
  bfr _b_3931(.a(_w_5833),.q(_w_5834));
  or_bb g1194(.a(n1184_0),.b(n1193_0),.q(n1194));
  bfr _b_5569(.a(_w_7471),.q(_w_7472));
  spl2 g529_s_0(.a(n529),.q0(n529_0),.q1(n529_1));
  bfr _b_4260(.a(_w_6162),.q(_w_6163));
  spl2 g817_s_0(.a(n817),.q0(n817_0),.q1(n817_1));
  spl2 g1321_s_0(.a(n1321),.q0(n1321_0),.q1(_w_12442));
  bfr _b_5012(.a(_w_6914),.q(_w_6915));
  bfr _b_14152(.a(_w_16054),.q(_w_16055));
  and_bb g864(.a(n843_1),.b(n862_1),.q(_w_8778));
  and_bi g896(.a(n895_0),.b(n832_0),.q(n896));
  spl2 g1373_s_0(.a(n1373),.q0(n1373_0),.q1(n1373_1));
  or_bb g814(.a(n713_0),.b(n813_0),.q(n814));
  bfr _b_3864(.a(_w_5766),.q(_w_5767));
  and_bi g340(.a(n298_1),.b(n338_1),.q(_w_15309));
  spl2 g320_s_0(.a(n320),.q0(n320_0),.q1(n320_1));
  spl2 g1172_s_0(.a(n1172),.q0(n1172_0),.q1(n1172_1));
  spl2 g783_s_0(.a(n783),.q0(n783_0),.q1(n783_1));
  spl2 g1838_s_0(.a(n1838),.q0(n1838_0),.q1(n1838_1));
  spl2 g643_s_0(.a(n643),.q0(n643_0),.q1(n643_1));
  spl2 g1534_s_0(.a(n1534),.q0(n1534_0),.q1(n1534_1));
  and_bb g1383(.a(N239_10),.b(N375_18),.q(_w_13544));
  bfr _b_7410(.a(_w_9312),.q(_w_9313));
  spl2 g330_s_0(.a(n330),.q0(n330_0),.q1(_w_8127));
  bfr _b_4677(.a(_w_6579),.q(_w_6580));
  bfr _b_9191(.a(_w_11093),.q(_w_11094));
  spl2 g332_s_0(.a(n332),.q0(n332_0),.q1(n332_1));
  bfr _b_8903(.a(_w_10805),.q(_w_10806));
  bfr _b_14371(.a(_w_16273),.q(_w_16274));
  spl2 g703_s_0(.a(n703),.q0(n703_0),.q1(n703_1));
  spl2 g147_s_0(.a(n147),.q0(n147_0),.q1(n147_1));
  bfr _b_4988(.a(_w_6890),.q(_w_6891));
  bfr _b_4420(.a(_w_6322),.q(n108_1));
  bfr _b_8713(.a(_w_10615),.q(_w_10616));
  spl2 g1389_s_0(.a(n1389),.q0(n1389_0),.q1(n1389_1));
  bfr _b_4595(.a(_w_6497),.q(_w_6498));
  bfr _b_4055(.a(_w_5957),.q(_w_5958));
  bfr _b_12635(.a(_w_14537),.q(_w_14538));
  and_bi g73(.a(n66_1),.b(n69_1),.q(n73));
  bfr _b_6302(.a(_w_8204),.q(n1429));
  spl2 g143_s_0(.a(n143),.q0(n143_0),.q1(n143_1));
  bfr _b_4846(.a(_w_6748),.q(_w_6749));
  spl2 g977_s_0(.a(n977),.q0(n977_0),.q1(n977_1));
  bfr _b_5019(.a(_w_6921),.q(_w_6922));
  spl2 g722_s_0(.a(n722),.q0(n722_0),.q1(n722_1));
  spl2 g1734_s_0(.a(n1734),.q0(n1734_0),.q1(n1734_1));
  bfr _b_12966(.a(_w_14868),.q(_w_14869));
  spl2 g1215_s_0(.a(n1215),.q0(n1215_0),.q1(n1215_1));
  bfr _b_7661(.a(_w_9563),.q(_w_9564));
  bfr _b_4162(.a(_w_6064),.q(_w_6065));
  spl2 g363_s_0(.a(n363),.q0(n363_0),.q1(n363_1));
  bfr _b_6052(.a(_w_7954),.q(_w_7955));
  bfr _b_13077(.a(_w_14979),.q(_w_14980));
  bfr _b_11204(.a(_w_13106),.q(_w_13107));
  spl2 g364_s_0(.a(n364),.q0(n364_0),.q1(n364_1));
  spl2 g176_s_0(.a(n176),.q0(n176_0),.q1(n176_1));
  bfr _b_4173(.a(_w_6075),.q(_w_6076));
  bfr _b_14275(.a(_w_16177),.q(_w_16178));
  bfr _b_6060(.a(_w_7962),.q(_w_7963));
  spl2 N222_s_5(.a(N222_19),.q0(_w_7575),.q1(N222_21));
  bfr _b_7642(.a(_w_9544),.q(_w_9545));
  spl2 g366_s_0(.a(n366),.q0(n366_0),.q1(n366_1));
  spl2 g648_s_0(.a(n648),.q0(n648_0),.q1(n648_1));
  bfr _b_9207(.a(_w_11109),.q(_w_11110));
  bfr _b_4053(.a(_w_5955),.q(_w_5956));
  bfr _b_12374(.a(_w_14276),.q(n1745));
  bfr _b_4993(.a(_w_6895),.q(_w_6896));
  spl2 g976_s_0(.a(n976),.q0(n976_0),.q1(n976_1));
  bfr _b_4198(.a(_w_6100),.q(N171_13));
  spl2 g986_s_0(.a(n986),.q0(n986_0),.q1(_w_8139));
  bfr _b_13355(.a(_w_15257),.q(_w_15258));
  bfr _b_6830(.a(_w_8732),.q(_w_8733));
  spl2 g130_s_0(.a(n130),.q0(n130_0),.q1(_w_8143));
  bfr _b_11831(.a(_w_13733),.q(_w_13734));
  bfr _b_11217(.a(_w_13119),.q(_w_13120));
  or_bb g1721(.a(n1719_0),.b(n1720),.q(_w_14123));
  spl2 g1347_s_0(.a(n1347),.q0(n1347_0),.q1(n1347_1));
  and_bi g1139(.a(n1137_0),.b(n1138),.q(n1139));
  bfr _b_5026(.a(_w_6928),.q(_w_6929));
  bfr _b_4443(.a(_w_6345),.q(n214_1));
  spl4L N392_s_4(.a(N392_3),.q0(N392_16),.q1(N392_17),.q2(N392_18),.q3(_w_8147));
  bfr _b_12572(.a(_w_14474),.q(_w_14475));
  or_bb g248(.a(n191_1),.b(n247_0),.q(_w_8151));
  bfr _b_3903(.a(_w_5805),.q(_w_5806));
  and_bi g1133(.a(n1131_0),.b(n1132),.q(n1133));
  spl2 g1199_s_0(.a(n1199),.q0(n1199_0),.q1(n1199_1));
  spl4L N341_s_1(.a(N341_0),.q0(N341_4),.q1(N341_5),.q2(N341_6),.q3(N341_7));
  and_bi g1780(.a(n1759_1),.b(n1762_1),.q(n1780));
  bfr _b_14167(.a(_w_16069),.q(_w_16070));
  bfr _b_11121(.a(_w_13023),.q(_w_13024));
  bfr _b_4674(.a(_w_6576),.q(_w_6577));
  bfr _b_13798(.a(_w_15700),.q(_w_15701));
  and_bi g1744(.a(n1743_0),.b(n1738_0),.q(n1744));
  bfr _b_9775(.a(_w_11677),.q(_w_11678));
  and_bi g1343(.a(n1272_1),.b(n1341_1),.q(_w_13431));
  bfr _b_6504(.a(_w_8406),.q(_w_8407));
  bfr _b_10139(.a(_w_12041),.q(_w_12042));
  bfr _b_3862(.a(_w_5764),.q(_w_5765));
  and_bi g1347(.a(n1345_0),.b(n1346),.q(n1347));
  bfr _b_3555(.a(_w_5457),.q(_w_5458));
  and_bi g1669(.a(n1606_1),.b(n1667_1),.q(_w_8153));
  or_bb g1039(.a(n1037_0),.b(n1038),.q(n1039));
  bfr _b_3664(.a(_w_5566),.q(_w_5567));
  bfr _b_8326(.a(_w_10228),.q(_w_10229));
  and_bb g607(.a(n521_1),.b(n605_1),.q(_w_8154));
  bfr _b_13298(.a(_w_15200),.q(_w_15201));
  spl2 g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1));
  and_bi g613(.a(n606_1),.b(n609_1),.q(n613));
  bfr _b_9914(.a(_w_11816),.q(_w_11817));
  bfr _b_4291(.a(_w_6193),.q(_w_6194));
  spl2 g846_s_0(.a(n846),.q0(n846_0),.q1(n846_1));
  spl2 g1291_s_0(.a(n1291),.q0(n1291_0),.q1(_w_9562));
  bfr _b_14178(.a(_w_16080),.q(_w_16081));
  bfr _b_10351(.a(_w_12253),.q(_w_12254));
  spl4L N528_s_2(.a(N528_1),.q0(N528_8),.q1(N528_9),.q2(N528_10),.q3(N528_11));
  or_bb g1119(.a(n1061_0),.b(n1118_0),.q(n1119));
  or_bb g1552(.a(n1550_0),.b(n1551_0),.q(n1552));
  bfr _b_7717(.a(_w_9619),.q(_w_9620));
  bfr _b_13755(.a(_w_15657),.q(_w_15658));
  bfr _b_8958(.a(_w_10860),.q(_w_10861));
  spl2 g181_s_0(.a(n181),.q0(n181_0),.q1(n181_1));
  and_bb g1114(.a(n1063_1),.b(n1112_1),.q(_w_8179));
  bfr _b_6296(.a(_w_8198),.q(n1123));
  or_bb g1113(.a(n1063_0),.b(n1112_0),.q(n1113));
  and_bi g1244(.a(n1242_0),.b(n1243),.q(n1244));
  and_bb g1108(.a(n1065_1),.b(n1106_1),.q(_w_8180));
  or_bb g173(.a(n171_0),.b(n172),.q(n173));
  bfr _b_5289(.a(_w_7191),.q(_w_7192));
  and_bi g260(.a(n242_1),.b(n258_1),.q(_w_8181));
  bfr _b_9721(.a(_w_11623),.q(n1254_1));
  bfr _b_14266(.a(_w_16168),.q(_w_16169));
  bfr _b_7362(.a(_w_9264),.q(_w_9265));
  or_bb g1106(.a(n1104_0),.b(n1105),.q(n1106));
  and_bi g1123(.a(n1060_1),.b(n1121_1),.q(_w_8198));
  bfr _b_3748(.a(_w_5650),.q(_w_5651));
  bfr _b_6212(.a(_w_8114),.q(_w_8115));
  bfr _b_6654(.a(_w_8556),.q(_w_8557));
  bfr _b_6349(.a(_w_8251),.q(_w_8252));
  bfr _b_8989(.a(_w_10891),.q(_w_10892));
  bfr _b_8658(.a(_w_10560),.q(n163));
  bfr _b_10514(.a(_w_12416),.q(_w_12417));
  bfr _b_4217(.a(_w_6119),.q(_w_6120));
  and_bi g1093(.a(n1070_1),.b(n1091_1),.q(_w_8200));
  bfr _b_3647(.a(_w_5549),.q(_w_5550));
  and_bi g625(.a(n570_1),.b(n573_1),.q(n625));
  and_bb g1739(.a(N256_10),.b(N443_19),.q(_w_8731));
  and_bi g1092(.a(n1091_0),.b(n1070_0),.q(n1092));
  bfr _b_13908(.a(_w_15810),.q(_w_15811));
  bfr _b_3690(.a(_w_5592),.q(_w_5593));
  or_bb g1089(.a(n1071_0),.b(n1088_0),.q(n1089));
  or_bb g587(.a(n585_0),.b(n586),.q(n587));
  and_bi g198(.a(n196_0),.b(n197),.q(n198));
  bfr _b_3540(.a(_w_5442),.q(_w_5443));
  bfr _b_13334(.a(_w_15236),.q(_w_15237));
  bfr _b_12109(.a(_w_14011),.q(_w_14012));
  bfr _b_7667(.a(_w_9569),.q(_w_9570));
  spl2 g1021_s_0(.a(n1021),.q0(n1021_0),.q1(n1021_1));
  bfr _b_14299(.a(_w_16201),.q(_w_16202));
  and_bi g947(.a(n893_1),.b(n896_1),.q(n947));
  and_bb g1660(.a(n1609_1),.b(n1658_1),.q(_w_8203));
  bfr _b_3893(.a(_w_5795),.q(_w_5796));
  spl2 g49_s_0(.a(n49),.q0(n49_0),.q1(n49_1));
  bfr _b_11618(.a(_w_13520),.q(n1369));
  and_bi g1168(.a(n1131_1),.b(n1134_1),.q(n1168));
  bfr _b_8678(.a(_w_10580),.q(_w_10581));
  bfr _b_4157(.a(_w_6059),.q(_w_6060));
  and_bb g1429(.a(n1370_1),.b(n1427_1),.q(_w_8204));
  spl2 g904_s_0(.a(n904),.q0(n904_0),.q1(n904_1));
  bfr _b_4559(.a(_w_6461),.q(N154_15));
  bfr _b_12627(.a(_w_14529),.q(_w_14530));
  spl2 g375_s_0(.a(n375),.q0(n375_0),.q1(n375_1));
  bfr _b_6980(.a(_w_8882),.q(_w_8883));
  spl2 g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1));
  and_bi g1081(.a(n1074_1),.b(n1079_1),.q(_w_8205));
  bfr _b_9274(.a(_w_11176),.q(_w_11177));
  bfr _b_11635(.a(_w_13537),.q(_w_13538));
  bfr _b_4159(.a(_w_6061),.q(_w_6062));
  bfr _b_9713(.a(_w_11615),.q(_w_11616));
  spl2 g1625_s_0(.a(n1625),.q0(n1625_0),.q1(n1625_1));
  spl2 g1171_s_0(.a(n1171),.q0(n1171_0),.q1(n1171_1));
  bfr _b_4180(.a(_w_6082),.q(_w_6083));
  and_bb g1549(.a(N239_12),.b(N409_18),.q(n1549));
  bfr _b_12994(.a(_w_14896),.q(_w_14897));
  spl2 g1479_s_0(.a(n1479),.q0(n1479_0),.q1(_w_13934));
  bfr _b_5424(.a(_w_7326),.q(_w_7327));
  bfr _b_8322(.a(_w_10224),.q(_w_10225));
  bfr _b_13988(.a(_w_15890),.q(_w_15891));
  and_bb g184(.a(N35_9),.b(N358_6),.q(_w_8208));
  bfr _b_3409(.a(_w_5311),.q(_w_5312));
  bfr _b_6939(.a(_w_8841),.q(_w_8842));
  spl2 g917_s_0(.a(n917),.q0(n917_0),.q1(_w_8216));
  bfr _b_8254(.a(_w_10156),.q(_w_10157));
  and_bi g1293(.a(n1291_0),.b(n1292),.q(n1293));
  bfr _b_10315(.a(_w_12217),.q(_w_12218));
  bfr _b_4185(.a(_w_6087),.q(_w_6088));
  bfr _b_12959(.a(_w_14861),.q(_w_14862));
  and_bb g1066(.a(N171_11),.b(N392_14),.q(n1066));
  bfr _b_12662(.a(_w_14564),.q(n1824));
  and_bi g1065(.a(n992_1),.b(n995_1),.q(n1065));
  bfr _b_5403(.a(_w_7305),.q(_w_7306));
  spl2 g1077_s_0(.a(n1077),.q0(n1077_0),.q1(_w_8220));
  bfr _b_11919(.a(_w_13821),.q(_w_13822));
  bfr _b_4949(.a(_w_6851),.q(_w_6852));
  bfr _b_6682(.a(_w_8584),.q(_w_8585));
  bfr _b_4256(.a(_w_6158),.q(_w_6159));
  bfr _b_10538(.a(_w_12440),.q(_w_12441));
  bfr _b_9133(.a(_w_11035),.q(_w_11036));
  bfr _b_9971(.a(_w_11873),.q(_w_11874));
  and_bi g187(.a(n156_1),.b(n159_1),.q(n187));
  and_bi g1294(.a(n1293_0),.b(n1288_0),.q(n1294));
  and_bi g1053(.a(n1028_1),.b(n1031_1),.q(n1053));
  and_bb g1468(.a(N222_12),.b(N409_17),.q(n1468));
  bfr _b_6804(.a(_w_8706),.q(_w_8707));
  bfr _b_9610(.a(_w_11512),.q(_w_11513));
  or_bb g1398(.a(n1380_0),.b(n1397_0),.q(n1398));
  and_bi g322(.a(n304_1),.b(n320_1),.q(_w_8228));
  bfr _b_13120(.a(_w_15022),.q(_w_15023));
  bfr _b_3536(.a(_w_5438),.q(_w_5439));
  and_bi g1051(.a(n1034_1),.b(n1037_1),.q(n1051));
  bfr _b_12851(.a(_w_14753),.q(_w_14754));
  bfr _b_12651(.a(_w_14553),.q(_w_14554));
  spl2 g505_s_0(.a(n505),.q0(n505_0),.q1(n505_1));
  bfr _b_4881(.a(_w_6783),.q(_w_6784));
  and_bb g1062(.a(N137_13),.b(N426_12),.q(n1062));
  and_bb g1050(.a(N35_19),.b(N528_6),.q(_w_8273));
  bfr _b_5382(.a(_w_7284),.q(_w_7285));
  bfr _b_3843(.a(_w_5745),.q(_w_5746));
  and_bi g1190(.a(n1188_0),.b(n1189),.q(_w_8297));
  and_bi g1049(.a(n1040_1),.b(n1043_1),.q(n1049));
  and_bb g401(.a(n371_1),.b(n399_1),.q(_w_10201));
  bfr _b_4600(.a(_w_6502),.q(_w_6503));
  and_bb g520(.a(N1_16),.b(N477_4),.q(n520));
  and_bi g1048(.a(n1047),.b(n1046_0),.q(_w_8300));
  bfr _b_8441(.a(_w_10343),.q(_w_10344));
  or_bb g1045(.a(n1043_0),.b(n1044),.q(_w_8354));
  spl4L N137_s_2(.a(N137_1),.q0(N137_8),.q1(N137_9),.q2(N137_10),.q3(_w_8833));
  and_bi g1037(.a(n1036_0),.b(n938_0),.q(n1037));
  bfr _b_9065(.a(_w_10967),.q(_w_10968));
  spl2 g538_s_0(.a(n538),.q0(n538_0),.q1(n538_1));
  bfr _b_4726(.a(_w_6628),.q(_w_6629));
  and_bi g1026(.a(n942_1),.b(n1024_1),.q(_w_8356));
  bfr _b_9696(.a(_w_11598),.q(n392));
  bfr _b_4380(.a(_w_6282),.q(_w_6283));
  or_bb g875(.a(n839_0),.b(n874_0),.q(n875));
  spl2 g831_s_0(.a(n831),.q0(n831_0),.q1(n831_1));
  bfr _b_4015(.a(_w_5917),.q(_w_5918));
  and_bi g1442(.a(n1440_0),.b(n1441),.q(n1442));
  and_bb g1630(.a(n1619_1),.b(n1628_1),.q(_w_9161));
  and_bb g54(.a(N18_6),.b(N307_5),.q(_w_12067));
  bfr _b_13935(.a(_w_15837),.q(_w_15838));
  and_bb g701(.a(n615_1),.b(n699_1),.q(_w_9291));
  bfr _b_4821(.a(_w_6723),.q(_w_6724));
  and_bi g283(.a(n282_0),.b(n234_0),.q(n283));
  bfr _b_13451(.a(_w_15353),.q(_w_15354));
  and_bb g1865(.a(n1854_1),.b(n1863_1),.q(_w_8358));
  bfr _b_4424(.a(_w_6326),.q(_w_6327));
  bfr _b_9327(.a(_w_11229),.q(_w_11230));
  bfr _b_11746(.a(_w_13648),.q(_w_13649));
  bfr _b_4156(.a(_w_6058),.q(_w_6059));
  bfr _b_13044(.a(_w_14946),.q(n1887_1));
  spl2 g63_s_0(.a(n63),.q0(n63_0),.q1(n63_1));
  bfr _b_12886(.a(_w_14788),.q(_w_14789));
  and_bi g691(.a(n690_0),.b(n618_0),.q(n691));
  bfr _b_8807(.a(_w_10709),.q(_w_10710));
  or_bb g991(.a(n989_0),.b(n990),.q(n991));
  bfr _b_3856(.a(_w_5758),.q(_w_5759));
  bfr _b_3441(.a(_w_5343),.q(_w_5344));
  spl2 g139_s_0(.a(n139),.q0(n139_0),.q1(n139_1));
  bfr _b_8710(.a(_w_10612),.q(_w_10613));
  bfr _b_11907(.a(_w_13809),.q(_w_13810));
  spl2 g1439_s_0(.a(n1439),.q0(n1439_0),.q1(n1439_1));
  bfr _b_5669(.a(_w_7571),.q(_w_7572));
  bfr _b_13397(.a(_w_15299),.q(n56_2));
  and_bb g624(.a(N103_11),.b(N392_10),.q(n624));
  bfr _b_8524(.a(_w_10426),.q(_w_10427));
  spl2 g1773_s_0(.a(n1773),.q0(n1773_0),.q1(n1773_1));
  and_bi g1639(.a(n1616_1),.b(n1637_1),.q(_w_13582));
  bfr _b_5725(.a(_w_7627),.q(_w_7628));
  spl2 g501_s_0(.a(n501),.q0(n501_0),.q1(n501_1));
  or_bb g1010(.a(n1009_0),.b(n947_0),.q(n1010));
  bfr _b_12985(.a(_w_14887),.q(_w_14888));
  bfr _b_8687(.a(_w_10589),.q(_w_10590));
  and_bi g1337(.a(n1274_1),.b(n1335_1),.q(_w_13425));
  spl2 g1241_s_0(.a(n1241),.q0(n1241_0),.q1(n1241_1));
  and_bi g1002(.a(n950_1),.b(n1000_1),.q(_w_8362));
  spl2 g129_s_0(.a(n129),.q0(n129_0),.q1(n129_1));
  and_bi g1128(.a(n1127_0),.b(n1058_0),.q(n1128));
  spl2 g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1));
  bfr _b_13076(.a(_w_14978),.q(_w_14979));
  and_bb g999(.a(n951_1),.b(n997_1),.q(_w_8363));
  and_bi g567(.a(n566_0),.b(n534_0),.q(n567));
  or_bb g967(.a(n965_0),.b(n966),.q(_w_8370));
  spl2 g1599_s_0(.a(n1599),.q0(n1599_0),.q1(n1599_1));
  bfr _b_7978(.a(_w_9880),.q(_w_9881));
  spl4L N528_s_1(.a(N528_0),.q0(N528_4),.q1(N528_5),.q2(N528_6),.q3(N528_7));
  bfr _b_10365(.a(_w_12267),.q(_w_12268));
  and_bb g858(.a(n845_1),.b(n856_1),.q(_w_9363));
  spl2 g448_s_0(.a(n448),.q0(n448_0),.q1(n448_1));
  bfr _b_6181(.a(_w_8083),.q(_w_8084));
  bfr _b_13568(.a(_w_15470),.q(_w_15471));
  and_bb g964(.a(N239_6),.b(N307_18),.q(_w_8381));
  bfr _b_4149(.a(_w_6051),.q(_w_6052));
  and_bb g962(.a(N256_20),.b(N290_19),.q(n962));
  and_bi g825(.a(n802_1),.b(n805_1),.q(n825));
  spl2 g1637_s_0(.a(n1637),.q0(n1637_0),.q1(n1637_1));
  spl2 g679_s_0(.a(n679),.q0(n679_0),.q1(n679_1));
  bfr _b_12532(.a(_w_14434),.q(_w_14435));
  spl2 g1860_s_0(.a(n1860),.q0(n1860_0),.q1(n1860_1));
  bfr _b_4735(.a(_w_6637),.q(_w_6638));
  and_bi g867(.a(n842_1),.b(n865_1),.q(_w_8776));
  bfr _b_11292(.a(_w_13194),.q(_w_13195));
  spl2 g1684_s_0(.a(n1684),.q0(n1684_0),.q1(n1684_1));
  bfr _b_9566(.a(_w_11468),.q(_w_11469));
  spl2 g593_s_0(.a(n593),.q0(n593_0),.q1(n593_1));
  bfr _b_7855(.a(_w_9757),.q(_w_9758));
  and_bb g958(.a(N205_8),.b(N341_16),.q(n958));
  bfr _b_10798(.a(_w_12700),.q(_w_12701));
  spl2 g1440_s_0(.a(n1440),.q0(n1440_0),.q1(_w_8385));
  bfr _b_10718(.a(_w_12620),.q(_w_12621));
  bfr _b_4417(.a(_w_6319),.q(_w_6320));
  bfr _b_8559(.a(_w_10461),.q(_w_10462));
  bfr _b_8793(.a(_w_10695),.q(_w_10696));
  and_bi g290(.a(n232_1),.b(n288_1),.q(_w_8390));
  bfr _b_8244(.a(_w_10146),.q(_w_10147));
  bfr _b_7508(.a(_w_9410),.q(_w_9411));
  and_bi g949(.a(n887_1),.b(n890_1),.q(n949));
  bfr _b_13590(.a(_w_15492),.q(_w_15493));
  bfr _b_11233(.a(_w_13135),.q(_w_13136));
  and_bi g1099(.a(n1068_1),.b(n1097_1),.q(_w_8559));
  and_bi g437(.a(n430_1),.b(n433_1),.q(n437));
  bfr _b_3693(.a(_w_5595),.q(_w_5596));
  bfr _b_7048(.a(_w_8950),.q(n1322));
  bfr _b_11081(.a(_w_12983),.q(_w_12984));
  bfr _b_10053(.a(_w_11955),.q(_w_11956));
  or_bb g789(.a(n787_0),.b(n788),.q(n789));
  bfr _b_4900(.a(_w_6802),.q(_w_6803));
  and_bi g941(.a(n911_1),.b(n914_1),.q(n941));
  and_bi g963(.a(n962_0),.b(n739_1),.q(n963));
  bfr _b_3649(.a(_w_5551),.q(_w_5552));
  bfr _b_4817(.a(_w_6719),.q(_w_6720));
  bfr _b_8580(.a(_w_10482),.q(_w_10483));
  and_bb g1516(.a(n1457_1),.b(n1514_1),.q(_w_11017));
  and_bi g729(.a(n658_1),.b(n661_1),.q(n729));
  bfr _b_7385(.a(_w_9287),.q(_w_9288));
  bfr _b_4723(.a(_w_6625),.q(_w_6626));
  bfr _b_4255(.a(_w_6157),.q(_w_6158));
  and_bi g935(.a(n929_1),.b(n932_1),.q(_w_8619));
  bfr _b_9825(.a(_w_11727),.q(_w_11728));
  and_bi g932(.a(n931_0),.b(n820_0),.q(n932));
  bfr _b_10632(.a(_w_12534),.q(_w_12535));
  and_bb g797(.a(n719_1),.b(n795_1),.q(_w_8943));
  bfr _b_6175(.a(_w_8077),.q(_w_8078));
  bfr _b_12211(.a(_w_14113),.q(n1690));
  spl4L N222_s_3(.a(N222_2),.q0(_w_8621),.q1(N222_13),.q2(_w_8677),.q3(_w_8701));
  and_bi g931(.a(n929_0),.b(n930),.q(n931));
  spl4L N154_s_2(.a(N154_1),.q0(N154_8),.q1(N154_9),.q2(N154_10),.q3(_w_7547));
  bfr _b_4795(.a(_w_6697),.q(n192_2));
  bfr _b_4531(.a(_w_6433),.q(_w_6434));
  bfr _b_9203(.a(_w_11105),.q(_w_11106));
  and_bb g1237(.a(n1170_1),.b(n1235_1),.q(_w_8726));
  and_bi g1013(.a(n1012_0),.b(n946_0),.q(n1013));
  spl2 g1674_s_0(.a(n1674),.q0(n1674_0),.q1(n1674_1));
  bfr _b_5002(.a(_w_6904),.q(_w_6905));
  and_bi g927(.a(n822_1),.b(n925_1),.q(_w_8727));
  spl4L N188_s_4(.a(N188_3),.q0(N188_16),.q1(N188_17),.q2(N188_18),.q3(N188_19));
  and_bb g1078(.a(n1075_1),.b(n1076_1),.q(_w_8728));
  bfr _b_9480(.a(_w_11382),.q(_w_11383));
  and_bi g1262(.a(n1260_0),.b(n1261),.q(n1262));
  bfr _b_9770(.a(_w_11672),.q(_w_11673));
  spl2 g621_s_0(.a(n621),.q0(n621_0),.q1(n621_1));
  bfr _b_12908(.a(_w_14810),.q(_w_14811));
  bfr _b_9738(.a(_w_11640),.q(_w_11641));
  bfr _b_10743(.a(_w_12645),.q(_w_12646));
  bfr _b_10425(.a(_w_12327),.q(_w_12328));
  and_bi g921(.a(n824_1),.b(n919_1),.q(_w_8729));
  bfr _b_13533(.a(_w_15435),.q(_w_15436));
  bfr _b_7498(.a(_w_9400),.q(_w_9401));
  bfr _b_7143(.a(_w_9045),.q(_w_9046));
  or_bb g916(.a(n914_0),.b(n915),.q(n916));
  or_bb g466(.a(n453_0),.b(n465_0),.q(n466));
  and_bb g100(.a(N1_9),.b(N358_4),.q(_w_8740));
  and_bi g913(.a(n911_0),.b(n912),.q(n913));
  bfr _b_10499(.a(_w_12401),.q(_w_12402));
  spl2 g821_s_0(.a(n821),.q0(n821_0),.q1(n821_1));
  bfr _b_8103(.a(_w_10005),.q(_w_10006));
  bfr _b_4901(.a(_w_6803),.q(_w_6804));
  and_bb g732(.a(N171_8),.b(N341_14),.q(n732));
  bfr _b_12586(.a(_w_14488),.q(_w_14489));
  and_bi g901(.a(n899_0),.b(n900),.q(n901));
  bfr _b_6109(.a(_w_8011),.q(_w_8012));
  or_bb g1137(.a(n1055_0),.b(n1136_0),.q(n1137));
  bfr _b_4202(.a(_w_6104),.q(_w_6105));
  bfr _b_6424(.a(_w_8326),.q(_w_8327));
  and_bi g721(.a(n682_1),.b(n685_1),.q(n721));
  bfr _b_5133(.a(_w_7035),.q(_w_7036));
  bfr _b_5533(.a(_w_7435),.q(_w_7436));
  bfr _b_7440(.a(_w_9342),.q(n1623_1));
  bfr _b_7931(.a(_w_9833),.q(_w_9834));
  or_bb g899(.a(n831_0),.b(n898_0),.q(n899));
  and_bb g838(.a(N154_10),.b(N375_13),.q(_w_8749));
  bfr _b_14149(.a(_w_16051),.q(_w_16052));
  bfr _b_5764(.a(_w_7666),.q(_w_7667));
  and_bb g846(.a(N222_20),.b(N307_17),.q(_w_8765));
  bfr _b_3849(.a(_w_5751),.q(_w_5752));
  and_bi g505(.a(n504_0),.b(n440_0),.q(n505));
  bfr _b_7257(.a(_w_9159),.q(_w_9160));
  bfr _b_14123(.a(_w_16025),.q(_w_16026));
  and_bi g897(.a(n832_1),.b(n895_1),.q(_w_8771));
  and_bi g1465(.a(n1404_1),.b(n1407_1),.q(n1465));
  bfr _b_5060(.a(_w_6962),.q(_w_6963));
  bfr _b_13893(.a(_w_15795),.q(_w_15796));
  bfr _b_9880(.a(_w_11782),.q(_w_11783));
  bfr _b_8542(.a(_w_10444),.q(_w_10445));
  and_bi g885(.a(n836_1),.b(n883_1),.q(_w_8772));
  and_bi g884(.a(n883_0),.b(n836_0),.q(n884));
  or_bb g112(.a(n111_0),.b(n78_1),.q(n112));
  bfr _b_9671(.a(_w_11573),.q(_w_11574));
  and_bb g1070(.a(N205_9),.b(N358_16),.q(_w_10443));
  or_bb g1497(.a(n1463_0),.b(n1496_0),.q(n1497));
  spl2 g1680_s_0(.a(n1680),.q0(n1680_0),.q1(n1680_1));
  bfr _b_5609(.a(_w_7511),.q(_w_7512));
  bfr _b_7026(.a(_w_8928),.q(_w_8929));
  and_bi g1301(.a(n1286_1),.b(n1299_1),.q(_w_8773));
  and_bi g367(.a(n336_1),.b(n339_1),.q(n367));
  bfr _b_8323(.a(_w_10225),.q(_w_10226));
  or_bb g1107(.a(n1065_0),.b(n1106_0),.q(n1107));
  bfr _b_7285(.a(_w_9187),.q(_w_9188));
  and_bi g1036(.a(n1034_0),.b(n1035),.q(n1036));
  bfr _b_4574(.a(_w_6476),.q(_w_6477));
  and_bi g1240(.a(n1169_1),.b(n1238_1),.q(_w_8775));
  bfr _b_14222(.a(_w_16124),.q(_w_16125));
  and_bi g872(.a(n871_0),.b(n840_0),.q(n872));
  bfr _b_4022(.a(_w_5924),.q(_w_5925));
  bfr _b_6439(.a(_w_8341),.q(_w_8342));
  bfr _b_10154(.a(_w_12056),.q(_w_12057));
  spl2 g1173_s_0(.a(n1173),.q0(n1173_0),.q1(n1173_1));
  and_bb g1132(.a(n1057_1),.b(n1130_1),.q(_w_8152));
  and_bb g131(.a(n101_1),.b(n129_1),.q(_w_8777));
  bfr _b_10272(.a(_w_12174),.q(_w_12175));
  spl2 g453_s_0(.a(n453),.q0(n453_0),.q1(n453_1));
  spl2 g1006_s_0(.a(n1006),.q0(n1006_0),.q1(n1006_1));
  or_bb g1440(.a(n1366_0),.b(n1439_0),.q(n1440));
  bfr _b_6716(.a(_w_8618),.q(n936));
  spl2 g1870_s_0(.a(n1870),.q0(n1870_0),.q1(_w_8781));
  and_bi g860(.a(n859_0),.b(n844_0),.q(n860));
  bfr _b_6907(.a(_w_8809),.q(_w_8810));
  and_bi g579(.a(n578_0),.b(n530_0),.q(n579));
  bfr _b_3962(.a(_w_5864),.q(_w_5865));
  bfr _b_9933(.a(_w_11835),.q(n899_1));
  spl2 g832_s_0(.a(n832),.q0(n832_0),.q1(n832_1));
  spl2 g543_s_0(.a(n543),.q0(n543_0),.q1(n543_1));
  spl2 g324_s_0(.a(n324),.q0(n324_0),.q1(_w_8789));
  bfr _b_13789(.a(_w_15691),.q(_w_15692));
  spl2 g1341_s_0(.a(n1341),.q0(n1341_0),.q1(n1341_1));
  and_bb g844(.a(N205_7),.b(N324_16),.q(_w_8793));
  bfr _b_7309(.a(_w_9211),.q(_w_9212));
  and_bb g842(.a(N188_8),.b(N341_15),.q(n842));
  bfr _b_5150(.a(_w_7052),.q(_w_7053));
  bfr _b_3454(.a(_w_5356),.q(_w_5357));
  bfr _b_5367(.a(_w_7269),.q(_w_7270));
  spl2 g1211_s_0(.a(n1211),.q0(n1211_0),.q1(n1211_1));
  bfr _b_13502(.a(_w_15404),.q(_w_15405));
  and_bb g836(.a(N137_11),.b(N392_12),.q(n836));
  and_bi g833(.a(n778_1),.b(n781_1),.q(n833));
  bfr _b_11444(.a(_w_13346),.q(n1319));
  or_bb g1832(.a(n1830_0),.b(n1831),.q(n1832));
  bfr _b_6185(.a(_w_8087),.q(_w_8088));
  and_bb g1636(.a(n1617_1),.b(n1634_1),.q(_w_8808));
  bfr _b_14075(.a(_w_15977),.q(_w_15978));
  bfr _b_13665(.a(_w_15567),.q(_w_15568));
  bfr _b_12646(.a(_w_14548),.q(_w_14549));
  and_bi g199(.a(n198_0),.b(n190_0),.q(n199));
  bfr _b_10258(.a(_w_12160),.q(_w_12161));
  bfr _b_6544(.a(_w_8446),.q(_w_8447));
  or_bb g819(.a(n817_0),.b(n818),.q(_w_8857));
  bfr _b_11207(.a(_w_13109),.q(_w_13110));
  spl2 g733_s_0(.a(n733),.q0(n733_0),.q1(n733_1));
  bfr _b_12128(.a(_w_14030),.q(_w_14031));
  bfr _b_7418(.a(_w_9320),.q(_w_9321));
  bfr _b_11541(.a(_w_13443),.q(_w_13444));
  and_bi g810(.a(n808_0),.b(n809),.q(n810));
  or_bb g1224(.a(n1174_0),.b(n1223_0),.q(n1224));
  bfr _b_4171(.a(_w_6073),.q(_w_6074));
  bfr _b_13979(.a(_w_15881),.q(_w_15882));
  bfr _b_3735(.a(_w_5637),.q(_w_5638));
  bfr _b_9337(.a(_w_11239),.q(_w_11240));
  or_bb g1484(.a(n1482_0),.b(n1483),.q(n1484));
  and_bb g803(.a(n717_1),.b(n801_1),.q(_w_8926));
  spl2 g1487_s_0(.a(n1487),.q0(n1487_0),.q1(n1487_1));
  and_bi g1071(.a(n974_1),.b(n977_1),.q(n1071));
  spl2 g1251_s_0(.a(n1251),.q0(n1251_0),.q1(n1251_1));
  bfr _b_10003(.a(_w_11905),.q(_w_11906));
  spl2 g514_s_0(.a(n514),.q0(n514_0),.q1(_w_8939));
  bfr _b_12820(.a(_w_14722),.q(_w_14723));
  bfr _b_6142(.a(_w_8044),.q(_w_8045));
  bfr _b_14172(.a(_w_16074),.q(_w_16075));
  bfr _b_7479(.a(_w_9381),.q(_w_9382));
  and_bi g1025(.a(n1024_0),.b(n942_0),.q(n1025));
  bfr _b_12166(.a(_w_14068),.q(_w_14069));
  spl2 g1415_s_0(.a(n1415),.q0(n1415_0),.q1(n1415_1));
  bfr _b_9056(.a(_w_10958),.q(_w_10959));
  bfr _b_11864(.a(_w_13766),.q(_w_13767));
  or_bb g796(.a(n719_0),.b(n795_0),.q(n796));
  bfr _b_8081(.a(_w_9983),.q(_w_9984));
  bfr _b_3479(.a(_w_5381),.q(_w_5382));
  bfr _b_6822(.a(_w_8724),.q(N222_15));
  bfr _b_7182(.a(_w_9084),.q(_w_9085));
  bfr _b_11238(.a(_w_13140),.q(_w_13141));
  bfr _b_5776(.a(_w_7678),.q(_w_7679));
  spl2 g274_s_0(.a(n274),.q0(n274_0),.q1(_w_8944));
  and_bi g794(.a(n720_1),.b(n792_1),.q(_w_8948));
  bfr _b_5841(.a(_w_7743),.q(_w_7744));
  spl2 g953_s_0(.a(n953),.q0(n953_0),.q1(n953_1));
  spl2 g716_s_0(.a(n716),.q0(n716_0),.q1(n716_1));
  bfr _b_8645(.a(_w_10547),.q(_w_10548));
  and_bi g470(.a(n452_1),.b(n468_1),.q(_w_8949));
  or_bb g1827(.a(n1825_0),.b(n1826_0),.q(n1827));
  and_bi g1406(.a(n1404_0),.b(n1405),.q(n1406));
  bfr _b_6650(.a(_w_8552),.q(_w_8553));
  bfr _b_4307(.a(_w_6209),.q(_w_6210));
  spl2 g594_s_0(.a(n594),.q0(n594_0),.q1(_w_8119));
  bfr _b_4464(.a(_w_6366),.q(_w_6367));
  or_bb g790(.a(n721_0),.b(n789_0),.q(n790));
  and_bi g204(.a(n202_0),.b(n203),.q(n204));
  bfr _b_14187(.a(_w_16089),.q(_w_16090));
  spl2 g433_s_0(.a(n433),.q0(n433_0),.q1(n433_1));
  and_bi g817(.a(n816_0),.b(n712_0),.q(n817));
  bfr _b_6096(.a(_w_7998),.q(_w_7999));
  bfr _b_3545(.a(_w_5447),.q(_w_5448));
  spl2 g599_s_0(.a(n599),.q0(n599_0),.q1(n599_1));
  bfr _b_6308(.a(_w_8210),.q(_w_8211));
  or_bb g1338(.a(n1336_0),.b(n1337),.q(n1338));
  bfr _b_7719(.a(_w_9621),.q(n894));
  bfr _b_13487(.a(_w_15389),.q(_w_15390));
  bfr _b_3839(.a(_w_5741),.q(_w_5742));
  and_bi g786(.a(n784_0),.b(n785),.q(n786));
  and_bi g1849(.a(n1818_1),.b(n1847_1),.q(_w_11133));
  bfr _b_11439(.a(_w_13341),.q(_w_13342));
  bfr _b_4626(.a(_w_6528),.q(_w_6529));
  and_bb g1367(.a(N103_18),.b(N511_10),.q(_w_13496));
  bfr _b_8003(.a(_w_9905),.q(_w_9906));
  spl2 g1230_s_0(.a(n1230),.q0(n1230_0),.q1(_w_8951));
  and_bi g965(.a(n963_0),.b(n964_0),.q(n965));
  bfr _b_4117(.a(_w_6019),.q(_w_6020));
  bfr _b_9654(.a(_w_11556),.q(_w_11557));
  spl2 g43_s_0(.a(n43),.q0(n43_0),.q1(n43_1));
  bfr _b_4072(.a(_w_5974),.q(_w_5975));
  and_bi g252(.a(n250_0),.b(n251),.q(n252));
  and_bi g1837(.a(n1822_1),.b(n1835_1),.q(_w_14572));
  bfr _b_7477(.a(_w_9379),.q(_w_9380));
  bfr _b_7424(.a(_w_9326),.q(_w_9327));
  and_bi g782(.a(n724_1),.b(n780_1),.q(_w_8955));
  and_bb g830(.a(N443_9),.b(N86_14),.q(_w_8956));
  or_bb g783(.a(n781_0),.b(n782),.q(n783));
  bfr _b_3891(.a(_w_5793),.q(_w_5794));
  and_bi g780(.a(n778_0),.b(n779),.q(n780));
  bfr _b_6323(.a(_w_8225),.q(_w_8226));
  spl2 g602_s_0(.a(n602),.q0(n602_0),.q1(n602_1));
  bfr _b_4728(.a(_w_6630),.q(_w_6631));
  bfr _b_4693(.a(_w_6595),.q(_w_6596));
  bfr _b_4401(.a(_w_6303),.q(n564_1));
  bfr _b_8033(.a(_w_9935),.q(_w_9936));
  bfr _b_12148(.a(_w_14050),.q(_w_14051));
  bfr _b_10846(.a(_w_12748),.q(_w_12749));
  bfr _b_8814(.a(_w_10716),.q(_w_10717));
  bfr _b_6591(.a(_w_8493),.q(_w_8494));
  bfr _b_9319(.a(_w_11221),.q(_w_11222));
  and_bi g573(.a(n572_0),.b(n532_0),.q(n573));
  and_bi g1117(.a(n1062_1),.b(n1115_1),.q(_w_8960));
  bfr _b_9321(.a(_w_11223),.q(_w_11224));
  spl4L N188_s_0(.a(_w_15531),.q0(N188_0),.q1(_w_8961),.q2(_w_8985),.q3(_w_9041));
  bfr _b_3451(.a(_w_5353),.q(_w_5354));
  bfr _b_7136(.a(_w_9038),.q(_w_9039));
  or_bb g1628(.a(n1626_0),.b(n1627),.q(n1628));
  spl2 g101_s_0(.a(n101),.q0(n101_0),.q1(n101_1));
  bfr _b_12722(.a(_w_14624),.q(_w_14625));
  bfr _b_4063(.a(_w_5965),.q(_w_5966));
  and_bi g776(.a(n726_1),.b(n774_1),.q(_w_9129));
  bfr _b_5561(.a(_w_7463),.q(_w_7464));
  bfr _b_6735(.a(_w_8637),.q(_w_8638));
  spl2 g1391_s_0(.a(n1391),.q0(n1391_0),.q1(n1391_1));
  bfr _b_10897(.a(_w_12799),.q(_w_12800));
  spl2 g1385_s_0(.a(n1385),.q0(n1385_0),.q1(n1385_1));
  and_bi g1728(.a(n1722_1),.b(n1725_1),.q(n1728));
  and_bi g775(.a(n774_0),.b(n726_0),.q(n775));
  spl2 g959_s_0(.a(n959),.q0(n959_0),.q1(n959_1));
  bfr _b_10433(.a(_w_12335),.q(_w_12336));
  and_bi g1530(.a(n1529_0),.b(n1452_0),.q(n1530));
  and_bi g1407(.a(n1406_0),.b(n1377_0),.q(n1407));
  bfr _b_5374(.a(_w_7276),.q(_w_7277));
  bfr _b_13344(.a(_w_15246),.q(_w_15247));
  bfr _b_8637(.a(_w_10539),.q(_w_10540));
  bfr _b_4845(.a(_w_6747),.q(_w_6748));
  and_bb g1023(.a(n1021_1),.b(n943_1),.q(_w_9132));
  and_bi g397(.a(n396_0),.b(n372_0),.q(n397));
  bfr _b_12317(.a(_w_14219),.q(_w_14220));
  bfr _b_11608(.a(_w_13510),.q(_w_13511));
  bfr _b_5596(.a(_w_7498),.q(N69_14));
  bfr _b_13062(.a(_w_14964),.q(_w_14965));
  and_bi g1258(.a(n1163_1),.b(n1256_1),.q(_w_9133));
  bfr _b_13761(.a(_w_15663),.q(_w_15664));
  or_bb g1303(.a(n1285_0),.b(n1302_0),.q(n1303));
  and_bi g1661(.a(n1659_0),.b(n1660),.q(n1661));
  and_bi g1263(.a(n1262_0),.b(n1161_0),.q(n1263));
  bfr _b_7877(.a(_w_9779),.q(_w_9780));
  or_bb g765(.a(n763_0),.b(n764),.q(n765));
  or_bb g1759(.a(n1733_0),.b(n1758_0),.q(n1759));
  and_bb g755(.a(n733_1),.b(n753_1),.q(_w_9137));
  bfr _b_3535(.a(_w_5437),.q(_w_5438));
  bfr _b_3447(.a(_w_5349),.q(_w_5350));
  bfr _b_4013(.a(_w_5915),.q(_w_5916));
  bfr _b_6089(.a(_w_7991),.q(_w_7992));
  bfr _b_5493(.a(_w_7395),.q(_w_7396));
  bfr _b_3883(.a(_w_5785),.q(_w_5786));
  spl2 g463_s_0(.a(n463),.q0(n463_0),.q1(n463_1));
  and_bi g752(.a(n734_1),.b(n750_1),.q(_w_9138));
  and_bi g475(.a(n474_0),.b(n450_0),.q(n475));
  and_bi g855(.a(n846_1),.b(n853_1),.q(_w_10572));
  bfr _b_3654(.a(_w_5556),.q(_w_5557));
  bfr _b_3632(.a(_w_5534),.q(_w_5535));
  and_bi g1355(.a(n1268_1),.b(n1353_1),.q(_w_13435));
  bfr _b_10211(.a(_w_12113),.q(_w_12114));
  or_bb g747(.a(n745_0),.b(n746),.q(n747));
  bfr _b_13703(.a(_w_15605),.q(_w_15606));
  bfr _b_6464(.a(_w_8366),.q(_w_8367));
  bfr _b_8692(.a(_w_10594),.q(n1414));
  and_bi g818(.a(n712_1),.b(n816_1),.q(_w_9139));
  bfr _b_3689(.a(_w_5591),.q(_w_5592));
  bfr _b_8733(.a(_w_10635),.q(_w_10636));
  and_bb g743(.a(n636_2),.b(n741_1),.q(_w_9140));
  spl2 g660_s_0(.a(n660),.q0(n660_0),.q1(n660_1));
  spl2 g521_s_0(.a(n521),.q0(n521_0),.q1(n521_1));
  bfr _b_13328(.a(_w_15230),.q(_w_15231));
  bfr _b_9895(.a(_w_11797),.q(_w_11798));
  or_bb g742(.a(n636_1),.b(n741_0),.q(n742));
  or_bb g1799(.a(n1797_0),.b(n1798),.q(n1799));
  bfr _b_13725(.a(_w_15627),.q(_w_15628));
  or_bb g740(.a(n635_1),.b(n739_0),.q(n740));
  bfr _b_5316(.a(_w_7218),.q(_w_7219));
  bfr _b_5947(.a(_w_7849),.q(_w_7850));
  bfr _b_10395(.a(_w_12297),.q(_w_12298));
  bfr _b_7970(.a(_w_9872),.q(_w_9873));
  bfr _b_8643(.a(_w_10545),.q(_w_10546));
  bfr _b_4165(.a(_w_6067),.q(_w_6068));
  and_bb g730(.a(N154_9),.b(N358_13),.q(_w_9177));
  bfr _b_9048(.a(_w_10950),.q(_w_10951));
  bfr _b_11429(.a(_w_13331),.q(_w_13332));
  bfr _b_11162(.a(_w_13064),.q(_w_13065));
  and_bi g933(.a(n820_1),.b(n931_1),.q(_w_9185));
  bfr _b_11523(.a(_w_13425),.q(n1337));
  bfr _b_4644(.a(_w_6546),.q(_w_6547));
  and_bb g726(.a(N120_11),.b(N392_11),.q(n726));
  bfr _b_12781(.a(_w_14683),.q(_w_14684));
  spl2 g1509_s_0(.a(n1509),.q0(n1509_0),.q1(_w_12820));
  bfr _b_6409(.a(_w_8311),.q(_w_8312));
  and_bb g712(.a(N1_18),.b(N511_4),.q(_w_9186));
  bfr _b_13992(.a(_w_15894),.q(_w_15895));
  and_bb g641(.a(n542_2),.b(n639_1),.q(_w_9202));
  bfr _b_7511(.a(_w_9413),.q(_w_9414));
  bfr _b_7628(.a(_w_9530),.q(_w_9531));
  and_bi g961(.a(n852_1),.b(n854_1),.q(n961));
  and_bi g725(.a(n670_1),.b(n673_1),.q(n725));
  and_bi g1109(.a(n1107_0),.b(n1108),.q(n1109));
  bfr _b_12331(.a(_w_14233),.q(n1827_1));
  or_bb g1575(.a(n1573_0),.b(n1574),.q(n1575));
  bfr _b_7219(.a(_w_9121),.q(_w_9122));
  and_bb g1795(.a(n1784_1),.b(n1793_1),.q(_w_14522));
  and_bb g720(.a(N443_8),.b(N69_14),.q(_w_9204));
  bfr _b_6940(.a(_w_8842),.q(_w_8843));
  bfr _b_13733(.a(_w_15635),.q(_w_15636));
  bfr _b_4707(.a(_w_6609),.q(_w_6610));
  bfr _b_8243(.a(_w_10145),.q(_w_10146));
  bfr _b_3699(.a(_w_5601),.q(_w_5602));
  spl2 g79_s_0(.a(n79),.q0(n79_0),.q1(n79_1));
  spl2 g1584_s_0(.a(n1584),.q0(n1584_0),.q1(n1584_1));
  bfr _b_4236(.a(_w_6138),.q(_w_6139));
  bfr _b_6179(.a(_w_8081),.q(_w_8082));
  bfr _b_3660(.a(_w_5562),.q(_w_5563));
  bfr _b_13570(.a(_w_15472),.q(_w_15473));
  and_bi g1007(.a(n1006_0),.b(n948_0),.q(n1007));
  and_bi g1706(.a(n1704_0),.b(n1705),.q(n1706));
  bfr _b_10340(.a(_w_12242),.q(_w_12243));
  bfr _b_7928(.a(_w_9830),.q(_w_9831));
  bfr _b_3933(.a(_w_5835),.q(_w_5836));
  and_bi g1401(.a(n1400_0),.b(n1379_0),.q(n1401));
  spl2 g365_s_0(.a(n365),.q0(n365_0),.q1(n365_1));
  bfr _b_13896(.a(_w_15798),.q(_w_15799));
  or_bb g268(.a(n239_0),.b(n267_0),.q(n268));
  or_bb g1686(.a(n1684_0),.b(n1685_0),.q(n1686));
  bfr _b_4865(.a(_w_6767),.q(_w_6768));
  spl2 g738_s_0(.a(n738),.q0(n738_0),.q1(_w_6185));
  and_bi g715(.a(n700_1),.b(n703_1),.q(n715));
  bfr _b_6754(.a(_w_8656),.q(_w_8657));
  bfr _b_7272(.a(_w_9174),.q(_w_9175));
  bfr _b_4854(.a(_w_6756),.q(_w_6757));
  and_bi g115(.a(n114_0),.b(n106_0),.q(n115));
  and_bb g106(.a(N307_7),.b(N52_6),.q(_w_9211));
  bfr _b_7126(.a(_w_9028),.q(_w_9029));
  bfr _b_11351(.a(_w_13253),.q(_w_13254));
  and_bi g1613(.a(n1576_1),.b(n1579_1),.q(n1613));
  bfr _b_6063(.a(_w_7965),.q(_w_7966));
  bfr _b_9190(.a(_w_11092),.q(_w_11093));
  and_bb g707(.a(n613_1),.b(n705_1),.q(_w_9217));
  bfr _b_13250(.a(_w_15152),.q(_w_15153));
  bfr _b_8389(.a(_w_10291),.q(_w_10292));
  or_bb g605(.a(n603_0),.b(n604),.q(n605));
  bfr _b_4771(.a(_w_6673),.q(_w_6674));
  spl2 g1000_s_0(.a(n1000),.q0(n1000_0),.q1(n1000_1));
  spl2 g1475_s_0(.a(n1475),.q0(n1475_0),.q1(n1475_1));
  bfr _b_13135(.a(_w_15037),.q(_w_15038));
  spl2 g452_s_0(.a(n452),.q0(n452_0),.q1(n452_1));
  bfr _b_14211(.a(_w_16113),.q(_w_16114));
  bfr _b_6630(.a(_w_8532),.q(_w_8533));
  and_bi g703(.a(n702_0),.b(n614_0),.q(n703));
  or_bb g1704(.a(n1678_0),.b(n1703_0),.q(n1704));
  bfr _b_5836(.a(_w_7738),.q(_w_7739));
  bfr _b_3634(.a(_w_5536),.q(_w_5537));
  bfr _b_13661(.a(_w_15563),.q(_w_15564));
  bfr _b_8275(.a(_w_10177),.q(_w_10178));
  bfr _b_9789(.a(_w_11691),.q(_w_11692));
  bfr _b_11664(.a(_w_13566),.q(_w_13567));
  spl2 g1168_s_0(.a(n1168),.q0(n1168_0),.q1(n1168_1));
  bfr _b_8356(.a(_w_10258),.q(_w_10259));
  spl2 g836_s_0(.a(n836),.q0(n836_0),.q1(n836_1));
  or_bb g700(.a(n615_0),.b(n699_0),.q(n700));
  bfr _b_3930(.a(_w_5832),.q(_w_5833));
  bfr _b_9871(.a(_w_11773),.q(_w_11774));
  spl2 g786_s_0(.a(n786),.q0(n786_0),.q1(n786_1));
  spl2 g1835_s_0(.a(n1835),.q0(n1835_0),.q1(n1835_1));
  and_bi g698(.a(n616_1),.b(n696_1),.q(_w_9218));
  and_bi g334(.a(n300_1),.b(n332_1),.q(_w_13096));
  and_bi g1671(.a(n1665_1),.b(n1668_1),.q(n1671));
  bfr _b_11713(.a(_w_13615),.q(_w_13616));
  spl4L N392_s_2(.a(N392_1),.q0(N392_8),.q1(N392_9),.q2(N392_10),.q3(N392_11));
  and_bb g647(.a(n633_1),.b(n645_1),.q(_w_9219));
  spl4L N1_s_0(.a(_w_15522),.q0(N1_0),.q1(_w_13584),.q2(_w_13606),.q3(_w_13660));
  bfr _b_4358(.a(_w_6260),.q(_w_6261));
  spl2 g939_s_0(.a(n939),.q0(n939_0),.q1(n939_1));
  spl2 g303_s_0(.a(n303),.q0(n303_0),.q1(n303_1));
  and_bi g1572(.a(n1570_0),.b(n1571),.q(n1572));
  bfr _b_9152(.a(_w_11054),.q(_w_11055));
  bfr _b_4392(.a(_w_6294),.q(_w_6295));
  and_bi g1808(.a(n1806_0),.b(n1807),.q(n1808));
  and_bb g689(.a(n619_1),.b(n687_1),.q(_w_9221));
  bfr _b_8261(.a(_w_10163),.q(_w_10164));
  bfr _b_4381(.a(_w_6283),.q(n286_1));
  bfr _b_4152(.a(_w_6054),.q(_w_6055));
  bfr _b_10225(.a(_w_12127),.q(_w_12128));
  bfr _b_3407(.a(_w_5309),.q(_w_5310));
  and_bb g309(.a(N154_5),.b(N273_13),.q(n309));
  spl2 g173_s_0(.a(n173),.q0(n173_0),.q1(n173_1));
  bfr _b_11451(.a(_w_13353),.q(_w_13354));
  and_bi g1305(.a(n1303_0),.b(n1304),.q(n1305));
  and_bb g534(.a(N120_9),.b(N358_11),.q(_w_12721));
  bfr _b_7447(.a(_w_9349),.q(_w_9350));
  spl2 g1472_s_0(.a(n1472),.q0(n1472_0),.q1(n1472_1));
  spl2 g880_s_0(.a(n880),.q0(n880_0),.q1(n880_1));
  and_bi g1866(.a(n1864_0),.b(n1865),.q(n1866));
  bfr _b_4789(.a(_w_6691),.q(_w_6692));
  bfr _b_13105(.a(_w_15007),.q(_w_15008));
  bfr _b_11195(.a(_w_13097),.q(_w_13098));
  spl2 g1825_s_0(.a(n1825),.q0(n1825_0),.q1(n1825_1));
  bfr _b_9962(.a(_w_11864),.q(_w_11865));
  and_bi g686(.a(n620_1),.b(n684_1),.q(_w_9226));
  bfr _b_10361(.a(_w_12263),.q(_w_12264));
  bfr _b_4045(.a(_w_5947),.q(_w_5948));
  bfr _b_9472(.a(_w_11374),.q(_w_11375));
  bfr _b_14026(.a(_w_15928),.q(_w_15929));
  bfr _b_3563(.a(_w_5465),.q(_w_5466));
  and_bi g1209(.a(n1208_0),.b(n1179_0),.q(n1209));
  bfr _b_13189(.a(_w_15091),.q(_w_15092));
  bfr _b_7603(.a(_w_9505),.q(_w_9506));
  bfr _b_4860(.a(_w_6762),.q(_w_6763));
  bfr _b_5750(.a(_w_7652),.q(_w_7653));
  spl2 g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1));
  or_bb g892(.a(n890_0),.b(n891),.q(n892));
  and_bb g180(.a(N1_11),.b(N392_4),.q(n180));
  spl2 g1069_s_0(.a(n1069),.q0(n1069_0),.q1(n1069_1));
  and_bi g1330(.a(n1329_0),.b(n1276_0),.q(n1330));
  bfr _b_7145(.a(_w_9047),.q(_w_9048));
  spl2 g1443_s_0(.a(n1443),.q0(n1443_0),.q1(n1443_1));
  bfr _b_13428(.a(_w_15330),.q(_w_15331));
  bfr _b_3549(.a(_w_5451),.q(_w_5452));
  bfr _b_6266(.a(_w_8168),.q(_w_8169));
  and_bi g141(.a(n118_1),.b(n121_1),.q(n141));
  or_bb g194(.a(n145_1),.b(n193_0),.q(_w_9244));
  bfr _b_5637(.a(_w_7539),.q(_w_7540));
  bfr _b_5708(.a(_w_7610),.q(_w_7611));
  bfr _b_3791(.a(_w_5693),.q(_w_5694));
  bfr _b_3486(.a(_w_5388),.q(_w_5389));
  bfr _b_7632(.a(_w_9534),.q(_w_9535));
  bfr _b_6395(.a(_w_8297),.q(_w_8298));
  and_bb g773(.a(n727_1),.b(n771_1),.q(_w_9245));
  and_bi g680(.a(n622_1),.b(n678_1),.q(_w_9246));
  bfr _b_4431(.a(_w_6333),.q(n1028_1));
  bfr _b_11050(.a(_w_12952),.q(_w_12953));
  spl2 g1356_s_0(.a(n1356),.q0(n1356_0),.q1(n1356_1));
  spl2 g935_s_0(.a(n935),.q0(n935_0),.q1(n935_1));
  and_bi g596(.a(n594_0),.b(n595),.q(n596));
  or_bb g1765(.a(n1731_0),.b(n1764_0),.q(n1765));
  or_bb g980(.a(n957_0),.b(n979_0),.q(n980));
  bfr _b_5185(.a(_w_7087),.q(_w_7088));
  and_bi g678(.a(n676_0),.b(n677),.q(n678));
  spl2 g719_s_0(.a(n719),.q0(n719_0),.q1(n719_1));
  bfr _b_4221(.a(_w_6123),.q(_w_6124));
  and_bi g53(.a(n46_1),.b(n49_1),.q(n53));
  and_bi g673(.a(n672_0),.b(n624_0),.q(n673));
  bfr _b_6280(.a(_w_8182),.q(_w_8183));
  bfr _b_6455(.a(_w_8357),.q(n227));
  bfr _b_10445(.a(_w_12347),.q(_w_12348));
  and_bb g1138(.a(n1055_1),.b(n1136_1),.q(_w_9249));
  and_bi g1627(.a(n1620_1),.b(n1625_1),.q(_w_9250));
  bfr _b_4926(.a(_w_6828),.q(_w_6829));
  bfr _b_8017(.a(_w_9919),.q(_w_9920));
  bfr _b_6390(.a(_w_8292),.q(_w_8293));
  and_bb g1654(.a(n1611_1),.b(n1652_1),.q(_w_9251));
  bfr _b_14309(.a(_w_16211),.q(_w_16212));
  bfr _b_9179(.a(_w_11081),.q(n154));
  bfr _b_10621(.a(_w_12523),.q(n518));
  and_bi g667(.a(n666_0),.b(n626_0),.q(n667));
  bfr _b_7513(.a(_w_9415),.q(_w_9416));
  bfr _b_3474(.a(_w_5376),.q(_w_5377));
  or_bb g1125(.a(n1059_0),.b(n1124_0),.q(n1125));
  spl2 g899_s_0(.a(n899),.q0(n899_0),.q1(_w_11832));
  and_bb g113(.a(n111_1),.b(n78_2),.q(_w_8807));
  spl2 g967_s_0(.a(n967),.q0(n967_0),.q1(n967_1));
  and_bi g666(.a(n664_0),.b(n665),.q(n666));
  bfr _b_6779(.a(_w_8681),.q(_w_8682));
  spl2 g1794_s_0(.a(n1794),.q0(n1794_0),.q1(_w_14952));
  or_bb g348(.a(n295_0),.b(n347_0),.q(n348));
  bfr _b_9428(.a(_w_11330),.q(_w_11331));
  bfr _b_7012(.a(_w_8914),.q(_w_8915));
  spl2 g342_s_0(.a(n342),.q0(n342_0),.q1(_w_15312));
  and_bi g1685(.a(n1623_1),.b(n1626_1),.q(n1685));
  bfr _b_13974(.a(_w_15876),.q(_w_15877));
  bfr _b_11264(.a(_w_13166),.q(_w_13167));
  or_bb g1136(.a(n1134_0),.b(n1135),.q(n1136));
  bfr _b_11677(.a(_w_13579),.q(n1840));
  and_bi g1894(.a(n1881_1),.b(n1884_1),.q(n1894));
  or_bb g606(.a(n521_0),.b(n605_0),.q(n606));
  bfr _b_13329(.a(_w_15231),.q(_w_15232));
  bfr _b_3460(.a(_w_5362),.q(_w_5363));
  and_bi g660(.a(n658_0),.b(n659),.q(n660));
  bfr _b_14094(.a(_w_15996),.q(_w_15997));
  bfr _b_4363(.a(_w_6265),.q(_w_6266));
  spl2 g55_s_0(.a(n55),.q0(n55_0),.q1(n55_1));
  bfr _b_4953(.a(_w_6855),.q(_w_6856));
  bfr _b_4672(.a(_w_6574),.q(_w_6575));
  or_bb g658(.a(n629_0),.b(n657_0),.q(n658));
  bfr _b_14267(.a(_w_16169),.q(_w_16170));
  spl2 g183_s_0(.a(n183),.q0(n183_0),.q1(n183_1));
  and_bi g835(.a(n772_1),.b(n775_1),.q(n835));
  bfr _b_11137(.a(_w_13039),.q(_w_13040));
  bfr _b_4577(.a(_w_6479),.q(_w_6480));
  and_bi g656(.a(n630_1),.b(n654_1),.q(_w_9261));
  or_bb g60(.a(n42_1),.b(n59_0),.q(n60));
  and_bi g1803(.a(n1802_0),.b(n1781_0),.q(n1803));
  and_bb g1616(.a(N205_15),.b(N460_16),.q(_w_9262));
  and_bi g723(.a(n676_1),.b(n679_1),.q(n723));
  bfr _b_5951(.a(_w_7853),.q(_w_7854));
  bfr _b_3524(.a(_w_5426),.q(_w_5427));
  spl2 g1434_s_0(.a(n1434),.q0(n1434_0),.q1(_w_9274));
  spl2 g1059_s_0(.a(n1059),.q0(n1059_0),.q1(n1059_1));
  or_bb g250(.a(n192_1),.b(n249_0),.q(n250));
  bfr _b_5516(.a(_w_7418),.q(_w_7419));
  bfr _b_5594(.a(_w_7496),.q(_w_7497));
  bfr _b_7556(.a(_w_9458),.q(_w_9459));
  bfr _b_13652(.a(_w_15554),.q(_w_15555));
  bfr _b_4333(.a(_w_6235),.q(_w_6236));
  spl2 g551_s_0(.a(n551),.q0(n551_0),.q1(n551_1));
  and_bi g650(.a(n632_1),.b(n648_1),.q(_w_9290));
  spl2 g207_s_0(.a(n207),.q0(n207_0),.q1(n207_1));
  and_bi g1055(.a(n1022_1),.b(n1025_1),.q(n1055));
  or_bb g645(.a(n643_0),.b(n644),.q(n645));
  bfr _b_3665(.a(_w_5567),.q(_w_5568));
  and_bb g559(.a(n537_1),.b(n557_1),.q(_w_9292));
  and_bb g1601(.a(n1534_1),.b(n1599_1),.q(_w_9293));
  bfr _b_4759(.a(_w_6661),.q(_w_6662));
  or_bb g1634(.a(n1632_0),.b(n1633),.q(n1634));
  bfr _b_5046(.a(_w_6948),.q(_w_6949));
  and_bi g859(.a(n857_0),.b(n858),.q(n859));
  bfr _b_7011(.a(_w_8913),.q(_w_8914));
  bfr _b_8370(.a(_w_10272),.q(_w_10273));
  bfr _b_11220(.a(_w_13122),.q(_w_13123));
  bfr _b_3916(.a(_w_5818),.q(_w_5819));
  bfr _b_5620(.a(_w_7522),.q(_w_7523));
  bfr _b_6104(.a(_w_8006),.q(_w_8007));
  and_bi g639(.a(n638),.b(n636_0),.q(n639));
  bfr _b_4046(.a(_w_5948),.q(_w_5949));
  bfr _b_5236(.a(_w_7138),.q(_w_7139));
  bfr _b_6489(.a(_w_8391),.q(_w_8392));
  bfr _b_10678(.a(_w_12580),.q(_w_12581));
  bfr _b_8450(.a(_w_10352),.q(_w_10353));
  and_bb g952(.a(N154_11),.b(N392_13),.q(n952));
  bfr _b_3455(.a(_w_5357),.q(_w_5358));
  bfr _b_8835(.a(_w_10737),.q(_w_10738));
  and_bb g637(.a(N222_21),.b(N273_17),.q(n637));
  and_bi g299(.a(n268_1),.b(n271_1),.q(n299));
  bfr _b_8385(.a(_w_10287),.q(_w_10288));
  bfr _b_4914(.a(_w_6816),.q(_w_6817));
  bfr _b_4812(.a(_w_6714),.q(_w_6715));
  bfr _b_9577(.a(_w_11479),.q(_w_11480));
  bfr _b_11452(.a(_w_13354),.q(_w_13355));
  and_bb g1820(.a(N205_19),.b(N528_16),.q(_w_9314));
  bfr _b_8631(.a(_w_10533),.q(_w_10534));
  and_bb g1056(.a(N477_9),.b(N86_16),.q(n1056));
  bfr _b_4614(.a(_w_6516),.q(_w_6517));
  bfr _b_5601(.a(_w_7503),.q(_w_7504));
  or_bb g1034(.a(n1033_0),.b(n939_0),.q(n1034));
  and_bb g1447(.a(n1364_1),.b(n1445_1),.q(_w_9338));
  bfr _b_14251(.a(_w_16153),.q(_w_16154));
  or_bb g1800(.a(n1782_0),.b(n1799_0),.q(n1800));
  spl4L N358_s_1(.a(N358_0),.q0(N358_4),.q1(N358_5),.q2(N358_6),.q3(N358_7));
  spl2 g952_s_0(.a(n952),.q0(n952_0),.q1(n952_1));
  bfr _b_7452(.a(_w_9354),.q(_w_9355));
  bfr _b_6497(.a(_w_8399),.q(_w_8400));
  bfr _b_3694(.a(_w_5596),.q(_w_5597));
  and_bi g629(.a(n558_1),.b(n561_1),.q(n629));
  and_bi g1312(.a(n1311_0),.b(n1282_0),.q(n1312));
  bfr _b_8558(.a(_w_10460),.q(_w_10461));
  spl2 g1623_s_0(.a(n1623),.q0(n1623_0),.q1(_w_9339));
  and_bi g1208(.a(n1206_0),.b(n1207),.q(n1208));
  and_bi g805(.a(n804_0),.b(n716_0),.q(n805));
  spl2 g1239_s_0(.a(n1239),.q0(n1239_0),.q1(n1239_1));
  bfr _b_4479(.a(_w_6381),.q(n42_2));
  bfr _b_6567(.a(_w_8469),.q(_w_8470));
  bfr _b_10622(.a(_w_12524),.q(_w_12525));
  bfr _b_8199(.a(_w_10101),.q(_w_10102));
  spl2 g323_s_0(.a(n323),.q0(n323_0),.q1(n323_1));
  spl3L g636_s_0(.a(n636),.q0(n636_0),.q1(_w_9343),.q2(_w_9345));
  bfr _b_6514(.a(_w_8416),.q(_w_8417));
  bfr _b_13888(.a(_w_15790),.q(_w_15791));
  bfr _b_7101(.a(_w_9003),.q(_w_9004));
  and_bi g895(.a(n893_0),.b(n894),.q(n895));
  spl2 g1564_s_0(.a(n1564),.q0(n1564_0),.q1(_w_9364));
  or_bb g1253(.a(n1251_0),.b(n1252),.q(n1253));
  spl2 g1323_s_0(.a(n1323),.q0(n1323_0),.q1(n1323_1));
  spl2 g1526_s_0(.a(n1526),.q0(n1526_0),.q1(n1526_1));
  and_bi g621(.a(n582_1),.b(n585_1),.q(n621));
  bfr _b_13670(.a(_w_15572),.q(_w_15573));
  and_bi g746(.a(n736_1),.b(n744_1),.q(_w_9372));
  spl2 g1679_s_0(.a(n1679),.q0(n1679_0),.q1(n1679_1));
  and_bi g939(.a(n917_1),.b(n920_1),.q(n939));
  bfr _b_11839(.a(_w_13741),.q(_w_13742));
  and_bb g1075(.a(N256_18),.b(N307_19),.q(_w_9541));
  and_bb g767(.a(n729_1),.b(n765_1),.q(_w_9548));
  bfr _b_5760(.a(_w_7662),.q(_w_7663));
  bfr _b_8494(.a(_w_10396),.q(_w_10397));
  bfr _b_4556(.a(_w_6458),.q(_w_6459));
  bfr _b_9399(.a(_w_11301),.q(_w_11302));
  bfr _b_10219(.a(_w_12121),.q(_w_12122));
  bfr _b_10631(.a(_w_12533),.q(_w_12534));
  spl2 g202_s_0(.a(n202),.q0(n202_0),.q1(_w_6284));
  or_bb g1027(.a(n1025_0),.b(n1026),.q(n1027));
  and_bb g616(.a(N35_15),.b(N460_6),.q(_w_9549));
  spl4L N375_s_4(.a(N375_3),.q0(N375_16),.q1(N375_17),.q2(N375_18),.q3(N375_19));
  bfr _b_9529(.a(_w_11431),.q(_w_11432));
  and_bi g615(.a(n600_1),.b(n603_1),.q(n615));
  bfr _b_8549(.a(_w_10451),.q(n785));
  and_bi g1105(.a(n1066_1),.b(n1103_1),.q(_w_9561));
  spl2 g1220_s_0(.a(n1220),.q0(n1220_0),.q1(n1220_1));
  spl2 g1611_s_0(.a(n1611),.q0(n1611_0),.q1(n1611_1));
  or_bb g813(.a(n811_0),.b(n812),.q(n813));
  bfr _b_14230(.a(_w_16132),.q(_w_16133));
  or_bb g507(.a(n505_0),.b(n506),.q(n507));
  and_bb g614(.a(N18_16),.b(N477_5),.q(n614));
  and_bb g1334(.a(n1275_1),.b(n1332_1),.q(_w_10780));
  bfr _b_11016(.a(_w_12918),.q(_w_12919));
  bfr _b_6334(.a(_w_8236),.q(_w_8237));
  bfr _b_3896(.a(_w_5798),.q(_w_5799));
  bfr _b_6874(.a(_w_8776),.q(n867));
  bfr _b_12329(.a(_w_14231),.q(_w_14232));
  bfr _b_7277(.a(_w_9179),.q(_w_9180));
  spl2 g578_s_0(.a(n578),.q0(n578_0),.q1(n578_1));
  and_bi g39(.a(n38),.b(n35_0),.q(_w_11406));
  spl2 g936_s_0(.a(n936),.q0(n936_0),.q1(n936_1));
  bfr _b_5860(.a(_w_7762),.q(_w_7763));
  and_bi g608(.a(n606_0),.b(n607),.q(n608));
  bfr _b_4288(.a(_w_6190),.q(_w_6191));
  and_bi g757(.a(n756_0),.b(n732_0),.q(n757));
  bfr _b_4780(.a(_w_6682),.q(_w_6683));
  and_bi g160(.a(n142_1),.b(n158_1),.q(_w_9567));
  bfr _b_8303(.a(_w_10205),.q(n1641_1));
  spl2 g940_s_0(.a(n940),.q0(n940_0),.q1(n940_1));
  bfr _b_6320(.a(_w_8222),.q(_w_8223));
  spl2 g1413_s_0(.a(n1413),.q0(n1413_0),.q1(n1413_1));
  bfr _b_10012(.a(_w_11914),.q(_w_11915));
  bfr _b_4027(.a(_w_5929),.q(_w_5930));
  bfr _b_3758(.a(_w_5660),.q(_w_5661));
  bfr _b_14056(.a(_w_15958),.q(_w_15959));
  bfr _b_9360(.a(_w_11262),.q(_w_11263));
  spl2 g1575_s_0(.a(n1575),.q0(n1575_0),.q1(n1575_1));
  bfr _b_10245(.a(_w_12147),.q(_w_12148));
  spl2 g1858_s_0(.a(n1858),.q0(n1858_0),.q1(_w_9574));
  bfr _b_4925(.a(_w_6827),.q(_w_6828));
  bfr _b_3861(.a(_w_5763),.q(_w_5764));
  bfr _b_5690(.a(_w_7592),.q(_w_7593));
  or_bb g599(.a(n597_0),.b(n598),.q(n599));
  bfr _b_13109(.a(_w_15011),.q(_w_15012));
  and_bb g1185(.a(N239_8),.b(N341_18),.q(n1185));
  and_bi g254(.a(n244_1),.b(n252_1),.q(_w_10954));
  or_bb g1112(.a(n1110_0),.b(n1111),.q(n1112));
  or_bb g310(.a(n245_1),.b(n309_0),.q(_w_9583));
  spl2 g1790_s_0(.a(n1790),.q0(n1790_0),.q1(n1790_1));
  bfr _b_4489(.a(_w_6391),.q(_w_6392));
  spl2 g962_s_0(.a(n962),.q0(n962_0),.q1(_w_9584));
  bfr _b_12366(.a(_w_14268),.q(_w_14269));
  and_bi g1059(.a(n1010_1),.b(n1013_1),.q(n1059));
  and_bb g383(.a(n308_2),.b(n381_1),.q(_w_9588));
  and_bi g597(.a(n596_0),.b(n524_0),.q(n597));
  or_bb g754(.a(n733_0),.b(n753_0),.q(n754));
  bfr _b_7612(.a(_w_9514),.q(_w_9515));
  spl4L N239_s_3(.a(N239_2),.q0(N239_12),.q1(_w_5853),.q2(_w_5861),.q3(_w_5873));
  spl2 g296_s_0(.a(n296),.q0(n296_0),.q1(n296_1));
  and_bi g1042(.a(n1040_0),.b(n1041),.q(n1042));
  bfr _b_8551(.a(_w_10453),.q(_w_10454));
  bfr _b_3442(.a(_w_5344),.q(_w_5345));
  or_bb g1605(.a(n1603_0),.b(n1604),.q(_w_9589));
  or_bb g664(.a(n627_0),.b(n663_0),.q(n664));
  bfr _b_7455(.a(_w_9357),.q(_w_9358));
  or_bb g593(.a(n591_0),.b(n592),.q(n593));
  bfr _b_11495(.a(_w_13397),.q(_w_13398));
  bfr _b_6757(.a(_w_8659),.q(_w_8660));
  bfr _b_7736(.a(_w_9638),.q(n674));
  bfr _b_8063(.a(_w_9965),.q(_w_9966));
  bfr _b_4866(.a(_w_6768),.q(_w_6769));
  or_bb g1422(.a(n1372_0),.b(n1421_0),.q(n1422));
  bfr _b_5787(.a(_w_7689),.q(_w_7690));
  and_bi g831(.a(n784_1),.b(n787_1),.q(n831));
  bfr _b_6208(.a(_w_8110),.q(_w_8111));
  and_bi g63(.a(n62_0),.b(n54_0),.q(n63));
  bfr _b_9628(.a(_w_11530),.q(_w_11531));
  bfr _b_13530(.a(_w_15432),.q(_w_15433));
  bfr _b_10195(.a(_w_12097),.q(n1687));
  bfr _b_3456(.a(_w_5358),.q(_w_5359));
  and_bi g976(.a(n974_0),.b(n975),.q(n976));
  bfr _b_7737(.a(_w_9639),.q(n583));
  and_bb g294(.a(N18_12),.b(N409_5),.q(n294));
  bfr _b_5320(.a(_w_7222),.q(_w_7223));
  bfr _b_12412(.a(_w_14314),.q(_w_14315));
  bfr _b_4594(.a(_w_6496),.q(_w_6497));
  bfr _b_3707(.a(_w_5609),.q(_w_5610));
  bfr _b_8533(.a(_w_10435),.q(_w_10436));
  bfr _b_6134(.a(_w_8036),.q(_w_8037));
  and_bb g930(.a(n821_1),.b(n928_1),.q(_w_8725));
  and_bb g894(.a(n833_1),.b(n892_1),.q(_w_9621));
  bfr _b_12786(.a(_w_14688),.q(n1874));
  and_bi g592(.a(n526_1),.b(n590_1),.q(_w_9622));
  bfr _b_4661(.a(_w_6563),.q(_w_6564));
  bfr _b_10089(.a(_w_11991),.q(_w_11992));
  bfr _b_4449(.a(_w_6351),.q(_w_6352));
  bfr _b_4939(.a(_w_6841),.q(_w_6842));
  and_bi g591(.a(n590_0),.b(n526_0),.q(n591));
  and_bb g1460(.a(N154_16),.b(N477_13),.q(n1460));
  bfr _b_4777(.a(_w_6679),.q(_w_6680));
  and_bb g300(.a(N358_8),.b(N69_9),.q(_w_9629));
  bfr _b_4719(.a(_w_6621),.q(_w_6622));
  bfr _b_12796(.a(_w_14698),.q(_w_14699));
  and_bb g589(.a(n527_1),.b(n587_1),.q(_w_9637));
  bfr _b_8599(.a(_w_10501),.q(_w_10502));
  and_bi g823(.a(n808_1),.b(n811_1),.q(n823));
  and_bb g815(.a(n713_1),.b(n813_1),.q(_w_9883));
  bfr _b_5972(.a(_w_7874),.q(N222_2));
  bfr _b_9990(.a(_w_11892),.q(_w_11893));
  and_bi g756(.a(n754_0),.b(n755),.q(n756));
  and_bi g1702(.a(n1679_1),.b(n1700_1),.q(_w_14116));
  bfr _b_5732(.a(_w_7634),.q(_w_7635));
  bfr _b_3490(.a(_w_5392),.q(_w_5393));
  spl2 g1100_s_0(.a(n1100),.q0(n1100_0),.q1(n1100_1));
  bfr _b_10060(.a(_w_11962),.q(_w_11963));
  bfr _b_5147(.a(_w_7049),.q(_w_7050));
  spl2 g1278_s_0(.a(n1278),.q0(n1278_0),.q1(n1278_1));
  bfr _b_13868(.a(_w_15770),.q(_w_15771));
  bfr _b_12123(.a(_w_14025),.q(_w_14026));
  bfr _b_10174(.a(_w_12076),.q(n1316));
  bfr _b_10345(.a(_w_12247),.q(_w_12248));
  and_bb g227(.a(n181_1),.b(n225_1),.q(_w_8357));
  spl2 g492_s_0(.a(n492),.q0(n492_0),.q1(n492_1));
  and_bi g1394(.a(n1392_0),.b(n1393),.q(n1394));
  bfr _b_4999(.a(_w_6901),.q(_w_6902));
  bfr _b_12111(.a(_w_14013),.q(_w_14014));
  spl2 g1703_s_0(.a(n1703),.q0(n1703_0),.q1(n1703_1));
  bfr _b_8799(.a(_w_10701),.q(_w_10702));
  bfr _b_3696(.a(_w_5598),.q(_w_5599));
  or_bb g80(.a(n55_1),.b(n79_0),.q(_w_13198));
  or_bb g581(.a(n579_0),.b(n580),.q(n581));
  and_bi g1001(.a(n1000_0),.b(n950_0),.q(n1001));
  bfr _b_14197(.a(_w_16099),.q(_w_16100));
  bfr _b_9601(.a(_w_11503),.q(_w_11504));
  and_bi g793(.a(n792_0),.b(n720_0),.q(n793));
  spl2 g896_s_0(.a(n896),.q0(n896_0),.q1(n896_1));
  bfr _b_5854(.a(_w_7756),.q(_w_7757));
  bfr _b_3457(.a(_w_5359),.q(_w_5360));
  spl2 g141_s_0(.a(n141),.q0(n141_0),.q1(n141_1));
  bfr _b_13201(.a(_w_15103),.q(_w_15104));
  or_bb g1593(.a(n1591_0),.b(n1592),.q(n1593));
  and_bb g1298(.a(n1287_1),.b(n1296_1),.q(_w_9640));
  and_bi g69(.a(n68_0),.b(n52_0),.q(n69));
  bfr _b_12394(.a(_w_14296),.q(_w_14297));
  bfr _b_10712(.a(_w_12614),.q(_w_12615));
  bfr _b_4170(.a(_w_6072),.q(_w_6073));
  bfr _b_8770(.a(_w_10672),.q(_w_10673));
  bfr _b_4840(.a(_w_6742),.q(_w_6743));
  bfr _b_5897(.a(_w_7799),.q(_w_7800));
  and_bb g632(.a(N171_7),.b(N324_14),.q(_w_9641));
  bfr _b_8652(.a(_w_10554),.q(_w_10555));
  and_bi g276(.a(n274_0),.b(n275),.q(n276));
  bfr _b_14268(.a(_w_16170),.q(_w_16171));
  bfr _b_6652(.a(_w_8554),.q(_w_8555));
  bfr _b_3427(.a(_w_5329),.q(_w_5330));
  spl2 g381_s_0(.a(n381),.q0(n381_0),.q1(n381_1));
  bfr _b_5687(.a(_w_7589),.q(_w_7590));
  bfr _b_7521(.a(_w_9423),.q(_w_9424));
  bfr _b_8449(.a(_w_10351),.q(_w_10352));
  and_bb g275(.a(n237_1),.b(n273_1),.q(_w_9659));
  bfr _b_10311(.a(_w_12213),.q(_w_12214));
  bfr _b_3990(.a(_w_5892),.q(_w_5893));
  spl2 g799_s_0(.a(n799),.q0(n799_0),.q1(n799_1));
  bfr _b_6931(.a(_w_8833),.q(_w_8834));
  and_bi g989(.a(n988_0),.b(n954_0),.q(n989));
  bfr _b_8756(.a(_w_10658),.q(_w_10659));
  and_bi g1250(.a(n1248_0),.b(n1249),.q(n1250));
  bfr _b_6177(.a(_w_8079),.q(_w_8080));
  bfr _b_7916(.a(_w_9818),.q(_w_9819));
  bfr _b_3844(.a(_w_5746),.q(_w_5747));
  bfr _b_9341(.a(_w_11243),.q(_w_11244));
  and_bb g526(.a(N426_7),.b(N52_13),.q(n526));
  bfr _b_12490(.a(_w_14392),.q(_w_14393));
  spl2 g298_s_0(.a(n298),.q0(n298_0),.q1(n298_1));
  bfr _b_9078(.a(_w_10980),.q(n749));
  bfr _b_11660(.a(_w_13562),.q(_w_13563));
  and_bi g1862(.a(n1855_1),.b(n1860_1),.q(_w_9684));
  bfr _b_4864(.a(_w_6766),.q(_w_6767));
  bfr _b_4694(.a(_w_6596),.q(_w_6597));
  spl2 g1082_s_0(.a(n1082),.q0(n1082_0),.q1(n1082_1));
  bfr _b_6198(.a(_w_8100),.q(_w_8101));
  or_bb g267(.a(n265_0),.b(n266),.q(n267));
  bfr _b_6612(.a(_w_8514),.q(_w_8515));
  bfr _b_8188(.a(_w_10090),.q(_w_10091));
  or_bb g546(.a(n456_1),.b(n545_0),.q(n546));
  and_bb g583(.a(n529_1),.b(n581_1),.q(_w_9639));
  and_bb g34(.a(N1_4),.b(N273_4),.q(N545_0));
  spl2 g409_s_0(.a(n409),.q0(n409_0),.q1(n409_1));
  bfr _b_8258(.a(_w_10160),.q(_w_10161));
  bfr _b_9463(.a(_w_11365),.q(_w_11366));
  bfr _b_4573(.a(_w_6475),.q(_w_6476));
  bfr _b_5054(.a(_w_6956),.q(_w_6957));
  bfr _b_4500(.a(_w_6402),.q(_w_6403));
  spl2 g910_s_0(.a(n910),.q0(n910_0),.q1(n910_1));
  bfr _b_6572(.a(_w_8474),.q(_w_8475));
  bfr _b_5193(.a(_w_7095),.q(_w_7096));
  bfr _b_5600(.a(_w_7502),.q(_w_7503));
  and_bi g282(.a(n280_0),.b(n281),.q(n282));
  spl2 g1311_s_0(.a(n1311),.q0(n1311_0),.q1(n1311_1));
  and_bi g1778(.a(n1765_1),.b(n1768_1),.q(n1778));
  bfr _b_14220(.a(_w_16122),.q(_w_16123));
  bfr _b_10328(.a(_w_12230),.q(_w_12231));
  and_bi g1655(.a(n1653_0),.b(n1654),.q(n1655));
  and_bi g97(.a(n96_0),.b(n72_0),.q(n97));
  bfr _b_4249(.a(_w_6151),.q(_w_6152));
  or_bb g262(.a(n241_0),.b(n261_0),.q(n262));
  bfr _b_5748(.a(_w_7650),.q(_w_7651));
  bfr _b_7861(.a(_w_9763),.q(_w_9764));
  and_bi g120(.a(n118_0),.b(n119),.q(n120));
  bfr _b_4422(.a(_w_6324),.q(n108_2));
  and_bi g654(.a(n652_0),.b(n653),.q(n654));
  bfr _b_10995(.a(_w_12897),.q(_w_12898));
  spl2 g158_s_0(.a(n158),.q0(n158_0),.q1(n158_1));
  bfr _b_6465(.a(_w_8367),.q(n1552_1));
  bfr _b_6912(.a(_w_8814),.q(_w_8815));
  bfr _b_11902(.a(_w_13804),.q(_w_13805));
  bfr _b_8476(.a(_w_10378),.q(_w_10379));
  and_bi g713(.a(n706_1),.b(n709_1),.q(n713));
  and_bb g724(.a(N103_12),.b(N409_10),.q(n724));
  bfr _b_12772(.a(_w_14674),.q(_w_14675));
  bfr _b_5887(.a(_w_7789),.q(_w_7790));
  and_bi g1578(.a(n1576_0),.b(n1577),.q(n1578));
  spl2 g1045_s_0(.a(n1045),.q0(n1045_0),.q1(n1045_1));
  bfr _b_4663(.a(_w_6565),.q(_w_6566));
  bfr _b_5930(.a(_w_7832),.q(_w_7833));
  bfr _b_6426(.a(_w_8328),.q(_w_8329));
  bfr _b_9756(.a(_w_11658),.q(_w_11659));
  and_bi g1546(.a(n1485_1),.b(n1488_1),.q(n1546));
  and_bi g827(.a(n796_1),.b(n799_1),.q(n827));
  bfr _b_11781(.a(_w_13683),.q(_w_13684));
  bfr _b_10422(.a(_w_12324),.q(_w_12325));
  and_bb g1813(.a(n1778_1),.b(n1811_1),.q(_w_9701));
  and_bi g1006(.a(n1004_0),.b(n1005),.q(n1006));
  bfr _b_6264(.a(_w_8166),.q(_w_8167));
  bfr _b_7059(.a(_w_8961),.q(_w_8962));
  bfr _b_4776(.a(_w_6678),.q(_w_6679));
  bfr _b_6533(.a(_w_8435),.q(_w_8436));
  spl2 g1286_s_0(.a(n1286),.q0(n1286_0),.q1(n1286_1));
  and_bi g369(.a(n330_1),.b(n333_1),.q(n369));
  and_bb g530(.a(N392_9),.b(N86_11),.q(n530));
  and_bi g1531(.a(n1452_1),.b(n1529_1),.q(_w_9738));
  spl2 g1847_s_0(.a(n1847),.q0(n1847_0),.q1(n1847_1));
  and_bb g454(.a(N154_6),.b(N307_13),.q(_w_9753));
  bfr _b_5559(.a(_w_7461),.q(_w_7462));
  bfr _b_7412(.a(_w_9314),.q(_w_9315));
  bfr _b_10530(.a(_w_12432),.q(_w_12433));
  or_bb g551(.a(n549_0),.b(n550),.q(n551));
  spl2 g396_s_0(.a(n396),.q0(n396_0),.q1(n396_1));
  and_bi g1792(.a(n1785_1),.b(n1790_1),.q(_w_14369));
  and_bi g631(.a(n552_1),.b(n555_1),.q(n631));
  and_bb g542(.a(n457_1),.b(n541_0),.q(n542));
  bfr _b_11988(.a(_w_13890),.q(_w_13891));
  or_bb g1247(.a(n1245_0),.b(n1246),.q(n1247));
  spl4L N443_s_1(.a(N443_0),.q0(N443_4),.q1(N443_5),.q2(N443_6),.q3(N443_7));
  or_bb g748(.a(n735_0),.b(n747_0),.q(n748));
  spl2 g750_s_0(.a(n750),.q0(n750_0),.q1(n750_1));
  bfr _b_12226(.a(_w_14128),.q(_w_14129));
  and_bb g1411(.a(n1376_1),.b(n1409_1),.q(_w_14824));
  bfr _b_4293(.a(_w_6195),.q(n694_1));
  bfr _b_12712(.a(_w_14614),.q(_w_14615));
  and_bi g449(.a(n394_1),.b(n397_1),.q(n449));
  spl2 g1671_s_0(.a(n1671),.q0(n1671_0),.q1(n1671_1));
  or_bb g513(.a(n511_0),.b(n512),.q(n513));
  or_bb g1118(.a(n1116_0),.b(n1117),.q(n1118));
  bfr _b_7158(.a(_w_9060),.q(_w_9061));
  and_bb g1666(.a(n1607_1),.b(n1664_1),.q(_w_9916));
  spl4L N290_s_1(.a(N290_0),.q0(N290_4),.q1(_w_9941),.q2(N290_6),.q3(N290_7));
  or_bb g694(.a(n617_0),.b(n693_0),.q(n694));
  bfr _b_6763(.a(_w_8665),.q(_w_8666));
  and_bb g192(.a(n147_1),.b(n191_0),.q(n192));
  bfr _b_9670(.a(_w_11572),.q(_w_11573));
  and_bb g1595(.a(n1536_1),.b(n1593_1),.q(_w_13956));
  bfr _b_4069(.a(_w_5971),.q(_w_5972));
  and_bi g619(.a(n588_1),.b(n591_1),.q(n619));
  spl2 g871_s_0(.a(n871),.q0(n871_0),.q1(n871_1));
  and_bi g277(.a(n276_0),.b(n236_0),.q(n277));
  spl2 g1469_s_0(.a(n1469),.q0(n1469_0),.q1(n1469_1));
  bfr _b_5182(.a(_w_7084),.q(_w_7085));
  bfr _b_9123(.a(_w_11025),.q(n86));
  bfr _b_4338(.a(_w_6240),.q(_w_6241));
  and_bi g1638(.a(n1637_0),.b(n1616_0),.q(n1638));
  bfr _b_7852(.a(_w_9754),.q(_w_9755));
  spl2 g721_s_0(.a(n721),.q0(n721_0),.q1(n721_1));
  bfr _b_6732(.a(_w_8634),.q(_w_8635));
  and_bi g229(.a(n228_0),.b(n180_0),.q(n229));
  bfr _b_5202(.a(_w_7104),.q(_w_7105));
  and_bi g101(.a(n94_1),.b(n97_1),.q(n101));
  bfr _b_7620(.a(_w_9522),.q(_w_9523));
  and_bb g1871(.a(n1852_1),.b(n1869_1),.q(_w_9947));
  spl2 g504_s_0(.a(n504),.q0(n504_0),.q1(n504_1));
  and_bb g221(.a(n183_1),.b(n219_1),.q(_w_9948));
  bfr _b_10458(.a(_w_12360),.q(_w_12361));
  bfr _b_8130(.a(_w_10032),.q(_w_10033));
  and_bi g116(.a(n106_1),.b(n114_1),.q(_w_9950));
  bfr _b_5612(.a(_w_7514),.q(_w_7515));
  and_bb g1474(.a(n1471_1),.b(n1472_1),.q(_w_9951));
  bfr _b_8797(.a(_w_10699),.q(_w_10700));
  spl2 g1119_s_0(.a(n1119),.q0(n1119_0),.q1(_w_9952));
  and_bi g1256(.a(n1254_0),.b(n1255),.q(n1256));
  bfr _b_7958(.a(_w_9860),.q(_w_9861));
  or_bb g1003(.a(n1001_0),.b(n1002),.q(n1003));
  bfr _b_3998(.a(_w_5900),.q(_w_5901));
  bfr _b_8535(.a(_w_10437),.q(_w_10438));
  and_bi g384(.a(n382_0),.b(n383),.q(n384));
  spl2 g572_s_0(.a(n572),.q0(n572_0),.q1(n572_1));
  bfr _b_4930(.a(_w_6832),.q(_w_6833));
  or_bb g1131(.a(n1057_0),.b(n1130_0),.q(n1131));
  bfr _b_7536(.a(_w_9438),.q(_w_9439));
  bfr _b_3440(.a(_w_5342),.q(_w_5343));
  bfr _b_13949(.a(_w_15851),.q(_w_15852));
  bfr _b_11458(.a(_w_13360),.q(_w_13361));
  spl2 g121_s_0(.a(n121),.q0(n121_0),.q1(n121_1));
  bfr _b_11653(.a(_w_13555),.q(_w_13556));
  and_bi g1349(.a(n1270_1),.b(n1347_1),.q(_w_9957));
  bfr _b_5922(.a(_w_7824),.q(_w_7825));
  and_bb g67(.a(n53_1),.b(n65_1),.q(_w_9958));
  bfr _b_14216(.a(_w_16118),.q(_w_16119));
  bfr _b_10522(.a(_w_12424),.q(n1405));
  bfr _b_6259(.a(_w_8161),.q(_w_8162));
  and_bb g1035(.a(n1033_1),.b(n939_1),.q(_w_11600));
  spl2 g869_s_0(.a(n869),.q0(n869_0),.q1(_w_9961));
  bfr _b_8517(.a(_w_10419),.q(_w_10420));
  bfr _b_4583(.a(_w_6485),.q(_w_6486));
  bfr _b_5923(.a(_w_7825),.q(_w_7826));
  spl2 g1780_s_0(.a(n1780),.q0(n1780_0),.q1(n1780_1));
  bfr _b_4065(.a(_w_5967),.q(_w_5968));
  and_bb g77(.a(N290_8),.b(N69_4),.q(n77));
  bfr _b_10946(.a(_w_12848),.q(n714));
  bfr _b_7435(.a(_w_9337),.q(n1820));
  bfr _b_9949(.a(_w_11851),.q(_w_11852));
  bfr _b_12296(.a(_w_14198),.q(_w_14199));
  and_bb g1379(.a(N205_12),.b(N409_16),.q(n1379));
  and_bi g159(.a(n158_0),.b(n142_0),.q(n159));
  bfr _b_7573(.a(_w_9475),.q(_w_9476));
  bfr _b_9451(.a(_w_11353),.q(_w_11354));
  and_bi g978(.a(n958_1),.b(n976_1),.q(_w_12301));
  bfr _b_14145(.a(_w_16047),.q(_w_16048));
  bfr _b_11877(.a(_w_13779),.q(_w_13780));
  bfr _b_6004(.a(_w_7906),.q(_w_7907));
  and_bi g210(.a(n208_0),.b(n209),.q(n210));
  bfr _b_11753(.a(_w_13655),.q(_w_13656));
  bfr _b_5014(.a(_w_6916),.q(_w_6917));
  bfr _b_11565(.a(_w_13467),.q(_w_13468));
  bfr _b_3925(.a(_w_5827),.q(_w_5828));
  bfr _b_6094(.a(_w_7996),.q(_w_7997));
  bfr _b_5036(.a(_w_6938),.q(_w_6939));
  and_bb g595(.a(n525_1),.b(n593_1),.q(_w_9973));
  and_bb g74(.a(N18_7),.b(N324_5),.q(_w_9974));
  bfr _b_9287(.a(_w_11189),.q(_w_11190));
  bfr _b_3889(.a(_w_5791),.q(_w_5792));
  or_bb g1028(.a(n1027_0),.b(n941_0),.q(n1028));
  bfr _b_12846(.a(_w_14748),.q(_w_14749));
  or_bb g1514(.a(n1512_0),.b(n1513),.q(n1514));
  bfr _b_10844(.a(_w_12746),.q(_w_12747));
  bfr _b_7934(.a(_w_9836),.q(_w_9837));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(_w_9988));
  and_bi g206(.a(n188_1),.b(n204_1),.q(_w_9992));
  bfr _b_3854(.a(_w_5756),.q(_w_5757));
  bfr _b_9574(.a(_w_11476),.q(_w_11477));
  bfr _b_4892(.a(_w_6794),.q(_w_6795));
  or_bb g71(.a(n69_0),.b(n70),.q(_w_9993));
  or_bb g1864(.a(n1854_0),.b(n1863_0),.q(n1864));
  bfr _b_12800(.a(_w_14702),.q(_w_14703));
  bfr _b_3493(.a(_w_5395),.q(_w_5396));
  bfr _b_4341(.a(_w_6243),.q(N120_15));
  and_bi g655(.a(n654_0),.b(n630_0),.q(n655));
  bfr _b_8605(.a(_w_10507),.q(_w_10508));
  and_bi g390(.a(n388_0),.b(n389),.q(n390));
  and_bi g1061(.a(n1004_1),.b(n1007_1),.q(n1061));
  bfr _b_8795(.a(_w_10697),.q(_w_10698));
  bfr _b_10935(.a(_w_12837),.q(_w_12838));
  or_bb g705(.a(n703_0),.b(n704),.q(n705));
  and_bb g987(.a(n955_1),.b(n985_1),.q(_w_10181));
  bfr _b_9838(.a(_w_11740),.q(_w_11741));
  and_bi g48(.a(n46_0),.b(n47),.q(n48));
  and_bi g172(.a(n138_1),.b(n170_1),.q(_w_10182));
  spl2 g223_s_0(.a(n223),.q0(n223_0),.q1(n223_1));
  bfr _b_10379(.a(_w_12281),.q(_w_12282));
  bfr _b_9223(.a(_w_11125),.q(_w_11126));
  or_bb g226(.a(n181_0),.b(n225_0),.q(n226));
  and_bi g506(.a(n440_1),.b(n504_1),.q(_w_11814));
  bfr _b_9690(.a(_w_11592),.q(N6260));
  spl2 g1404_s_0(.a(n1404),.q0(n1404_0),.q1(_w_10184));
  bfr _b_5819(.a(_w_7721),.q(_w_7722));
  bfr _b_4755(.a(_w_6657),.q(_w_6658));
  and_bb g1384(.a(N256_15),.b(N358_19),.q(_w_10188));
  bfr _b_12925(.a(_w_14827),.q(_w_14828));
  and_bb g888(.a(n835_1),.b(n886_1),.q(_w_10200));
  or_bb g1869(.a(n1867_0),.b(n1868),.q(_w_8229));
  and_bi g925(.a(n923_0),.b(n924),.q(n925));
  bfr _b_7044(.a(_w_8946),.q(_w_8947));
  bfr _b_7218(.a(_w_9120),.q(_w_9121));
  and_bi g690(.a(n688_0),.b(n689),.q(n690));
  bfr _b_8616(.a(_w_10518),.q(_w_10519));
  bfr _b_4124(.a(_w_6026),.q(_w_6027));
  bfr _b_6451(.a(_w_8353),.q(N6150));
  bfr _b_8877(.a(_w_10779),.q(n494));
  spl2 g1641_s_0(.a(n1641),.q0(n1641_0),.q1(_w_10202));
  and_bb g1537(.a(N137_18),.b(N511_12),.q(_w_13907));
  spl2 g1511_s_0(.a(n1511),.q0(n1511_0),.q1(n1511_1));
  and_bb g157(.a(n143_1),.b(n155_1),.q(_w_10206));
  spl2 g1209_s_0(.a(n1209),.q0(n1209_0),.q1(n1209_1));
  spl2 g768_s_0(.a(n768),.q0(n768_0),.q1(n768_1));
  or_bb g1599(.a(n1597_0),.b(n1598),.q(n1599));
  bfr _b_7906(.a(_w_9808),.q(_w_9809));
  bfr _b_6896(.a(_w_8798),.q(_w_8799));
  bfr _b_4223(.a(_w_6125),.q(_w_6126));
  spl2 g549_s_0(.a(n549),.q0(n549_0),.q1(n549_1));
  bfr _b_14373(.a(_w_16275),.q(_w_16276));
  and_bi g1590(.a(n1588_0),.b(n1589),.q(n1590));
  and_bi g462(.a(n460_0),.b(n461),.q(n462));
  bfr _b_7283(.a(_w_9185),.q(n933));
  bfr _b_7018(.a(_w_8920),.q(_w_8921));
  and_bi g1500(.a(n1499_0),.b(n1462_0),.q(n1500));
  bfr _b_9198(.a(_w_11100),.q(_w_11101));
  bfr _b_9798(.a(_w_11700),.q(_w_11701));
  bfr _b_4584(.a(_w_6486),.q(_w_6487));
  bfr _b_4411(.a(_w_6313),.q(_w_6314));
  and_bb g622(.a(N409_9),.b(N86_12),.q(n622));
  spl2 g1634_s_0(.a(n1634),.q0(n1634_0),.q1(n1634_1));
  bfr _b_9221(.a(_w_11123),.q(_w_11124));
  bfr _b_3726(.a(_w_5628),.q(_w_5629));
  bfr _b_3829(.a(_w_5731),.q(_w_5732));
  spl2 g1098_s_0(.a(n1098),.q0(n1098_0),.q1(n1098_1));
  and_bi g1111(.a(n1064_1),.b(n1109_1),.q(_w_8199));
  or_bb g58(.a(n41_1),.b(n57_0),.q(_w_12487));
  bfr _b_14282(.a(_w_16184),.q(_w_16185));
  bfr _b_5278(.a(_w_7180),.q(_w_7181));
  bfr _b_9681(.a(_w_11583),.q(_w_11584));
  bfr _b_5966(.a(_w_7868),.q(_w_7869));
  spl4L N426_s_1(.a(N426_0),.q0(N426_4),.q1(N426_5),.q2(N426_6),.q3(N426_7));
  and_bb g1231(.a(n1172_1),.b(n1229_1),.q(_w_10283));
  spl2 g1569_s_0(.a(n1569),.q0(n1569_0),.q1(n1569_1));
  bfr _b_6984(.a(_w_8886),.q(_w_8887));
  and_bi g584(.a(n582_0),.b(n583),.q(n584));
  spl2 g807_s_0(.a(n807),.q0(n807_0),.q1(n807_1));
  spl2 g1572_s_0(.a(n1572),.q0(n1572_0),.q1(n1572_1));
  bfr _b_4273(.a(_w_6175),.q(_w_6176));
  bfr _b_7801(.a(_w_9703),.q(_w_9704));
  bfr _b_12007(.a(_w_13909),.q(_w_13910));
  bfr _b_9691(.a(_w_11593),.q(_w_11594));
  and_bi g1116(.a(n1115_0),.b(n1062_0),.q(n1116));
  and_bb g188(.a(N324_8),.b(N69_7),.q(_w_10284));
  bfr _b_10684(.a(_w_12586),.q(_w_12587));
  and_bi g668(.a(n626_1),.b(n666_1),.q(_w_10298));
  and_bb g634(.a(N188_6),.b(N307_15),.q(_w_10299));
  bfr _b_12152(.a(_w_14054),.q(_w_14055));
  and_bb g107(.a(N290_9),.b(N86_4),.q(n107));
  bfr _b_7384(.a(_w_9286),.q(_w_9287));
  and_bi g264(.a(n262_0),.b(n263),.q(n264));
  and_bi g346(.a(n296_1),.b(n344_1),.q(_w_10305));
  bfr _b_3874(.a(_w_5776),.q(_w_5777));
  spl2 g1762_s_0(.a(n1762),.q0(n1762_0),.q1(n1762_1));
  bfr _b_6811(.a(_w_8713),.q(_w_8714));
  bfr _b_9377(.a(_w_11279),.q(_w_11280));
  and_bi g545(.a(n544),.b(n542_0),.q(n545));
  bfr _b_7898(.a(_w_9800),.q(_w_9801));
  spl2 g132_s_0(.a(n132),.q0(n132_0),.q1(n132_1));
  bfr _b_12540(.a(_w_14442),.q(_w_14443));
  bfr _b_8079(.a(_w_9981),.q(_w_9982));
  or_bb g1235(.a(n1233_0),.b(n1234),.q(n1235));
  spl2 g732_s_0(.a(n732),.q0(n732_0),.q1(n732_1));
  bfr _b_9517(.a(_w_11419),.q(_w_11420));
  bfr _b_10222(.a(_w_12124),.q(_w_12125));
  and_bi g982(.a(n980_0),.b(n981),.q(n982));
  bfr _b_12176(.a(_w_14078),.q(n281));
  and_bi g1631(.a(n1629_0),.b(n1630),.q(n1631));
  bfr _b_11078(.a(_w_12980),.q(_w_12981));
  bfr _b_9982(.a(_w_11884),.q(_w_11885));
  and_bi g1432(.a(n1369_1),.b(n1430_1),.q(_w_14613));
  bfr _b_14272(.a(_w_16174),.q(_w_16175));
  or_bb g974(.a(n959_0),.b(n973_0),.q(n974));
  bfr _b_5661(.a(_w_7563),.q(_w_7564));
  bfr _b_11326(.a(_w_13228),.q(_w_13229));
  bfr _b_9761(.a(_w_11663),.q(_w_11664));
  and_bb g257(.a(n243_1),.b(n255_1),.q(_w_10306));
  bfr _b_4228(.a(_w_6130),.q(_w_6131));
  bfr _b_10287(.a(_w_12189),.q(_w_12190));
  bfr _b_4487(.a(_w_6389),.q(n1137_1));
  and_bb g349(.a(n295_1),.b(n347_1),.q(_w_12077));
  bfr _b_5255(.a(_w_7157),.q(_w_7158));
  bfr _b_4059(.a(_w_5961),.q(_w_5962));
  spl2 g1397_s_0(.a(n1397),.q0(n1397_0),.q1(n1397_1));
  bfr _b_3835(.a(_w_5737),.q(_w_5738));
  bfr _b_8321(.a(_w_10223),.q(_w_10224));
  and_bi g1400(.a(n1398_0),.b(n1399),.q(n1400));
  bfr _b_4399(.a(_w_6301),.q(_w_6302));
  and_bb g479(.a(n449_1),.b(n477_1),.q(_w_10439));
  bfr _b_8340(.a(_w_10242),.q(_w_10243));
  bfr _b_8263(.a(_w_10165),.q(_w_10166));
  and_bb g456(.a(n379_1),.b(n455_0),.q(n456));
  or_bb g766(.a(n729_0),.b(n765_0),.q(n766));
  spl2 g1484_s_0(.a(n1484),.q0(n1484_0),.q1(n1484_1));
  bfr _b_5335(.a(_w_7237),.q(_w_7238));
  bfr _b_12918(.a(_w_14820),.q(_w_14821));
  and_bi g1103(.a(n1101_0),.b(n1102),.q(n1103));
  and_bb g175(.a(n137_1),.b(n173_1),.q(_w_10440));
  bfr _b_5808(.a(_w_7710),.q(_w_7711));
  or_bb g992(.a(n953_0),.b(n991_0),.q(n992));
  spl2 g85_s_0(.a(n85),.q0(n85_0),.q1(n85_1));
  and_bi g1798(.a(n1783_1),.b(n1796_1),.q(_w_12514));
  and_bi g562(.a(n536_1),.b(n560_1),.q(_w_10442));
  bfr _b_4648(.a(_w_6550),.q(_w_6551));
  spl2 g712_s_0(.a(n712),.q0(n712_0),.q1(n712_1));
  bfr _b_12642(.a(_w_14544),.q(_w_14545));
  bfr _b_10977(.a(_w_12879),.q(_w_12880));
  spl2 g84_s_0(.a(n84),.q0(n84_0),.q1(n84_1));
  bfr _b_7348(.a(_w_9250),.q(n1627));
  bfr _b_4612(.a(_w_6514),.q(_w_6515));
  spl2 g1602_s_0(.a(n1602),.q0(n1602_0),.q1(n1602_1));
  or_bb g706(.a(n613_0),.b(n705_0),.q(n706));
  bfr _b_3941(.a(_w_5843),.q(_w_5844));
  bfr _b_5554(.a(_w_7456),.q(_w_7457));
  bfr _b_5227(.a(_w_7129),.q(_w_7130));
  or_bb g1009(.a(n1007_0),.b(n1008),.q(n1009));
  and_bb g1711(.a(n1676_1),.b(n1709_1),.q(_w_10452));
  and_bb g306(.a(N120_6),.b(N307_11),.q(_w_10453));
  bfr _b_9976(.a(_w_11878),.q(_w_11879));
  bfr _b_5696(.a(_w_7598),.q(_w_7599));
  and_bi g750(.a(n748_0),.b(n749),.q(n750));
  bfr _b_12979(.a(_w_14881),.q(_w_14882));
  bfr _b_4265(.a(_w_6167),.q(_w_6168));
  and_bb g209(.a(n187_1),.b(n207_1),.q(_w_10559));
  bfr _b_13516(.a(_w_15418),.q(_w_15419));
  and_bb g1064(.a(N154_12),.b(N409_13),.q(n1064));
  and_bi g1431(.a(n1430_0),.b(n1369_0),.q(n1431));
  bfr _b_3450(.a(_w_5352),.q(_w_5353));
  spl2 g510_s_0(.a(n510),.q0(n510_0),.q1(n510_1));
  spl4L N392_s_1(.a(N392_0),.q0(N392_4),.q1(N392_5),.q2(N392_6),.q3(N392_7));
  bfr _b_6354(.a(_w_8256),.q(_w_8257));
  bfr _b_7413(.a(_w_9315),.q(_w_9316));
  spl2 g925_s_0(.a(n925),.q0(n925_0),.q1(n925_1));
  bfr _b_9175(.a(_w_11077),.q(_w_11078));
  bfr _b_10105(.a(_w_12007),.q(_w_12008));
  and_bb g89(.a(n75_1),.b(n87_1),.q(_w_10565));
  bfr _b_4485(.a(_w_6387),.q(_w_6388));
  spl2 g1730_s_0(.a(n1730),.q0(n1730_0),.q1(n1730_1));
  bfr _b_10329(.a(_w_12231),.q(_w_12232));
  and_bi g134(.a(n100_1),.b(n132_1),.q(_w_10566));
  bfr _b_3945(.a(_w_5847),.q(_w_5848));
  spl2 g1692_s_0(.a(n1692),.q0(n1692_0),.q1(_w_10567));
  and_bi g1476(.a(n1475_0),.b(n1470_0),.q(n1476));
  or_bb g1805(.a(n1803_0),.b(n1804),.q(n1805));
  bfr _b_4929(.a(_w_6831),.q(_w_6832));
  and_bi g416(.a(n366_1),.b(n414_1),.q(_w_10571));
  bfr _b_8550(.a(_w_10452),.q(n1711));
  bfr _b_13353(.a(_w_15255),.q(_w_15256));
  bfr _b_10772(.a(_w_12674),.q(_w_12675));
  and_bi g233(.a(n226_1),.b(n229_1),.q(n233));
  bfr _b_3684(.a(_w_5586),.q(_w_5587));
  bfr _b_10407(.a(_w_12309),.q(n1288));
  bfr _b_4310(.a(_w_6212),.q(_w_6213));
  spl2 g1419_s_0(.a(n1419),.q0(n1419_0),.q1(n1419_1));
  bfr _b_9955(.a(_w_11857),.q(_w_11858));
  and_bi g1145(.a(n1143_0),.b(n1144),.q(n1145));
  or_bb g772(.a(n727_0),.b(n771_0),.q(n772));
  spl2 g763_s_0(.a(n763),.q0(n763_0),.q1(n763_1));
  or_bb g1392(.a(n1382_0),.b(n1391_0),.q(n1392));
  bfr _b_4330(.a(_w_6232),.q(_w_6233));
  bfr _b_3934(.a(_w_5836),.q(n739_1));
  and_bi g493(.a(n492_0),.b(n444_0),.q(n493));
  bfr _b_12947(.a(_w_14849),.q(_w_14850));
  and_bi g480(.a(n478_0),.b(n479),.q(n480));
  bfr _b_8736(.a(_w_10638),.q(_w_10639));
  bfr _b_8204(.a(_w_10106),.q(_w_10107));
  bfr _b_12313(.a(_w_14215),.q(_w_14216));
  and_bi g1414(.a(n1375_1),.b(n1412_1),.q(_w_10594));
  bfr _b_13365(.a(_w_15267),.q(_w_15268));
  and_bi g806(.a(n716_1),.b(n804_1),.q(_w_10595));
  spl4L N120_s_0(.a(_w_15526),.q0(N120_0),.q1(_w_9373),.q2(_w_9397),.q3(_w_9453));
  spl2 g546_s_0(.a(n546),.q0(n546_0),.q1(_w_10596));
  bfr _b_4819(.a(_w_6721),.q(_w_6722));
  and_bb g76(.a(N307_6),.b(N35_6),.q(_w_10600));
  spl2 g728_s_0(.a(n728),.q0(n728_0),.q1(n728_1));
  bfr _b_3426(.a(_w_5328),.q(_w_5329));
  spl2 g1554_s_0(.a(n1554),.q0(n1554_0),.q1(n1554_1));
  and_bb g1748(.a(n1737_1),.b(n1746_1),.q(_w_15052));
  bfr _b_5517(.a(_w_7419),.q(_w_7420));
  bfr _b_12807(.a(_w_14709),.q(_w_14710));
  bfr _b_10927(.a(_w_12829),.q(_w_12830));
  bfr _b_4542(.a(_w_6444),.q(_w_6445));
  and_bb g1550(.a(N256_4),.b(N392_19),.q(n1550));
  bfr _b_13653(.a(_w_15555),.q(_w_15556));
  bfr _b_11981(.a(_w_13883),.q(_w_13884));
  bfr _b_7335(.a(_w_9237),.q(_w_9238));
  and_bb g52(.a(N1_7),.b(N324_4),.q(_w_10606));
  bfr _b_6331(.a(_w_8233),.q(_w_8234));
  spl2 g581_s_0(.a(n581),.q0(n581_0),.q1(n581_1));
  spl2 g249_s_0(.a(n249),.q0(n249_0),.q1(n249_1));
  or_bb g484(.a(n447_0),.b(n483_0),.q(n484));
  bfr _b_9407(.a(_w_11309),.q(_w_11310));
  bfr _b_8123(.a(_w_10025),.q(_w_10026));
  or_bb g279(.a(n277_0),.b(n278),.q(n279));
  bfr _b_13612(.a(_w_15514),.q(_w_15515));
  spl2 g1523_s_0(.a(n1523),.q0(n1523_0),.q1(n1523_1));
  bfr _b_13954(.a(_w_15856),.q(_w_15857));
  spl2 g397_s_0(.a(n397),.q0(n397_0),.q1(n397_1));
  spl2 g859_s_0(.a(n859),.q0(n859_0),.q1(n859_1));
  bfr _b_8520(.a(_w_10422),.q(_w_10423));
  spl2 g1330_s_0(.a(n1330),.q0(n1330_0),.q1(n1330_1));
  and_bb g659(.a(n629_1),.b(n657_1),.q(_w_10620));
  bfr _b_6326(.a(_w_8228),.q(n322));
  and_bi g764(.a(n730_1),.b(n762_1),.q(_w_9135));
  spl2 g1318_s_0(.a(n1318),.q0(n1318_0),.q1(n1318_1));
  bfr _b_4367(.a(_w_6269),.q(N120_6));
  spl2 g1384_s_0(.a(n1384),.q0(n1384_0),.q1(n1384_1));
  bfr _b_6617(.a(_w_8519),.q(_w_8520));
  bfr _b_6880(.a(_w_8782),.q(_w_8783));
  spl2 g1497_s_0(.a(n1497),.q0(n1497_0),.q1(_w_7535));
  bfr _b_8908(.a(_w_10810),.q(_w_10811));
  and_bi g132(.a(n130_0),.b(n131),.q(n132));
  bfr _b_14241(.a(_w_16143),.q(_w_16144));
  bfr _b_6522(.a(_w_8424),.q(_w_8425));
  spl2 g1481_s_0(.a(n1481),.q0(n1481_0),.q1(n1481_1));
  bfr _b_10849(.a(_w_12751),.q(_w_12752));
  bfr _b_8109(.a(_w_10011),.q(_w_10012));
  bfr _b_7582(.a(_w_9484),.q(_w_9485));
  spl2 g138_s_0(.a(n138),.q0(n138_0),.q1(n138_1));
  bfr _b_5006(.a(_w_6908),.q(_w_6909));
  and_bi g1619(.a(n1558_1),.b(n1561_1),.q(n1619));
  bfr _b_14235(.a(_w_16137),.q(_w_16138));
  and_bi g358(.a(n292_1),.b(n356_1),.q(_w_10621));
  and_bi g762(.a(n760_0),.b(n761),.q(n762));
  and_bi g166(.a(n140_1),.b(n164_1),.q(_w_10623));
  bfr _b_11615(.a(_w_13517),.q(_w_13518));
  and_bb g287(.a(n233_1),.b(n285_1),.q(_w_10624));
  and_bi g889(.a(n887_0),.b(n888),.q(n889));
  bfr _b_9637(.a(_w_11539),.q(_w_11540));
  and_bi g741(.a(n740),.b(n738_0),.q(n741));
  or_bb g393(.a(n391_0),.b(n392),.q(n393));
  bfr _b_10544(.a(_w_12446),.q(_w_12447));
  bfr _b_6306(.a(_w_8208),.q(_w_8209));
  or_bb g923(.a(n823_0),.b(n922_0),.q(n923));
  and_bi g396(.a(n394_0),.b(n395),.q(n396));
  bfr _b_8509(.a(_w_10411),.q(_w_10412));
  or_bb g1478(.a(n1476_0),.b(n1477),.q(n1478));
  bfr _b_10864(.a(_w_12766),.q(_w_12767));
  spl2 g1229_s_0(.a(n1229),.q0(n1229_0),.q1(n1229_1));
  bfr _b_7221(.a(_w_9123),.q(_w_9124));
  and_bi g972(.a(n960_1),.b(n970_1),.q(_w_10625));
  bfr _b_10036(.a(_w_11938),.q(_w_11939));
  bfr _b_9115(.a(_w_11017),.q(n1516));
  bfr _b_4362(.a(_w_6264),.q(_w_6265));
  bfr _b_11172(.a(_w_13074),.q(_w_13075));
  spl2 g1066_s_0(.a(n1066),.q0(n1066_0),.q1(n1066_1));
  spl2 g1354_s_0(.a(n1354),.q0(n1354_0),.q1(n1354_1));
  bfr _b_4631(.a(_w_6533),.q(_w_6534));
  or_bb g66(.a(n53_0),.b(n65_0),.q(n66));
  bfr _b_5230(.a(_w_7132),.q(_w_7133));
  and_bi g1038(.a(n938_1),.b(n1036_1),.q(_w_10626));
  and_bb g1011(.a(n1009_1),.b(n947_1),.q(_w_8359));
  spl2 g1536_s_0(.a(n1536),.q0(n1536_0),.q1(n1536_1));
  bfr _b_6368(.a(_w_8270),.q(_w_8271));
  spl2 g267_s_0(.a(n267),.q0(n267_0),.q1(n267_1));
  bfr _b_8919(.a(_w_10821),.q(n1126));
  spl2 g1335_s_0(.a(n1335),.q0(n1335_0),.q1(n1335_1));
  and_bi g91(.a(n90_0),.b(n74_0),.q(n91));
  or_bb g156(.a(n143_0),.b(n155_0),.q(n156));
  bfr _b_4248(.a(_w_6150),.q(N171_6));
  bfr _b_10819(.a(_w_12721),.q(_w_12722));
  and_bi g114(.a(n112_0),.b(n113),.q(n114));
  bfr _b_8300(.a(_w_10202),.q(_w_10203));
  bfr _b_14353(.a(_w_16255),.q(_w_16256));
  bfr _b_10878(.a(_w_12780),.q(_w_12781));
  bfr _b_9821(.a(_w_11723),.q(_w_11724));
  bfr _b_4624(.a(_w_6526),.q(_w_6527));
  bfr _b_4578(.a(_w_6480),.q(_w_6481));
  bfr _b_8272(.a(_w_10174),.q(_w_10175));
  bfr _b_10357(.a(_w_12259),.q(_w_12260));
  and_bi g385(.a(n384_0),.b(n376_0),.q(n385));
  bfr _b_5490(.a(_w_7392),.q(_w_7393));
  bfr _b_6995(.a(_w_8897),.q(_w_8898));
  bfr _b_7992(.a(_w_9894),.q(_w_9895));
  bfr _b_8078(.a(_w_9980),.q(_w_9981));
  bfr _b_13089(.a(_w_14991),.q(_w_14992));
  bfr _b_3698(.a(_w_5600),.q(_w_5601));
  spl2 g1548_s_0(.a(n1548),.q0(n1548_0),.q1(n1548_1));
  spl2 g311_s_0(.a(n311),.q0(n311_0),.q1(n311_1));
  bfr _b_5178(.a(_w_7080),.q(_w_7081));
  spl2 g1418_s_0(.a(n1418),.q0(n1418_0),.q1(n1418_1));
  and_bi g1814(.a(n1812_0),.b(n1813),.q(n1814));
  bfr _b_5959(.a(_w_7861),.q(_w_7862));
  and_bb g191(.a(N120_4),.b(N290_11),.q(n191));
  bfr _b_7605(.a(_w_9507),.q(_w_9508));
  and_bi g153(.a(n152_0),.b(n144_0),.q(n153));
  and_bb g182(.a(N18_10),.b(N375_5),.q(_w_10645));
  spl2 g1701_s_0(.a(n1701),.q0(n1701_0),.q1(n1701_1));
  bfr _b_10208(.a(_w_12110),.q(_w_12111));
  spl2 g513_s_0(.a(n513),.q0(n513_0),.q1(n513_1));
  bfr _b_8265(.a(_w_10167),.q(_w_10168));
  spl2 g1518_s_0(.a(n1518),.q0(n1518_0),.q1(n1518_1));
  bfr _b_9188(.a(_w_11090),.q(_w_11091));
  spl2 g276_s_0(.a(n276),.q0(n276_0),.q1(n276_1));
  bfr _b_12998(.a(_w_14900),.q(_w_14901));
  bfr _b_4442(.a(_w_6344),.q(_w_6345));
  bfr _b_9500(.a(_w_11402),.q(_w_11403));
  bfr _b_4869(.a(_w_6771),.q(_w_6772));
  bfr _b_12132(.a(_w_14034),.q(_w_14035));
  and_bi g1438(.a(n1367_1),.b(n1436_1),.q(_w_13756));
  bfr _b_4168(.a(_w_6070),.q(_w_6071));
  and_bb g41(.a(N290_6),.b(N35_4),.q(n41));
  spl2 g1704_s_0(.a(n1704),.q0(n1704_0),.q1(_w_13928));
  spl2 g1383_s_0(.a(n1383),.q0(n1383_0),.q1(n1383_1));
  bfr _b_4928(.a(_w_6830),.q(_w_6831));
  spl2 g377_s_0(.a(n377),.q0(n377_0),.q1(n377_1));
  and_bb g42(.a(n36_1),.b(n41_0),.q(n42));
  and_bi g504(.a(n502_0),.b(n503),.q(n504));
  bfr _b_4275(.a(_w_6177),.q(_w_6178));
  and_bi g811(.a(n810_0),.b(n714_0),.q(n811));
  and_bi g1363(.a(n1357_1),.b(n1360_1),.q(n1363));
  spl2 g496_s_0(.a(n496),.q0(n496_0),.q1(_w_15305));
  and_bi g241(.a(n202_1),.b(n205_1),.q(n241));
  bfr _b_3518(.a(_w_5420),.q(_w_5421));
  bfr _b_10107(.a(_w_12009),.q(_w_12010));
  bfr _b_5428(.a(_w_7330),.q(_w_7331));
  bfr _b_13514(.a(_w_15416),.q(_w_15417));
  bfr _b_10348(.a(_w_12250),.q(_w_12251));
  bfr _b_6673(.a(_w_8575),.q(_w_8576));
  and_bi g321(.a(n320_0),.b(n304_0),.q(n321));
  bfr _b_4813(.a(_w_6715),.q(_w_6716));
  bfr _b_4077(.a(_w_5979),.q(_w_5980));
  bfr _b_13457(.a(_w_15359),.q(_w_15360));
  and_bb g169(.a(n139_1),.b(n167_1),.q(_w_10778));
  and_bi g1852(.a(n1839_1),.b(n1842_1),.q(_w_14614));
  and_bi g81(.a(n80),.b(n78_0),.q(n81));
  and_bi g1164(.a(n1143_1),.b(n1146_1),.q(n1164));
  and_bb g541(.a(N205_4),.b(N290_16),.q(n541));
  bfr _b_9902(.a(_w_11804),.q(N171_3));
  bfr _b_4080(.a(_w_5982),.q(_w_5983));
  bfr _b_4245(.a(_w_6147),.q(_w_6148));
  spl2 g555_s_0(.a(n555),.q0(n555_0),.q1(n555_1));
  and_bi g1331(.a(n1276_1),.b(n1329_1),.q(_w_13015));
  and_bb g1754(.a(n1735_1),.b(n1752_1),.q(_w_14289));
  or_bb g471(.a(n469_0),.b(n470),.q(n471));
  and_bb g364(.a(N35_12),.b(N409_6),.q(n364));
  and_bi g727(.a(n664_1),.b(n667_1),.q(n727));
  or_bb g795(.a(n793_0),.b(n794),.q(n795));
  spl2 g790_s_0(.a(n790),.q0(n790_0),.q1(_w_13980));
  bfr _b_4247(.a(_w_6149),.q(_w_6150));
  spl4L N52_s_1(.a(N52_0),.q0(N52_4),.q1(N52_5),.q2(_w_10781),.q3(_w_10783));
  bfr _b_4678(.a(_w_6580),.q(_w_6581));
  spl2 g1424_s_0(.a(n1424),.q0(n1424_0),.q1(n1424_1));
  and_bb g1052(.a(N511_7),.b(N52_18),.q(_w_10785));
  bfr _b_10541(.a(_w_12443),.q(_w_12444));
  spl2 g1394_s_0(.a(n1394),.q0(n1394_0),.q1(n1394_1));
  or_bb g496(.a(n443_0),.b(n495_0),.q(n496));
  and_bb g1096(.a(n1069_1),.b(n1094_1),.q(_w_10801));
  and_bi g1336(.a(n1335_0),.b(n1274_0),.q(n1336));
  and_bb g1822(.a(N222_6),.b(N511_17),.q(_w_10802));
  and_bb g601(.a(n523_1),.b(n599_1),.q(_w_10818));
  bfr _b_6801(.a(_w_8703),.q(_w_8704));
  and_bb g119(.a(n105_1),.b(n117_1),.q(_w_9686));
  or_bb g676(.a(n623_0),.b(n675_0),.q(n676));
  bfr _b_13280(.a(_w_15182),.q(_w_15183));
  bfr _b_9064(.a(_w_10966),.q(_w_10967));
  or_bb g1496(.a(n1494_0),.b(n1495),.q(n1496));
  bfr _b_8805(.a(_w_10707),.q(_w_10708));
  spl2 g991_s_0(.a(n991),.q0(n991_0),.q1(n991_1));
  and_bi g1402(.a(n1379_1),.b(n1400_1),.q(_w_13577));
  bfr _b_9567(.a(_w_11469),.q(_w_11470));
  and_bi g812(.a(n714_1),.b(n810_1),.q(_w_10819));
  spl4L N222_s_0(.a(N222),.q0(_w_7760),.q1(_w_7809),.q2(_w_7874),.q3(N222_3));
  bfr _b_9930(.a(_w_11832),.q(_w_11833));
  and_bi g451(.a(n388_1),.b(n391_1),.q(n451));
  and_bi g381(.a(n380),.b(n378_0),.q(n381));
  spl2 g243_s_0(.a(n243),.q0(n243_0),.q1(n243_1));
  and_bi g633(.a(n546_1),.b(n549_1),.q(n633));
  spl2 g1797_s_0(.a(n1797),.q0(n1797_0),.q1(n1797_1));
  bfr _b_6564(.a(_w_8466),.q(_w_8467));
  or_bb g162(.a(n141_0),.b(n161_0),.q(n162));
  bfr _b_8209(.a(_w_10111),.q(_w_10112));
  bfr _b_7292(.a(_w_9194),.q(_w_9195));
  bfr _b_13396(.a(_w_15298),.q(_w_15299));
  and_bi g1008(.a(n948_1),.b(n1006_1),.q(_w_10820));
  bfr _b_7405(.a(_w_9307),.q(_w_9308));
  and_bb g630(.a(N154_8),.b(N341_13),.q(n630));
  bfr _b_10994(.a(_w_12896),.q(_w_12897));
  bfr _b_5020(.a(_w_6922),.q(_w_6923));
  bfr _b_12054(.a(_w_13956),.q(n1595));
  bfr _b_9778(.a(_w_11680),.q(_w_11681));
  and_bi g877(.a(n875_0),.b(n876),.q(n877));
  and_bi g604(.a(n522_1),.b(n602_1),.q(_w_9566));
  bfr _b_7604(.a(_w_9506),.q(_w_9507));
  and_bb g108(.a(n107_0),.b(n79_1),.q(n108));
  bfr _b_3888(.a(_w_5790),.q(_w_5791));
  bfr _b_6138(.a(_w_8040),.q(_w_8041));
  bfr _b_13118(.a(_w_15020),.q(_w_15021));
  bfr _b_6394(.a(_w_8296),.q(n1050));
  spl4L N443_s_3(.a(N443_2),.q0(N443_12),.q1(N443_13),.q2(N443_14),.q3(N443_15));
  bfr _b_6463(.a(_w_8365),.q(_w_8366));
  bfr _b_10018(.a(_w_11920),.q(_w_11921));
  bfr _b_10618(.a(_w_12520),.q(_w_12521));
  bfr _b_5630(.a(_w_7532),.q(_w_7533));
  spl2 g1364_s_0(.a(n1364),.q0(n1364_0),.q1(n1364_1));
  bfr _b_6015(.a(_w_7917),.q(_w_7918));
  bfr _b_11822(.a(_w_13724),.q(_w_13725));
  bfr _b_4297(.a(_w_6199),.q(n688_1));
  and_bb g728(.a(N137_10),.b(N375_12),.q(_w_10822));
  bfr _b_3808(.a(_w_5710),.q(_w_5711));
  bfr _b_5008(.a(_w_6910),.q(_w_6911));
  and_bi g1220(.a(n1218_0),.b(n1219),.q(n1220));
  spl2 g1296_s_0(.a(n1296),.q0(n1296_0),.q1(n1296_1));
  spl2 g1187_s_0(.a(n1187),.q0(n1187_0),.q1(n1187_1));
  bfr _b_8062(.a(_w_9964),.q(n869_1));
  and_bi g443(.a(n412_1),.b(n415_1),.q(n443));
  bfr _b_5129(.a(_w_7031),.q(_w_7032));
  bfr _b_4894(.a(_w_6796),.q(_w_6797));
  and_bb g1375(.a(N171_14),.b(N443_14),.q(_w_10839));
  bfr _b_9340(.a(_w_11242),.q(_w_11243));
  bfr _b_9145(.a(_w_11047),.q(_w_11048));
  or_bb g124(.a(n103_0),.b(n123_0),.q(n124));
  bfr _b_4018(.a(_w_5920),.q(_w_5921));
  bfr _b_5999(.a(_w_7901),.q(_w_7902));
  bfr _b_8044(.a(_w_9946),.q(n1621));
  and_bi g265(.a(n264_0),.b(n240_0),.q(n265));
  or_bb g93(.a(n91_0),.b(n92),.q(n93));
  bfr _b_7601(.a(_w_9503),.q(_w_9504));
  bfr _b_3768(.a(_w_5670),.q(_w_5671));
  and_bi g1020(.a(n944_1),.b(n1018_1),.q(_w_10859));
  or_bb g202(.a(n189_0),.b(n201_0),.q(n202));
  bfr _b_7383(.a(_w_9285),.q(_w_9286));
  bfr _b_8584(.a(_w_10486),.q(_w_10487));
  spl3L g146_s_0(.a(n146),.q0(n146_0),.q1(_w_13540),.q2(_w_13542));
  spl2 g886_s_0(.a(n886),.q0(n886_0),.q1(n886_1));
  bfr _b_3876(.a(_w_5778),.q(_w_5779));
  bfr _b_6615(.a(_w_8517),.q(_w_8518));
  bfr _b_11597(.a(_w_13499),.q(_w_13500));
  and_bi g469(.a(n468_0),.b(n452_0),.q(n469));
  bfr _b_11021(.a(_w_12923),.q(_w_12924));
  spl2 g1471_s_0(.a(n1471),.q0(n1471_0),.q1(n1471_1));
  spl2 g1749_s_0(.a(n1749),.q0(n1749_0),.q1(n1749_1));
  and_bi g566(.a(n564_0),.b(n565),.q(n566));
  and_bb g186(.a(N341_7),.b(N52_8),.q(n186));
  bfr _b_13414(.a(_w_15316),.q(n1834));
  and_bi g68(.a(n66_0),.b(n67),.q(n68));
  and_bi g205(.a(n204_0),.b(n188_0),.q(n205));
  bfr _b_3517(.a(_w_5419),.q(_w_5420));
  bfr _b_10190(.a(_w_12092),.q(n352));
  and_bb g851(.a(n848_1),.b(n850),.q(n851));
  bfr _b_14077(.a(_w_15979),.q(_w_15980));
  bfr _b_4200(.a(_w_6102),.q(_w_6103));
  bfr _b_13306(.a(_w_15208),.q(_w_15209));
  bfr _b_6584(.a(_w_8486),.q(_w_8487));
  bfr _b_10791(.a(_w_12693),.q(_w_12694));
  bfr _b_4697(.a(_w_6599),.q(_w_6600));
  bfr _b_3621(.a(_w_5523),.q(_w_5524));
  and_bi g316(.a(n306_1),.b(n314_1),.q(_w_10881));
  bfr _b_11861(.a(_w_13763),.q(_w_13764));
  bfr _b_10680(.a(_w_12582),.q(_w_12583));
  bfr _b_3671(.a(_w_5573),.q(_w_5574));
  bfr _b_14322(.a(_w_16224),.q(_w_16225));
  bfr _b_6794(.a(_w_8696),.q(_w_8697));
  bfr _b_7428(.a(_w_9330),.q(_w_9331));
  spl4L N1_s_4(.a(N1_3),.q0(N1_16),.q1(N1_17),.q2(N1_18),.q3(N1_19));
  and_bi g1097(.a(n1095_0),.b(n1096),.q(n1097));
  and_bb g452(.a(N137_7),.b(N324_12),.q(_w_10895));
  spl2 g1541_s_0(.a(n1541),.q0(n1541_0),.q1(n1541_1));
  bfr _b_7596(.a(_w_9498),.q(_w_9499));
  and_bi g45(.a(n44),.b(n42_0),.q(n45));
  and_bb g848(.a(N256_21),.b(N273_19),.q(n848));
  bfr _b_5218(.a(_w_7120),.q(_w_7121));
  bfr _b_5589(.a(_w_7491),.q(_w_7492));
  bfr _b_4502(.a(_w_6404),.q(_w_6405));
  bfr _b_8308(.a(_w_10210),.q(_w_10211));
  and_bi g500(.a(n442_1),.b(n498_1),.q(_w_10884));
  bfr _b_9220(.a(_w_11122),.q(_w_11123));
  and_bi g1656(.a(n1655_0),.b(n1610_0),.q(n1656));
  bfr _b_9816(.a(_w_11718),.q(_w_11719));
  spl2 g1365_s_0(.a(n1365),.q0(n1365_0),.q1(n1365_1));
  and_bb g56(.a(n43_1),.b(n55_0),.q(n56));
  and_bb g455(.a(N188_4),.b(N290_15),.q(n455));
  bfr _b_3655(.a(_w_5557),.q(_w_5558));
  and_bi g995(.a(n994_0),.b(n952_0),.q(n995));
  bfr _b_12247(.a(_w_14149),.q(_w_14150));
  bfr _b_9564(.a(_w_11466),.q(_w_11467));
  bfr _b_12398(.a(_w_14300),.q(_w_14301));
  spl2 g700_s_0(.a(n700),.q0(n700_0),.q1(_w_10889));
  and_bi g98(.a(n72_1),.b(n96_1),.q(_w_10893));
  and_bb g461(.a(n378_2),.b(n459_1),.q(_w_10894));
  and_bi g266(.a(n240_1),.b(n264_1),.q(_w_10909));
  or_bb g335(.a(n333_0),.b(n334),.q(n335));
  bfr _b_9365(.a(_w_11267),.q(_w_11268));
  and_bi g249(.a(n248),.b(n246_0),.q(n249));
  bfr _b_5744(.a(_w_7646),.q(_w_7647));
  bfr _b_8485(.a(_w_10387),.q(_w_10388));
  spl2 g432_s_0(.a(n432),.q0(n432_0),.q1(n432_1));
  and_bi g1773(.a(n1771_0),.b(n1772),.q(n1773));
  bfr _b_12289(.a(_w_14191),.q(_w_14192));
  bfr _b_8313(.a(_w_10215),.q(_w_10216));
  bfr _b_14341(.a(_w_16243),.q(_w_16244));
  bfr _b_7449(.a(_w_9351),.q(_w_9352));
  bfr _b_3708(.a(_w_5610),.q(_w_5611));
  bfr _b_4791(.a(_w_6693),.q(n156_1));
  spl2 g66_s_0(.a(n66),.q0(n66_0),.q1(_w_10910));
  spl2 g777_s_0(.a(n777),.q0(n777_0),.q1(n777_1));
  bfr _b_9766(.a(_w_11668),.q(_w_11669));
  bfr _b_12250(.a(_w_14152),.q(n1726));
  or_bb g934(.a(n932_0),.b(n933),.q(_w_12629));
  spl2 g307_s_0(.a(n307),.q0(n307_0),.q1(n307_1));
  or_bb g1451(.a(n1449_0),.b(n1450),.q(_w_10914));
  bfr _b_4673(.a(_w_6575),.q(_w_6576));
  and_bi g1604(.a(n1533_1),.b(n1602_1),.q(_w_10955));
  bfr _b_5070(.a(_w_6972),.q(_w_6973));
  bfr _b_4720(.a(_w_6622),.q(_w_6623));
  bfr _b_3554(.a(_w_5456),.q(_w_5457));
  and_bb g628(.a(N137_9),.b(N358_12),.q(_w_10956));
  bfr _b_6966(.a(_w_8868),.q(_w_8869));
  and_bi g239(.a(n208_1),.b(n211_1),.q(n239));
  bfr _b_12173(.a(_w_14075),.q(_w_14076));
  bfr _b_5636(.a(_w_7538),.q(n1497_1));
  spl2 g256_s_0(.a(n256),.q0(n256_0),.q1(_w_6390));
  and_bi g521(.a(n514_1),.b(n517_1),.q(n521));
  spl2 g666_s_0(.a(n666),.q0(n666_0),.q1(n666_1));
  spl2 g1446_s_0(.a(n1446),.q0(n1446_0),.q1(_w_10964));
  and_bi g1847(.a(n1845_0),.b(n1846),.q(n1847));
  spl2 g1844_s_0(.a(n1844),.q0(n1844_0),.q1(n1844_1));
  bfr _b_9642(.a(_w_11544),.q(_w_11545));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  and_bb g749(.a(n735_1),.b(n747_1),.q(_w_10980));
  and_bi g873(.a(n840_1),.b(n871_1),.q(_w_10981));
  and_bi g222(.a(n220_0),.b(n221),.q(n222));
  bfr _b_4242(.a(_w_6144),.q(_w_6145));
  and_bb g389(.a(n375_1),.b(n387_1),.q(_w_10982));
  and_bi g1672(.a(n1659_1),.b(n1662_1),.q(_w_10983));
  bfr _b_3508(.a(_w_5410),.q(_w_5411));
  and_bi g408(.a(n406_0),.b(n407),.q(n408));
  or_bb g868(.a(n866_0),.b(n867),.q(n868));
  spl2 g552_s_0(.a(n552),.q0(n552_0),.q1(_w_11011));
  bfr _b_10828(.a(_w_12730),.q(n284));
  spl2 g1557_s_0(.a(n1557),.q0(n1557_0),.q1(n1557_1));
  bfr _b_12981(.a(_w_14883),.q(_w_14884));
  bfr _b_7814(.a(_w_9716),.q(_w_9717));
  bfr _b_9021(.a(_w_10923),.q(_w_10924));
  or_bb g881(.a(n837_0),.b(n880_0),.q(n881));
  and_bb g1417(.a(n1374_1),.b(n1415_1),.q(_w_13580));
  spl2 g327_s_0(.a(n327),.q0(n327_0),.q1(n327_1));
  or_bb g110(.a(n109_0),.b(n77_1),.q(_w_11015));
  bfr _b_14012(.a(_w_15914),.q(_w_15915));
  or_bb g1004(.a(n1003_0),.b(n949_0),.q(n1004));
  bfr _b_12943(.a(_w_14845),.q(_w_14846));
  and_bi g1281(.a(n1212_1),.b(n1215_1),.q(n1281));
  bfr _b_4562(.a(_w_6464),.q(_w_6465));
  and_bi g70(.a(n52_1),.b(n68_1),.q(_w_11016));
  bfr _b_5645(.a(_w_7547),.q(_w_7548));
  spl2 g830_s_0(.a(n830),.q0(n830_0),.q1(n830_1));
  bfr _b_9325(.a(_w_11227),.q(n1645));
  spl2 g1375_s_0(.a(n1375),.q0(n1375_0),.q1(n1375_1));
  and_bi g1505(.a(n1503_0),.b(n1504),.q(n1505));
  bfr _b_11250(.a(_w_13152),.q(_w_13153));
  bfr _b_6192(.a(_w_8094),.q(_w_8095));
  bfr _b_9137(.a(_w_11039),.q(_w_11040));
  and_bb g946(.a(N103_14),.b(N443_10),.q(_w_11018));
  bfr _b_7112(.a(_w_9014),.q(_w_9015));
  bfr _b_4535(.a(_w_6437),.q(N154_13));
  spl2 g1130_s_0(.a(n1130),.q0(n1130_0),.q1(n1130_1));
  spl2 g1421_s_0(.a(n1421),.q0(n1421_0),.q1(n1421_1));
  or_bb g489(.a(n487_0),.b(n488),.q(n489));
  bfr _b_5412(.a(_w_7314),.q(_w_7315));
  or_bb g478(.a(n449_0),.b(n477_0),.q(n478));
  and_bi g1584(.a(n1582_0),.b(n1583),.q(n1584));
  spl2 g426_s_0(.a(n426),.q0(n426_0),.q1(n426_1));
  or_bb g118(.a(n105_0),.b(n117_0),.q(n118));
  bfr _b_7854(.a(_w_9756),.q(_w_9757));
  bfr _b_7319(.a(_w_9221),.q(n689));
  bfr _b_8351(.a(_w_10253),.q(_w_10254));
  bfr _b_14028(.a(N477),.q(_w_15931));
  bfr _b_4745(.a(_w_6647),.q(_w_6648));
  spl2 g483_s_0(.a(n483),.q0(n483_0),.q1(n483_1));
  or_bb g465(.a(n463_0),.b(n464),.q(n465));
  bfr _b_14037(.a(_w_15939),.q(_w_15940));
  bfr _b_3828(.a(_w_5730),.q(_w_5731));
  or_bb g1308(.a(n1306_0),.b(n1307),.q(n1308));
  bfr _b_7099(.a(_w_9001),.q(_w_9002));
  bfr _b_8296(.a(_w_10198),.q(_w_10199));
  and_bi g1178(.a(n1101_1),.b(n1104_1),.q(n1178));
  bfr _b_13525(.a(_w_15427),.q(_w_15428));
  bfr _b_6247(.a(_w_8149),.q(_w_8150));
  bfr _b_13906(.a(_w_15808),.q(_w_15809));
  bfr _b_9716(.a(_w_11618),.q(n1462));
  or_bb g1100(.a(n1098_0),.b(n1099),.q(n1100));
  and_bi g1830(.a(n1829_0),.b(n1824_0),.q(n1830));
  and_bi g356(.a(n354_0),.b(n355),.q(n356));
  bfr _b_9922(.a(_w_11824),.q(_w_11825));
  bfr _b_6749(.a(_w_8651),.q(_w_8652));
  spl2 g1820_s_0(.a(n1820),.q0(n1820_0),.q1(n1820_1));
  bfr _b_5383(.a(_w_7285),.q(_w_7286));
  and_bi g672(.a(n670_0),.b(n671),.q(n672));
  bfr _b_12463(.a(_w_14365),.q(_w_14366));
  and_bb g1840(.a(n1821_1),.b(n1838_1),.q(_w_13579));
  bfr _b_3559(.a(_w_5461),.q(_w_5462));
  spl2 g1721_s_0(.a(n1721),.q0(n1721_0),.q1(n1721_1));
  spl2 g1115_s_0(.a(n1115),.q0(n1115_0),.q1(n1115_1));
  and_bb g1017(.a(n1015_1),.b(n945_1),.q(_w_11023));
  bfr _b_10291(.a(_w_12193),.q(_w_12194));
  bfr _b_4474(.a(_w_6376),.q(_w_6377));
  spl2 g860_s_0(.a(n860),.q0(n860_0),.q1(n860_1));
  and_bi g86(.a(n76_1),.b(n84_1),.q(_w_11025));
  or_bb g887(.a(n835_0),.b(n886_0),.q(n887));
  bfr _b_7951(.a(_w_9853),.q(_w_9854));
  bfr _b_8050(.a(_w_9952),.q(_w_9953));
  bfr _b_8869(.a(_w_10771),.q(_w_10772));
  bfr _b_9665(.a(_w_11567),.q(_w_11568));
  and_bi g610(.a(n520_1),.b(n608_1),.q(_w_11027));
  and_bb g1535(.a(N120_19),.b(N528_11),.q(_w_11028));
  and_bi g1900(.a(n1895_1),.b(n1899_0),.q(N6287));
  and_bb g1486(.a(n1467_1),.b(n1484_1),.q(_w_13856));
  bfr _b_7747(.a(_w_9649),.q(_w_9650));
  and_bi g375(.a(n312_1),.b(n315_1),.q(n375));
  bfr _b_4687(.a(_w_6589),.q(_w_6590));
  and_bb g125(.a(n103_1),.b(n123_1),.q(_w_11060));
  spl2 g1191_s_0(.a(n1191),.q0(n1191_0),.q1(n1191_1));
  and_bi g126(.a(n124_0),.b(n125),.q(n126));
  and_bi g1724(.a(n1722_0),.b(n1723),.q(n1724));
  bfr _b_7403(.a(_w_9305),.q(_w_9306));
  bfr _b_4705(.a(_w_6607),.q(_w_6608));
  spl2 g942_s_0(.a(n942),.q0(n942_0),.q1(n942_1));
  bfr _b_5801(.a(_w_7703),.q(_w_7704));
  bfr _b_10963(.a(_w_12865),.q(_w_12866));
  or_bb g168(.a(n139_0),.b(n167_0),.q(n168));
  bfr _b_8820(.a(_w_10722),.q(_w_10723));
  and_bb g296(.a(N35_11),.b(N392_6),.q(n296));
  bfr _b_6691(.a(_w_8593),.q(_w_8594));
  bfr _b_12332(.a(_w_14234),.q(n1742));
  bfr _b_9280(.a(_w_11182),.q(_w_11183));
  and_bi g1221(.a(n1220_0),.b(n1175_0),.q(n1221));
  bfr _b_10183(.a(_w_12085),.q(_w_12086));
  spl2 g347_s_0(.a(n347),.q0(n347_0),.q1(n347_1));
  and_bi g1737(.a(n1692_1),.b(n1695_1),.q(n1737));
  and_bi g103(.a(n88_1),.b(n91_1),.q(n103));
  and_bb g1717(.a(n1674_1),.b(n1715_1),.q(_w_11062));
  bfr _b_6195(.a(_w_8097),.q(_w_8098));
  or_bb g388(.a(n375_0),.b(n387_0),.q(n388));
  and_bi g735(.a(n640_1),.b(n643_1),.q(n735));
  and_bb g1738(.a(N239_15),.b(N460_18),.q(_w_9278));
  and_bi g1184(.a(n1083_1),.b(n1086_1),.q(n1184));
  bfr _b_5491(.a(_w_7393),.q(_w_7394));
  spl2 g1884_s_0(.a(n1884),.q0(n1884_0),.q1(n1884_1));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(n153_1));
  or_bb g129(.a(n127_0),.b(n128),.q(n129));
  bfr _b_13943(.a(_w_15845),.q(_w_15846));
  and_bi g474(.a(n472_0),.b(n473),.q(n474));
  bfr _b_4849(.a(_w_6751),.q(_w_6752));
  bfr _b_12897(.a(_w_14799),.q(_w_14800));
  bfr _b_4201(.a(_w_6103),.q(_w_6104));
  bfr _b_11054(.a(_w_12956),.q(_w_12957));
  spl2 g1719_s_0(.a(n1719),.q0(n1719_0),.q1(n1719_1));
  spl2 g421_s_0(.a(n421),.q0(n421_0),.q1(n421_1));
  spl2 g1143_s_0(.a(n1143),.q0(n1143_0),.q1(_w_15291));
  spl4L N443_s_0(.a(_w_15792),.q0(N443_0),.q1(N443_1),.q2(N443_2),.q3(N443_3));
  bfr _b_13430(.a(_w_15332),.q(_w_15333));
  bfr _b_4734(.a(_w_6636),.q(_w_6637));
  or_bb g130(.a(n101_0),.b(n129_0),.q(n130));
  bfr _b_5222(.a(_w_7124),.q(_w_7125));
  bfr _b_9318(.a(_w_11220),.q(_w_11221));
  bfr _b_12423(.a(_w_14325),.q(_w_14326));
  and_bb g1614(.a(N188_16),.b(N477_15),.q(n1614));
  bfr _b_13495(.a(_w_15397),.q(_w_15398));
  and_bi g154(.a(n144_1),.b(n152_1),.q(_w_11081));
  and_bb g900(.a(n831_1),.b(n898_1),.q(_w_11082));
  bfr _b_12140(.a(_w_14042),.q(_w_14043));
  bfr _b_5108(.a(_w_7010),.q(_w_7011));
  or_bb g399(.a(n397_0),.b(n398),.q(n399));
  and_bi g137(.a(n130_1),.b(n133_1),.q(n137));
  bfr _b_12895(.a(_w_14797),.q(_w_14798));
  bfr _b_11465(.a(_w_13367),.q(_w_13368));
  and_bb g1608(.a(N137_19),.b(N528_12),.q(_w_11083));
  spl2 g1233_s_0(.a(n1233),.q0(n1233_0),.q1(n1233_1));
  bfr _b_3812(.a(_w_5714),.q(_w_5715));
  bfr _b_4875(.a(_w_6777),.q(_w_6778));
  spl2 g1140_s_0(.a(n1140),.q0(n1140_0),.q1(n1140_1));
  bfr _b_10338(.a(_w_12240),.q(n1779));
  spl2 g1275_s_0(.a(n1275),.q0(n1275_0),.q1(n1275_1));
  and_bi g1408(.a(n1377_1),.b(n1406_1),.q(_w_11107));
  spl2 g1691_s_0(.a(n1691),.q0(n1691_0),.q1(n1691_1));
  and_bi g751(.a(n750_0),.b(n734_0),.q(n751));
  bfr _b_9097(.a(_w_10999),.q(_w_11000));
  bfr _b_13639(.a(_w_15541),.q(_w_15539));
  bfr _b_11855(.a(_w_13757),.q(_w_13758));
  spl2 g1889_s_0(.a(n1889),.q0(n1889_0),.q1(n1889_1));
  spl2 g1821_s_0(.a(n1821),.q0(n1821_0),.q1(n1821_1));
  and_bb g1510(.a(n1459_1),.b(n1508_1),.q(_w_13868));
  bfr _b_11666(.a(_w_13568),.q(_w_13569));
  spl2 g1729_s_0(.a(n1729),.q0(n1729_0),.q1(n1729_1));
  or_bb g874(.a(n872_0),.b(n873),.q(n874));
  and_bb g140(.a(N341_6),.b(N35_8),.q(n140));
  bfr _b_7466(.a(_w_9368),.q(_w_9369));
  and_bi g1883(.a(n1881_0),.b(n1882),.q(n1883));
  and_bb g1274(.a(N120_16),.b(N477_11),.q(n1274));
  or_bb g857(.a(n845_0),.b(n856_0),.q(n857));
  spl2 g1449_s_0(.a(n1449),.q0(n1449_0),.q1(n1449_1));
  bfr _b_7973(.a(_w_9875),.q(_w_9876));
  spl2 g302_s_0(.a(n302),.q0(n302_0),.q1(n302_1));
  or_bb g318(.a(n305_0),.b(n317_0),.q(n318));
  bfr _b_5950(.a(_w_7852),.q(_w_7853));
  bfr _b_6540(.a(_w_8442),.q(_w_8443));
  bfr _b_7364(.a(_w_9266),.q(_w_9267));
  bfr _b_9731(.a(_w_11633),.q(_w_11634));
  spl2 g1336_s_0(.a(n1336),.q0(n1336_0),.q1(n1336_1));
  bfr _b_4335(.a(_w_6237),.q(_w_6238));
  and_bb g151(.a(n108_2),.b(n149_1),.q(_w_11226));
  bfr _b_4664(.a(_w_6566),.q(_w_6567));
  bfr _b_14033(.a(_w_15935),.q(_w_15936));
  or_bb g1088(.a(n1086_0),.b(n1087),.q(n1088));
  bfr _b_7564(.a(_w_9466),.q(_w_9467));
  bfr _b_12819(.a(_w_14721),.q(_w_14722));
  bfr _b_5010(.a(_w_6912),.q(_w_6913));
  spl4L N35_s_0(.a(_w_15570),.q0(N35_0),.q1(_w_11228),.q2(_w_11252),.q3(_w_11308));
  and_bi g1313(.a(n1282_1),.b(n1311_1),.q(_w_11400));
  bfr _b_5029(.a(_w_6931),.q(_w_6932));
  and_bb g509(.a(n439_1),.b(n507_1),.q(_w_11405));
  bfr _b_4390(.a(_w_6292),.q(_w_6293));
  bfr _b_5984(.a(_w_7886),.q(n456_1));
  bfr _b_13002(.a(_w_14904),.q(_w_14905));
  bfr _b_4235(.a(_w_6137),.q(_w_6138));
  and_bi g1821(.a(n1800_1),.b(n1803_1),.q(n1821));
  or_bb g1124(.a(n1122_0),.b(n1123),.q(n1124));
  bfr _b_11304(.a(_w_13206),.q(_w_13207));
  and_bb g145(.a(N103_4),.b(N290_10),.q(n145));
  or_bb g1508(.a(n1506_0),.b(n1507),.q(n1508));
  and_bi g289(.a(n288_0),.b(n232_0),.q(n289));
  and_bi g1477(.a(n1470_1),.b(n1475_1),.q(_w_11578));
  bfr _b_9249(.a(_w_11151),.q(_w_11152));
  spl2 g775_s_0(.a(n775),.q0(n775_0),.q1(n775_1));
  bfr _b_7489(.a(_w_9391),.q(_w_9392));
  and_bi g422(.a(n364_1),.b(n420_1),.q(_w_15304));
  and_bb g55(.a(N290_7),.b(N52_4),.q(n55));
  bfr _b_9846(.a(_w_11748),.q(_w_11749));
  and_bi g1513(.a(n1458_1),.b(n1511_1),.q(_w_11579));
  bfr _b_5795(.a(_w_7697),.q(_w_7698));
  and_bb g1559(.a(n1548_1),.b(n1557_1),.q(_w_11580));
  bfr _b_13543(.a(_w_15445),.q(_w_15446));
  spl2 g1165_s_0(.a(n1165),.q0(n1165_0),.q1(n1165_1));
  bfr _b_7429(.a(_w_9331),.q(_w_9332));
  bfr _b_7935(.a(_w_9837),.q(_w_9838));
  bfr _b_12175(.a(_w_14077),.q(N6240));
  or_bb g1850(.a(n1848_0),.b(n1849),.q(_w_11581));
  bfr _b_13004(.a(_w_14906),.q(_w_14907));
  bfr _b_4514(.a(_w_6416),.q(_w_6417));
  and_bi g1493(.a(n1491_0),.b(n1492),.q(n1493));
  spl2 g734_s_0(.a(n734),.q0(n734_0),.q1(n734_1));
  bfr _b_7007(.a(_w_8909),.q(_w_8910));
  and_bb g1276(.a(N137_15),.b(N460_12),.q(_w_12412));
  and_bb g834(.a(N120_12),.b(N409_11),.q(n834));
  bfr _b_7472(.a(_w_9374),.q(_w_9375));
  or_bb g638(.a(n541_1),.b(n637_0),.q(_w_11597));
  or_bb g1332(.a(n1330_0),.b(n1331),.q(n1332));
  bfr _b_7249(.a(_w_9151),.q(_w_9152));
  bfr _b_4083(.a(_w_5985),.q(_w_5986));
  bfr _b_6669(.a(_w_8571),.q(_w_8572));
  or_bb g652(.a(n631_0),.b(n651_0),.q(n652));
  and_bb g79(.a(N273_8),.b(N69_5),.q(n79));
  and_bi g463(.a(n462_0),.b(n454_0),.q(n463));
  bfr _b_4216(.a(_w_6118),.q(_w_6119));
  bfr _b_3567(.a(_w_5469),.q(_w_5470));
  bfr _b_9746(.a(_w_11648),.q(_w_11649));
  and_bb g102(.a(N18_8),.b(N341_5),.q(n102));
  bfr _b_7821(.a(_w_9723),.q(_w_9724));
  bfr _b_12681(.a(_w_14583),.q(_w_14584));
  spl2 g1179_s_0(.a(n1179),.q0(n1179_0),.q1(n1179_1));
  spl2 g204_s_0(.a(n204),.q0(n204_0),.q1(n204_1));
  bfr _b_8416(.a(_w_10318),.q(_w_10319));
  spl2 g661_s_0(.a(n661),.q0(n661_0),.q1(n661_1));
  and_bb g1785(.a(N239_16),.b(N477_18),.q(n1785));
  bfr _b_4947(.a(_w_6849),.q(_w_6850));
  bfr _b_3704(.a(_w_5606),.q(_w_5607));
  bfr _b_7760(.a(_w_9662),.q(_w_9663));
  and_bi g434(.a(n360_1),.b(n432_1),.q(_w_11601));
  bfr _b_11369(.a(_w_13271),.q(_w_13272));
  bfr _b_7985(.a(_w_9887),.q(_w_9888));
  or_bb g1211(.a(n1209_0),.b(n1210),.q(n1211));
  spl2 g511_s_0(.a(n511),.q0(n511_0),.q1(n511_1));
  bfr _b_9808(.a(_w_11710),.q(_w_11711));
  or_bb g423(.a(n421_0),.b(n422),.q(n423));
  bfr _b_6963(.a(_w_8865),.q(_w_8866));
  bfr _b_6945(.a(_w_8847),.q(_w_8848));
  bfr _b_4003(.a(_w_5905),.q(_w_5906));
  bfr _b_4882(.a(_w_6784),.q(_w_6785));
  and_bb g1462(.a(N171_15),.b(N460_14),.q(_w_11607));
  bfr _b_5681(.a(_w_7583),.q(_w_7584));
  spl2 g567_s_0(.a(n567),.q0(n567_0),.q1(n567_1));
  bfr _b_9631(.a(_w_11533),.q(_w_11534));
  spl2 g1508_s_0(.a(n1508),.q0(n1508_0),.q1(n1508_1));
  spl2 g998_s_0(.a(n998),.q0(n998_0),.q1(_w_5565));
  spl2 g1124_s_0(.a(n1124),.q0(n1124_0),.q1(n1124_1));
  and_bi g428(.a(n362_1),.b(n426_1),.q(_w_11619));
  bfr _b_10396(.a(_w_12298),.q(_w_12299));
  bfr _b_5371(.a(_w_7273),.q(_w_7274));
  bfr _b_12224(.a(_w_14126),.q(_w_14127));
  spl2 g1254_s_0(.a(n1254),.q0(n1254_0),.q1(_w_11620));
  bfr _b_9968(.a(_w_11870),.q(_w_11871));
  bfr _b_3588(.a(_w_5490),.q(_w_5491));
  bfr _b_9282(.a(_w_11184),.q(_w_11185));
  spl2 g778_s_0(.a(n778),.q0(n778_0),.q1(_w_6313));
  and_bb g948(.a(N120_13),.b(N426_11),.q(n948));
  and_bi g1141(.a(n1054_1),.b(n1139_1),.q(_w_11630));
  bfr _b_7816(.a(_w_9718),.q(_w_9719));
  bfr _b_13669(.a(N358),.q(_w_15572));
  spl2 g642_s_0(.a(n642),.q0(n642_0),.q1(n642_1));
  spl4L N171_s_0(.a(_w_15529),.q0(N171_0),.q1(_w_11637),.q2(_w_11661),.q3(_w_11717));
  bfr _b_9839(.a(_w_11741),.q(_w_11742));
  or_bb g711(.a(n709_0),.b(n710),.q(_w_10207));
  and_bb g431(.a(n361_1),.b(n429_1),.q(_w_11805));
  bfr _b_6293(.a(_w_8195),.q(_w_8196));
  bfr _b_8689(.a(_w_10591),.q(_w_10592));
  or_bb g1344(.a(n1342_0),.b(n1343),.q(n1344));
  bfr _b_10757(.a(_w_12659),.q(_w_12660));
  bfr _b_4589(.a(_w_6491),.q(_w_6492));
  and_bi g841(.a(n754_1),.b(n757_1),.q(n841));
  and_bi g158(.a(n156_0),.b(n157),.q(n158));
  bfr _b_3600(.a(_w_5502),.q(_w_5503));
  and_bi g1842(.a(n1841_0),.b(n1820_0),.q(n1842));
  bfr _b_8902(.a(_w_10804),.q(_w_10805));
  bfr _b_5197(.a(_w_7099),.q(_w_7100));
  spl2 g913_s_0(.a(n913),.q0(n913_0),.q1(n913_1));
  or_bb g917(.a(n825_0),.b(n916_0),.q(n917));
  bfr _b_3823(.a(_w_5725),.q(_w_5726));
  and_bi g1228(.a(n1173_1),.b(n1226_1),.q(_w_11806));
  bfr _b_12045(.a(_w_13947),.q(n992_1));
  and_bb g104(.a(N324_6),.b(N35_7),.q(_w_12012));
  bfr _b_7316(.a(_w_9218),.q(n698));
  bfr _b_7845(.a(_w_9747),.q(_w_9748));
  bfr _b_4670(.a(_w_6572),.q(_w_6573));
  bfr _b_4437(.a(_w_6339),.q(_w_6340));
  bfr _b_10254(.a(_w_12156),.q(_w_12157));
  and_bb g540(.a(N171_6),.b(N307_14),.q(_w_11807));
  and_bi g1524(.a(n1523_0),.b(n1454_0),.q(n1524));
  and_bi g1769(.a(n1730_1),.b(n1767_1),.q(_w_11813));
  bfr _b_14054(.a(_w_15956),.q(_w_15957));
  bfr _b_8327(.a(_w_10229),.q(_w_10230));
  bfr _b_4481(.a(_w_6383),.q(_w_6384));
  bfr _b_9802(.a(_w_11704),.q(_w_11705));
  bfr _b_4603(.a(_w_6505),.q(_w_6506));
  bfr _b_6419(.a(_w_8321),.q(_w_8322));
  bfr _b_3418(.a(_w_5320),.q(_w_5321));
  spl2 g1750_s_0(.a(n1750),.q0(n1750_0),.q1(n1750_1));
  spl2 g1289_s_0(.a(n1289),.q0(n1289_0),.q1(n1289_1));
  bfr _b_10905(.a(_w_12807),.q(_w_12808));
  and_bi g297(.a(n274_1),.b(n277_1),.q(n297));
  spl2 g1097_s_0(.a(n1097),.q0(n1097_0),.q1(n1097_1));
  bfr _b_4770(.a(_w_6672),.q(_w_6673));
  bfr _b_8870(.a(_w_10772),.q(_w_10773));
  and_bi g1110(.a(n1109_0),.b(n1064_0),.q(n1110));
  or_bb g1094(.a(n1092_0),.b(n1093),.q(n1094));
  bfr _b_3656(.a(_w_5558),.q(n1034_1));
  spl2 g1878_s_0(.a(n1878),.q0(n1878_0),.q1(n1878_1));
  bfr _b_3764(.a(_w_5666),.q(_w_5667));
  spl2 g228_s_0(.a(n228),.q0(n228_0),.q1(n228_1));
  and_bi g1523(.a(n1521_0),.b(n1522),.q(n1523));
  bfr _b_13262(.a(_w_15164),.q(_w_15165));
  and_bi g1157(.a(n1155_0),.b(n1156),.q(n1157));
  bfr _b_4082(.a(_w_5984),.q(_w_5985));
  and_bi g1483(.a(n1468_1),.b(n1481_1),.q(_w_11815));
  and_bi g1031(.a(n1030_0),.b(n940_0),.q(n1031));
  and_bb g298(.a(N375_7),.b(N52_10),.q(_w_11816));
  bfr _b_5007(.a(_w_6909),.q(N103_1));
  spl2 g1530_s_0(.a(n1530),.q0(n1530_0),.q1(n1530_1));
  bfr _b_3552(.a(_w_5454),.q(_w_5455));
  bfr _b_8726(.a(_w_10628),.q(n891));
  and_bb g1504(.a(n1461_1),.b(n1502_1),.q(_w_9130));
  bfr _b_6071(.a(_w_7973),.q(_w_7974));
  bfr _b_7356(.a(_w_9258),.q(_w_9259));
  bfr _b_12788(.a(_w_14690),.q(_w_14691));
  or_bb g417(.a(n415_0),.b(n416),.q(n417));
  bfr _b_4148(.a(_w_6050),.q(_w_6051));
  and_bi g586(.a(n528_1),.b(n584_1),.q(_w_9960));
  bfr _b_6991(.a(_w_8893),.q(_w_8894));
  and_bi g994(.a(n992_0),.b(n993),.q(n994));
  bfr _b_5294(.a(_w_7196),.q(_w_7197));
  bfr _b_4657(.a(_w_6559),.q(_w_6560));
  and_bi g486(.a(n484_0),.b(n485),.q(n486));
  bfr _b_8205(.a(_w_10107),.q(_w_10108));
  bfr _b_12564(.a(_w_14466),.q(_w_14467));
  bfr _b_6253(.a(_w_8155),.q(_w_8156));
  bfr _b_8991(.a(_w_10893),.q(n98));
  and_bb g379(.a(N171_5),.b(N273_14),.q(n379));
  bfr _b_10011(.a(_w_11913),.q(_w_11914));
  spl2 g1873_s_0(.a(n1873),.q0(n1873_0),.q1(n1873_1));
  bfr _b_11669(.a(_w_13571),.q(_w_13572));
  and_bi g1044(.a(n936_1),.b(n1042_1),.q(_w_11841));
  and_bb g1058(.a(N103_15),.b(N460_10),.q(_w_12335));
  bfr _b_4480(.a(_w_6382),.q(_w_6383));
  bfr _b_12496(.a(_w_14398),.q(_w_14399));
  bfr _b_3879(.a(_w_5781),.q(_w_5782));
  spl2 g576_s_0(.a(n576),.q0(n576_0),.q1(_w_11842));
  bfr _b_5423(.a(_w_7325),.q(_w_7326));
  and_bi g301(.a(n262_1),.b(n265_1),.q(n301));
  and_bi g926(.a(n925_0),.b(n822_0),.q(n926));
  and_bi g1650(.a(n1649_0),.b(n1612_0),.q(n1650));
  spl2 g265_s_0(.a(n265),.q0(n265_0),.q1(n265_1));
  or_bb g771(.a(n769_0),.b(n770),.q(n771));
  bfr _b_12145(.a(_w_14047),.q(_w_14048));
  bfr _b_7506(.a(_w_9408),.q(_w_9409));
  and_bi g1057(.a(n1016_1),.b(n1019_1),.q(n1057));
  bfr _b_4035(.a(_w_5937),.q(_w_5938));
  or_bb g1016(.a(n1015_0),.b(n945_0),.q(n1016));
  or_bb g1095(.a(n1069_0),.b(n1094_0),.q(n1095));
  bfr _b_12696(.a(_w_14598),.q(_w_14599));
  or_bb g802(.a(n717_0),.b(n801_0),.q(n802));
  bfr _b_13264(.a(_w_15166),.q(_w_15167));
  spl2 g190_s_0(.a(n190),.q0(n190_0),.q1(n190_1));
  bfr _b_6511(.a(_w_8413),.q(_w_8414));
  bfr _b_8025(.a(_w_9927),.q(_w_9928));
  bfr _b_12110(.a(_w_14012),.q(_w_14013));
  and_bb g307(.a(N154_4),.b(N290_13),.q(n307));
  and_bi g1360(.a(n1359_0),.b(n1266_0),.q(n1360));
  bfr _b_11362(.a(_w_13264),.q(_w_13265));
  and_bi g1489(.a(n1466_1),.b(n1487_1),.q(_w_11846));
  and_bi g293(.a(n286_1),.b(n289_1),.q(n293));
  bfr _b_4029(.a(_w_5931),.q(_w_5932));
  bfr _b_13720(.a(_w_15622),.q(_w_15623));
  bfr _b_11619(.a(_w_13521),.q(_w_13522));
  bfr _b_6457(.a(_w_8359),.q(n1011));
  bfr _b_3405(.a(_w_5307),.q(_w_5308));
  bfr _b_5373(.a(_w_7275),.q(_w_7276));
  and_bb g1195(.a(n1184_1),.b(n1193_1),.q(_w_12011));
  and_bb g1181(.a(N205_10),.b(N375_16),.q(_w_9227));
  bfr _b_6146(.a(_w_8048),.q(_w_8049));
  bfr _b_4992(.a(_w_6894),.q(_w_6895));
  and_bb g362(.a(N18_13),.b(N426_5),.q(n362));
  bfr _b_4271(.a(_w_6173),.q(_w_6174));
  bfr _b_10887(.a(_w_12789),.q(_w_12790));
  spl4L N426_s_2(.a(N426_1),.q0(N426_8),.q1(N426_9),.q2(N426_10),.q3(N426_11));
  bfr _b_8838(.a(_w_10740),.q(_w_10741));
  bfr _b_4110(.a(_w_6012),.q(_w_6013));
  or_bb g291(.a(n289_0),.b(n290),.q(_w_10662));
  bfr _b_8936(.a(_w_10838),.q(n47));
  spl2 g1351_s_0(.a(n1351),.q0(n1351_0),.q1(_w_12027));
  and_bi g278(.a(n236_1),.b(n276_1),.q(_w_12031));
  bfr _b_3803(.a(_w_5705),.q(_w_5706));
  or_bb g905(.a(n829_0),.b(n904_0),.q(n905));
  spl2 g982_s_0(.a(n982),.q0(n982_0),.q1(n982_1));
  spl2 g1743_s_0(.a(n1743),.q0(n1743_0),.q1(n1743_1));
  bfr _b_14000(.a(_w_15902),.q(_w_15903));
  bfr _b_6472(.a(_w_8374),.q(_w_8375));
  bfr _b_7467(.a(_w_9369),.q(_w_9370));
  bfr _b_10349(.a(_w_12251),.q(_w_12252));
  bfr _b_4299(.a(_w_6201),.q(_w_6202));
  or_bb g312(.a(n246_1),.b(n311_0),.q(n312));
  and_bb g1399(.a(n1380_1),.b(n1397_1),.q(_w_12033));
  and_bi g1283(.a(n1206_1),.b(n1209_1),.q(n1283));
  bfr _b_9972(.a(_w_11874),.q(_w_11875));
  and_bi g512(.a(n438_1),.b(n510_1),.q(_w_12034));
  and_bi g253(.a(n252_0),.b(n244_0),.q(n253));
  bfr _b_4465(.a(_w_6367),.q(_w_6368));
  bfr _b_11237(.a(_w_13139),.q(_w_13140));
  and_bi g96(.a(n94_0),.b(n95),.q(n96));
  bfr _b_10861(.a(_w_12763),.q(_w_12764));
  bfr _b_3685(.a(_w_5587),.q(_w_5588));
  spl2 g1425_s_0(.a(n1425),.q0(n1425_0),.q1(n1425_1));
  and_bi g1067(.a(n986_1),.b(n989_1),.q(n1067));
  and_bb g761(.a(n731_1),.b(n759_1),.q(_w_12060));
  spl2 g1128_s_0(.a(n1128),.q0(n1128_0),.q1(n1128_1));
  and_bi g498(.a(n496_0),.b(n497),.q(n498));
  and_bi g1449(.a(n1448_0),.b(n1363_0),.q(n1449));
  spl2 g1539_s_0(.a(n1539),.q0(n1539_0),.q1(n1539_1));
  bfr _b_14323(.a(_w_16225),.q(_w_16226));
  bfr _b_13134(.a(_w_15036),.q(_w_15037));
  bfr _b_10163(.a(_w_12065),.q(n328));
  and_bb g37(.a(N1_5),.b(N290_5),.q(n37));
  bfr _b_5303(.a(_w_7205),.q(_w_7206));
  bfr _b_12012(.a(_w_13914),.q(_w_13915));
  bfr _b_5746(.a(_w_7648),.q(_w_7649));
  and_bi g391(.a(n390_0),.b(n374_0),.q(n391));
  and_bb g360(.a(N1_14),.b(N443_4),.q(_w_12061));
  bfr _b_7172(.a(_w_9074),.q(_w_9075));
  bfr _b_4975(.a(_w_6877),.q(N137_3));
  spl2 g1370_s_0(.a(n1370),.q0(n1370_0),.q1(n1370_1));
  and_bi g402(.a(n400_0),.b(n401),.q(n402));
  bfr _b_12885(.a(_w_14787),.q(_w_14788));
  and_bi g763(.a(n762_0),.b(n730_0),.q(n763));
  spl2 g531_s_0(.a(n531),.q0(n531_0),.q1(n531_1));
  bfr _b_9944(.a(_w_11846),.q(n1489));
  bfr _b_6495(.a(_w_8397),.q(_w_8398));
  bfr _b_9042(.a(_w_10944),.q(_w_10945));
  bfr _b_10319(.a(_w_12221),.q(_w_12222));
  bfr _b_4350(.a(_w_6252),.q(_w_6253));
  or_bb g801(.a(n799_0),.b(n800),.q(n801));
  bfr _b_4306(.a(_w_6208),.q(_w_6209));
  bfr _b_5745(.a(_w_7647),.q(_w_7648));
  bfr _b_13844(.a(_w_15746),.q(_w_15747));
  spl2 g1088_s_0(.a(n1088),.q0(n1088_0),.q1(n1088_1));
  or_bb g922(.a(n920_0),.b(n921),.q(n922));
  and_bi g433(.a(n432_0),.b(n360_0),.q(n433));
  bfr _b_7438(.a(_w_9340),.q(_w_9341));
  bfr _b_8577(.a(_w_10479),.q(_w_10480));
  bfr _b_13752(.a(_w_15654),.q(_w_15655));
  bfr _b_8283(.a(_w_10185),.q(_w_10186));
  and_bi g327(.a(n326_0),.b(n302_0),.q(n327));
  and_bi g328(.a(n302_1),.b(n326_1),.q(_w_12065));
  spl2 g1661_s_0(.a(n1661),.q0(n1661_0),.q1(n1661_1));
  bfr _b_13310(.a(_w_15212),.q(_w_15213));
  spl2 g193_s_0(.a(n193),.q0(n193_0),.q1(n193_1));
  bfr _b_3635(.a(_w_5537),.q(_w_5538));
  bfr _b_6739(.a(_w_8641),.q(_w_8642));
  bfr _b_11459(.a(_w_13361),.q(_w_13362));
  spl4L N205_s_2(.a(N205_1),.q0(N205_8),.q1(N205_9),.q2(N205_10),.q3(_w_7996));
  bfr _b_7442(.a(_w_9344),.q(n636_1));
  bfr _b_3718(.a(_w_5620),.q(_w_5621));
  bfr _b_5869(.a(_w_7771),.q(_w_7772));
  and_bb g1304(.a(n1285_1),.b(n1302_1),.q(_w_12066));
  bfr _b_8719(.a(_w_10621),.q(n358));
  bfr _b_4548(.a(_w_6450),.q(_w_6451));
  bfr _b_13603(.a(_w_15505),.q(_w_15506));
  spl2 g1285_s_0(.a(n1285),.q0(n1285_0),.q1(n1285_1));
  bfr _b_13304(.a(_w_15206),.q(_w_15207));
  bfr _b_3797(.a(_w_5699),.q(_w_5700));
  bfr _b_4379(.a(_w_6281),.q(_w_6282));
  bfr _b_9045(.a(_w_10947),.q(_w_10948));
  or_bb g123(.a(n121_0),.b(n122),.q(n123));
  bfr _b_7680(.a(_w_9582),.q(n598));
  bfr _b_13362(.a(_w_15264),.q(_w_15265));
  and_bb g906(.a(n829_1),.b(n904_1),.q(_w_12073));
  bfr _b_5726(.a(_w_7628),.q(_w_7629));
  bfr _b_13622(.a(_w_15524),.q(_w_15522));
  bfr _b_10827(.a(_w_12729),.q(n882));
  bfr _b_3623(.a(_w_5525),.q(_w_5526));
  bfr _b_4764(.a(_w_6666),.q(_w_6667));
  and_bb g1464(.a(N188_14),.b(N443_15),.q(_w_12508));
  spl2 g1542_s_0(.a(n1542),.q0(n1542_0),.q1(n1542_1));
  bfr _b_3757(.a(_w_5659),.q(_w_5660));
  and_bb g343(.a(n297_1),.b(n341_1),.q(_w_12074));
  bfr _b_7965(.a(_w_9867),.q(_w_9868));
  or_bb g856(.a(n854_0),.b(n855),.q(n856));
  and_bb g413(.a(n367_1),.b(n411_1),.q(_w_12075));
  bfr _b_10057(.a(_w_11959),.q(_w_11960));
  and_bi g339(.a(n338_0),.b(n298_0),.q(n339));
  and_bb g246(.a(n193_1),.b(n245_0),.q(n246));
  bfr _b_5788(.a(_w_7690),.q(_w_7691));
  bfr _b_7374(.a(_w_9276),.q(_w_9277));
  bfr _b_3728(.a(_w_5630),.q(_w_5631));
  and_bb g1648(.a(n1613_1),.b(n1646_1),.q(_w_8207));
  bfr _b_4520(.a(_w_6422),.q(_w_6423));
  and_bi g183(.a(n168_1),.b(n171_1),.q(n183));
  bfr _b_10973(.a(_w_12875),.q(_w_12876));
  or_bb g1817(.a(n1815_0),.b(n1816),.q(_w_14541));
  and_bb g446(.a(N375_9),.b(N86_10),.q(_w_12491));
  bfr _b_7321(.a(_w_9223),.q(_w_9224));
  bfr _b_12343(.a(_w_14245),.q(_w_14246));
  bfr _b_12093(.a(_w_13995),.q(_w_13996));
  or_bb g1404(.a(n1378_0),.b(n1403_0),.q(n1404));
  bfr _b_5407(.a(_w_7309),.q(_w_7310));
  and_bi g459(.a(n458),.b(n456_0),.q(n459));
  or_bb g582(.a(n529_0),.b(n581_0),.q(n582));
  bfr _b_13333(.a(_w_15235),.q(_w_15236));
  and_bi g351(.a(n350_0),.b(n294_0),.q(n351));
  spl2 g1618_s_0(.a(n1618),.q0(n1618_0),.q1(n1618_1));
  bfr _b_4752(.a(_w_6654),.q(_w_6655));
  bfr _b_7784(.a(_w_9686),.q(n119));
  and_bb g36(.a(N18_5),.b(N273_5),.q(n36));
  bfr _b_4622(.a(_w_6524),.q(_w_6525));
  spl2 g487_s_0(.a(n487),.q0(n487_0),.q1(n487_1));
  spl2 g1864_s_0(.a(n1864),.q0(n1864_0),.q1(_w_12084));
  bfr _b_7163(.a(_w_9065),.q(_w_9066));
  bfr _b_8039(.a(_w_9941),.q(_w_9942));
  spl2 g1085_s_0(.a(n1085),.q0(n1085_0),.q1(n1085_1));
  bfr _b_8170(.a(_w_10072),.q(_w_10073));
  or_bb g1260(.a(n1162_0),.b(n1259_0),.q(_w_12088));
  and_bi g1819(.a(n1806_1),.b(n1809_1),.q(n1819));
  bfr _b_7659(.a(_w_9561),.q(n1105));
  or_bb g354(.a(n293_0),.b(n353_0),.q(n354));
  bfr _b_13195(.a(_w_15097),.q(_w_15098));
  spl4L N511_s_3(.a(N511_2),.q0(N511_12),.q1(N511_13),.q2(N511_14),.q3(N511_15));
  bfr _b_9183(.a(_w_11085),.q(_w_11086));
  and_bi g111(.a(n110),.b(n108_0),.q(n111));
  and_bi g1311(.a(n1309_0),.b(n1310),.q(n1311));
  or_bb g1033(.a(n1031_0),.b(n1032),.q(n1033));
  bfr _b_7537(.a(_w_9439),.q(_w_9440));
  and_bi g554(.a(n552_0),.b(n553),.q(n554));
  and_bb g1423(.a(n1372_1),.b(n1421_1),.q(_w_12093));
  bfr _b_7943(.a(_w_9845),.q(_w_9846));
  and_bb g355(.a(n293_1),.b(n353_1),.q(_w_12094));
  and_bi g1651(.a(n1612_1),.b(n1649_1),.q(_w_13979));
  and_bi g1227(.a(n1226_0),.b(n1173_0),.q(n1227));
  spl2 g637_s_0(.a(n637),.q0(n637_0),.q1(n637_1));
  bfr _b_5065(.a(_w_6967),.q(_w_6968));
  bfr _b_9034(.a(_w_10936),.q(_w_10937));
  bfr _b_9768(.a(_w_11670),.q(_w_11671));
  and_bi g1841(.a(n1839_0),.b(n1840),.q(n1841));
  bfr _b_3724(.a(_w_5626),.q(N256_5));
  and_bb g653(.a(n631_1),.b(n651_1),.q(_w_12096));
  spl2 g420_s_0(.a(n420),.q0(n420_0),.q1(n420_1));
  spl2 g1732_s_0(.a(n1732),.q0(n1732_0),.q1(n1732_1));
  bfr _b_9368(.a(_w_11270),.q(_w_11271));
  bfr _b_9496(.a(_w_11398),.q(_w_11399));
  or_bb g682(.a(n621_0),.b(n681_0),.q(n682));
  bfr _b_5139(.a(_w_7041),.q(_w_7042));
  or_bb g359(.a(n357_0),.b(n358),.q(_w_12098));
  bfr _b_14227(.a(_w_16129),.q(_w_16130));
  bfr _b_5962(.a(_w_7864),.q(_w_7865));
  and_bb g1213(.a(n1178_1),.b(n1211_1),.q(_w_12206));
  bfr _b_11418(.a(_w_13320),.q(_w_13321));
  and_bi g272(.a(n238_1),.b(n270_1),.q(_w_12211));
  spl2 g1004_s_0(.a(n1004),.q0(n1004_0),.q1(_w_12212));
  spl2 g104_s_0(.a(n104),.q0(n104_0),.q1(n104_1));
  bfr _b_3763(.a(_w_5665),.q(_w_5666));
  bfr _b_6898(.a(_w_8800),.q(_w_8801));
  and_bi g1129(.a(n1058_1),.b(n1127_1),.q(_w_9203));
  and_bi g421(.a(n420_0),.b(n364_0),.q(n421));
  bfr _b_8800(.a(_w_10702),.q(_w_10703));
  bfr _b_9041(.a(_w_10943),.q(_w_10944));
  bfr _b_3832(.a(_w_5734),.q(_w_5735));
  and_bb g1779(.a(N188_19),.b(N528_15),.q(_w_12217));
  bfr _b_6738(.a(_w_8640),.q(_w_8641));
  and_bb g524(.a(N35_14),.b(N443_6),.q(_w_12277));
  and_bi g648(.a(n646_0),.b(n647),.q(n648));
  bfr _b_9426(.a(_w_11328),.q(_w_11329));
  bfr _b_5712(.a(_w_7614),.q(_w_7615));
  spl2 g585_s_0(.a(n585),.q0(n585_0),.q1(n585_1));
  and_bi g883(.a(n881_0),.b(n882),.q(n883));
  and_bb g368(.a(N375_8),.b(N69_10),.q(_w_12281));
  and_bi g1019(.a(n1018_0),.b(n944_0),.q(n1019));
  spl2 g1184_s_0(.a(n1184),.q0(n1184_0),.q1(n1184_1));
  spl2 g1747_s_0(.a(n1747),.q0(n1747_0),.q1(_w_14761));
  spl2 g1131_s_0(.a(n1131),.q0(n1131_0),.q1(_w_12297));
  bfr _b_4962(.a(_w_6864),.q(_w_6865));
  and_bb g1288(.a(N239_9),.b(N358_18),.q(_w_12302));
  bfr _b_4407(.a(_w_6309),.q(_w_6310));
  bfr _b_3522(.a(_w_5424),.q(_w_5425));
  spl2 g1867_s_0(.a(n1867),.q0(n1867_0),.q1(n1867_1));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(n75_1));
  bfr _b_8055(.a(_w_9957),.q(n1349));
  bfr _b_10771(.a(_w_12673),.q(_w_12674));
  and_bb g337(.a(n299_1),.b(n335_1),.q(_w_12310));
  and_bb g370(.a(N358_9),.b(N86_9),.q(_w_12311));
  bfr _b_5169(.a(_w_7071),.q(_w_7072));
  bfr _b_9847(.a(_w_11749),.q(_w_11750));
  and_bb g242(.a(N324_9),.b(N86_7),.q(_w_12319));
  spl2 g1353_s_0(.a(n1353),.q0(n1353_0),.q1(n1353_1));
  bfr _b_7247(.a(_w_9149),.q(_w_9150));
  and_bi g371(.a(n324_1),.b(n327_1),.q(n371));
  bfr _b_6915(.a(_w_8817),.q(_w_8818));
  and_bb g372(.a(N103_8),.b(N341_10),.q(n372));
  bfr _b_7407(.a(_w_9309),.q(_w_9310));
  and_bi g1216(.a(n1177_1),.b(n1214_1),.q(_w_12334));
  bfr _b_4966(.a(_w_6868),.q(_w_6869));
  bfr _b_7590(.a(_w_9492),.q(_w_9493));
  bfr _b_8706(.a(_w_10608),.q(_w_10609));
  and_bi g1073(.a(n968_1),.b(n971_1),.q(n1073));
  bfr _b_12809(.a(_w_14711),.q(_w_14712));
  and_bi g492(.a(n490_0),.b(n491),.q(n492));
  spl2 g516_s_0(.a(n516),.q0(n516_0),.q1(n516_1));
  or_bb g406(.a(n369_0),.b(n405_0),.q(n406));
  and_bi g1361(.a(n1266_1),.b(n1359_1),.q(_w_13447));
  or_bb g387(.a(n385_0),.b(n386),.q(n387));
  bfr _b_13640(.a(N324),.q(_w_15543));
  and_bb g33(.a(N18_4),.b(N290_4),.q(n33));
  and_bi g866(.a(n865_0),.b(n842_0),.q(n866));
  and_bb g319(.a(n305_1),.b(n317_1),.q(_w_12515));
  bfr _b_3541(.a(_w_5443),.q(_w_5444));
  and_bb g366(.a(N392_7),.b(N52_11),.q(n366));
  bfr _b_9934(.a(_w_11836),.q(n695));
  or_bb g1082(.a(n1080_0),.b(n1081),.q(_w_12357));
  spl2 g1122_s_0(.a(n1122),.q0(n1122_0),.q1(n1122_1));
  bfr _b_4039(.a(_w_5941),.q(_w_5942));
  spl2 g1333_s_0(.a(n1333),.q0(n1333_0),.q1(_w_12360));
  and_bi g85(.a(n84_0),.b(n76_0),.q(n85));
  bfr _b_4415(.a(_w_6317),.q(_w_6318));
  bfr _b_6730(.a(_w_8632),.q(_w_8633));
  bfr _b_13407(.a(_w_15309),.q(n340));
  spl2 g813_s_0(.a(n813),.q0(n813_0),.q1(n813_1));
  bfr _b_8136(.a(_w_10038),.q(_w_10039));
  spl2 g1707_s_0(.a(n1707),.q0(n1707_0),.q1(n1707_1));
  bfr _b_5210(.a(_w_7112),.q(_w_7113));
  spl2 g1896_s_0(.a(n1896),.q0(n1896_0),.q1(n1896_1));
  bfr _b_8560(.a(_w_10462),.q(_w_10463));
  bfr _b_4796(.a(_w_6698),.q(_w_6699));
  spl2 g798_s_0(.a(n798),.q0(n798_0),.q1(n798_1));
  and_bi g1266(.a(n1260_1),.b(n1263_1),.q(n1266));
  bfr _b_11288(.a(_w_13190),.q(_w_13191));
  bfr _b_7847(.a(_w_9749),.q(_w_9750));
  bfr _b_6260(.a(_w_8162),.q(_w_8163));
  or_bb g1569(.a(n1567_0),.b(n1568),.q(n1569));
  bfr _b_7140(.a(_w_9042),.q(_w_9043));
  and_bi g850(.a(n737_2),.b(N222_18),.q(_w_12365));
  bfr _b_5849(.a(_w_7751),.q(_w_7752));
  bfr _b_4898(.a(_w_6800),.q(_w_6801));
  and_bi g1519(.a(n1456_1),.b(n1517_1),.q(_w_12367));
  and_bi g920(.a(n919_0),.b(n824_0),.q(n920));
  bfr _b_5974(.a(_w_7876),.q(N273_4));
  spl2 g582_s_0(.a(n582),.q0(n582_0),.q1(_w_6292));
  spl2 g429_s_0(.a(n429),.q0(n429_0),.q1(n429_1));
  and_bi g415(.a(n414_0),.b(n366_0),.q(n415));
  and_bi g798(.a(n796_0),.b(n797),.q(n798));
  and_bi g59(.a(n58),.b(n56_0),.q(n59));
  bfr _b_12196(.a(_w_14098),.q(_w_14099));
  spl4L N528_s_4(.a(N528_3),.q0(N528_16),.q1(N528_17),.q2(N528_18),.q3(N528_19));
  bfr _b_6528(.a(_w_8430),.q(_w_8431));
  and_bb g1893(.a(N256_5),.b(N528_19),.q(_w_12368));
  or_bb g1503(.a(n1461_0),.b(n1502_0),.q(n1503));
  bfr _b_4839(.a(_w_6741),.q(_w_6742));
  bfr _b_12154(.a(_w_14056),.q(_w_14057));
  bfr _b_5322(.a(_w_7224),.q(_w_7225));
  bfr _b_6844(.a(_w_8746),.q(_w_8747));
  bfr _b_11492(.a(_w_13394),.q(_w_13395));
  or_bb g418(.a(n365_0),.b(n417_0),.q(n418));
  spl2 g424_s_0(.a(n424),.q0(n424_0),.q1(_w_8135));
  spl2 g1736_s_0(.a(n1736),.q0(n1736_0),.q1(n1736_1));
  bfr _b_7763(.a(_w_9665),.q(_w_9666));
  and_bi g539(.a(n460_1),.b(n463_1),.q(n539));
  or_bb g424(.a(n363_0),.b(n423_0),.q(n424));
  or_bb g929(.a(n821_0),.b(n928_0),.q(n929));
  and_bi g1804(.a(n1781_1),.b(n1802_1),.q(_w_9209));
  spl2 g1453_s_0(.a(n1453),.q0(n1453_0),.q1(n1453_1));
  bfr _b_10983(.a(_w_12885),.q(_w_12886));
  and_bi g1085(.a(n1083_0),.b(n1084),.q(n1085));
  and_bb g1683(.a(N239_14),.b(N443_18),.q(_w_12397));
  and_bi g561(.a(n560_0),.b(n536_0),.q(n561));
  spl2 g1673_s_0(.a(n1673),.q0(n1673_0),.q1(n1673_1));
  bfr _b_11266(.a(_w_13168),.q(_w_13169));
  spl2 g508_s_0(.a(n508),.q0(n508_0),.q1(_w_12401));
  and_bb g425(.a(n363_1),.b(n423_1),.q(_w_12405));
  spl2 g1591_s_0(.a(n1591),.q0(n1591_0),.q1(n1591_1));
  bfr _b_3574(.a(_w_5476),.q(_w_5477));
  bfr _b_13268(.a(_w_15170),.q(_w_15171));
  and_bi g152(.a(n150_0),.b(n151),.q(n152));
  or_bb g1887(.a(n1877_0),.b(n1886_0),.q(n1887));
  bfr _b_3964(.a(_w_5866),.q(_w_5867));
  bfr _b_6843(.a(_w_8745),.q(_w_8746));
  bfr _b_8629(.a(_w_10531),.q(_w_10532));
  bfr _b_11688(.a(_w_13590),.q(_w_13591));
  and_bi g511(.a(n510_0),.b(n438_0),.q(n511));
  bfr _b_4718(.a(_w_6620),.q(_w_6621));
  bfr _b_6663(.a(_w_8565),.q(_w_8566));
  bfr _b_7686(.a(_w_9588),.q(n383));
  bfr _b_13856(.a(_w_15758),.q(_w_15759));
  bfr _b_13474(.a(_w_15376),.q(_w_15377));
  and_bb g1441(.a(n1366_1),.b(n1439_1),.q(_w_12410));
  spl2 g1824_s_0(.a(n1824),.q0(n1824_0),.q1(n1824_1));
  bfr _b_10158(.a(_w_12060),.q(n761));
  bfr _b_3422(.a(_w_5324),.q(_w_5325));
  bfr _b_10042(.a(_w_11944),.q(_w_11945));
  bfr _b_10687(.a(_w_12589),.q(_w_12590));
  and_bb g83(.a(n56_2),.b(n81_1),.q(_w_12411));
  bfr _b_5602(.a(_w_7504),.q(_w_7505));
  or_bb g490(.a(n445_0),.b(n489_0),.q(n490));
  bfr _b_4829(.a(_w_6731),.q(_w_6732));
  bfr _b_12648(.a(_w_14550),.q(_w_14551));
  bfr _b_8092(.a(_w_9994),.q(_w_9995));
  bfr _b_4126(.a(_w_6028),.q(_w_6029));
  and_bi g1264(.a(n1161_1),.b(n1262_1),.q(_w_13048));
  and_bi g623(.a(n576_1),.b(n579_1),.q(n623));
  bfr _b_3752(.a(_w_5654),.q(_w_5655));
  and_bi g679(.a(n678_0),.b(n622_0),.q(n679));
  bfr _b_7006(.a(_w_8908),.q(_w_8909));
  bfr _b_5310(.a(_w_7212),.q(_w_7213));
  bfr _b_9991(.a(_w_11893),.q(_w_11894));
  bfr _b_7865(.a(_w_9767),.q(_w_9768));
  bfr _b_9246(.a(_w_11148),.q(_w_11149));
  bfr _b_4628(.a(_w_6530),.q(_w_6531));
  bfr _b_8673(.a(_w_10575),.q(_w_10576));
  and_bb g302(.a(N341_9),.b(N86_8),.q(n302));
  and_bi g427(.a(n426_0),.b(n362_0),.q(n427));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  and_bb g1405(.a(n1378_1),.b(n1403_1),.q(_w_12424));
  bfr _b_3863(.a(_w_5765),.q(_w_5766));
  bfr _b_7390(.a(_w_9292),.q(n559));
  spl2 g1622_s_0(.a(n1622),.q0(n1622_0),.q1(n1622_1));
  and_bi g482(.a(n448_1),.b(n480_1),.q(_w_12425));
  bfr _b_13273(.a(_w_15175),.q(_w_15176));
  bfr _b_8152(.a(_w_10054),.q(_w_10055));
  bfr _b_8444(.a(_w_10346),.q(_w_10347));
  bfr _b_10185(.a(_w_12087),.q(n1864_1));
  bfr _b_4654(.a(_w_6556),.q(_w_6557));
  bfr _b_12500(.a(_w_14402),.q(_w_14403));
  spl2 g1206_s_0(.a(n1206),.q0(n1206_0),.q1(_w_15300));
  spl2 g336_s_0(.a(n336),.q0(n336_0),.q1(_w_12426));
  bfr _b_6310(.a(_w_8212),.q(_w_8213));
  spl2 g318_s_0(.a(n318),.q0(n318_0),.q1(_w_12430));
  bfr _b_10970(.a(_w_12872),.q(_w_12873));
  and_bi g1540(.a(n1503_1),.b(n1506_1),.q(n1540));
  bfr _b_7074(.a(_w_8976),.q(_w_8977));
  and_bb g240(.a(N341_8),.b(N69_8),.q(n240));
  spl2 g922_s_0(.a(n922),.q0(n922_0),.q1(n922_1));
  bfr _b_10295(.a(_w_12197),.q(_w_12198));
  spl2 g960_s_0(.a(n960),.q0(n960_0),.q1(n960_1));
  bfr _b_5885(.a(_w_7787),.q(_w_7788));
  spl2 g1731_s_0(.a(n1731),.q0(n1731_0),.q1(n1731_1));
  and_bi g1662(.a(n1661_0),.b(n1608_0),.q(n1662));
  spl2 g159_s_0(.a(n159),.q0(n159_0),.q1(n159_1));
  bfr _b_11989(.a(_w_13891),.q(_w_13892));
  bfr _b_4024(.a(_w_5926),.q(_w_5927));
  spl2 g87_s_0(.a(n87),.q0(n87_0),.q1(n87_1));
  and_bi g1615(.a(n1570_1),.b(n1573_1),.q(n1615));
  spl2 g1125_s_0(.a(n1125),.q0(n1125_0),.q1(_w_10860));
  and_bi g1517(.a(n1515_0),.b(n1516),.q(n1517));
  bfr _b_4611(.a(_w_6513),.q(_w_6514));
  bfr _b_4181(.a(_w_6083),.q(_w_6084));
  bfr _b_7444(.a(_w_9346),.q(n636_2));
  bfr _b_8816(.a(_w_10718),.q(_w_10719));
  bfr _b_6849(.a(_w_8751),.q(_w_8752));
  and_bb g450(.a(N120_8),.b(N341_11),.q(n450));
  bfr _b_4073(.a(_w_5975),.q(_w_5976));
  bfr _b_13704(.a(_w_15606),.q(_w_15607));
  bfr _b_10592(.a(_w_12494),.q(_w_12495));
  bfr _b_8765(.a(_w_10667),.q(_w_10668));
  and_bi g1134(.a(n1133_0),.b(n1056_0),.q(n1134));
  spl2 g1371_s_0(.a(n1371),.q0(n1371_0),.q1(n1371_1));
  bfr _b_5556(.a(_w_7458),.q(_w_7459));
  bfr _b_6758(.a(_w_8660),.q(_w_8661));
  and_bb g824(.a(N35_17),.b(N494_6),.q(_w_12478));
  bfr _b_7265(.a(_w_9167),.q(_w_9168));
  and_bi g352(.a(n294_1),.b(n350_1),.q(_w_12092));
  or_bb g460(.a(n378_1),.b(n459_0),.q(n460));
  bfr _b_4091(.a(_w_5993),.q(_w_5994));
  and_bi g1239(.a(n1238_0),.b(n1169_0),.q(n1239));
  spl2 g462_s_0(.a(n462),.q0(n462_0),.q1(n462_1));
  bfr _b_5856(.a(_w_7758),.q(_w_7759));
  bfr _b_5009(.a(_w_6911),.q(_w_6912));
  spl2 g1459_s_0(.a(n1459),.q0(n1459_0),.q1(n1459_1));
  and_bi g230(.a(n180_1),.b(n228_1),.q(_w_12488));
  bfr _b_13054(.a(_w_14956),.q(_w_14957));
  bfr _b_7245(.a(_w_9147),.q(_w_9148));
  and_bi g139(.a(n124_1),.b(n127_1),.q(n139));
  or_bb g155(.a(n153_0),.b(n154),.q(n155));
  and_bb g1120(.a(n1061_1),.b(n1118_1),.q(_w_12489));
  spl2 g1315_s_0(.a(n1315),.q0(n1315_0),.q1(_w_11401));
  bfr _b_7796(.a(_w_9698),.q(_w_9699));
  bfr _b_7941(.a(_w_9843),.q(_w_9844));
  bfr _b_4286(.a(_w_6188),.q(_w_6189));
  or_bb g1259(.a(n1257_0),.b(n1258),.q(n1259));
  and_bi g181(.a(n174_1),.b(n177_1),.q(n181));
  bfr _b_6914(.a(_w_8816),.q(_w_8817));
  bfr _b_9083(.a(_w_10985),.q(_w_10986));
  and_bi g481(.a(n480_0),.b(n448_0),.q(n481));
  and_bb g378(.a(n309_1),.b(n377_0),.q(n378));
  bfr _b_9061(.a(_w_10963),.q(n628));
  bfr _b_13914(.a(_w_15816),.q(_w_15817));
  bfr _b_13852(.a(_w_15754),.q(_w_15755));
  spl2 g1468_s_0(.a(n1468),.q0(n1468_0),.q1(n1468_1));
  and_bi g488(.a(n446_1),.b(n486_1),.q(_w_12507));
  or_bb g495(.a(n493_0),.b(n494),.q(n495));
  bfr _b_4820(.a(_w_6722),.q(_w_6723));
  and_bb g503(.a(n441_1),.b(n501_1),.q(_w_12512));
  bfr _b_3880(.a(_w_5782),.q(_w_5783));
  spl2 g53_s_0(.a(n53),.q0(n53_0),.q1(n53_1));
  bfr _b_3448(.a(_w_5350),.q(_w_5351));
  bfr _b_12192(.a(_w_14094),.q(_w_14095));
  or_bb g760(.a(n731_0),.b(n759_0),.q(n760));
  and_bb g136(.a(N1_10),.b(N375_4),.q(_w_10629));
  and_bb g497(.a(n443_1),.b(n495_1),.q(_w_12516));
  and_bi g1079(.a(n1077_0),.b(n1078),.q(n1079));
  bfr _b_5043(.a(_w_6945),.q(_w_6946));
  bfr _b_7252(.a(_w_9154),.q(_w_9155));
  spl2 g606_s_0(.a(n606),.q0(n606_0),.q1(_w_6305));
  or_bb g508(.a(n439_0),.b(n507_0),.q(n508));
  and_bb g636(.a(n543_1),.b(n635_0),.q(n636));
  bfr _b_4428(.a(_w_6330),.q(_w_6331));
  bfr _b_4210(.a(_w_6112),.q(N171_14));
  bfr _b_11376(.a(_w_13278),.q(_w_13279));
  bfr _b_3675(.a(_w_5577),.q(_w_5578));
  and_bi g75(.a(n60_1),.b(n63_1),.q(n75));
  bfr _b_9366(.a(_w_11268),.q(_w_11269));
  and_bi g1561(.a(n1560_0),.b(n1547_0),.q(n1561));
  and_bb g515(.a(n437_1),.b(n513_1),.q(_w_12518));
  bfr _b_12616(.a(_w_14518),.q(_w_14519));
  spl2 g1833_s_0(.a(n1833),.q0(n1833_0),.q1(_w_12519));
  bfr _b_4079(.a(_w_5981),.q(_w_5982));
  bfr _b_4546(.a(_w_6448),.q(_w_6449));
  bfr _b_7406(.a(_w_9308),.q(_w_9309));
  bfr _b_6454(.a(_w_8356),.q(n1026));
  bfr _b_6408(.a(_w_8310),.q(_w_8311));
  bfr _b_4150(.a(_w_6052),.q(_w_6053));
  bfr _b_6026(.a(_w_7928),.q(_w_7929));
  spl2 g781_s_0(.a(n781),.q0(n781_0),.q1(n781_1));
  bfr _b_6205(.a(_w_8107),.q(_w_8108));
  bfr _b_11525(.a(_w_13427),.q(_w_13428));
  bfr _b_3412(.a(_w_5314),.q(n1083_1));
  bfr _b_8704(.a(_w_10606),.q(_w_10607));
  or_bb g519(.a(n517_0),.b(n518),.q(_w_12524));
  bfr _b_4615(.a(_w_6517),.q(_w_6518));
  bfr _b_4509(.a(_w_6411),.q(_w_6412));
  bfr _b_7675(.a(_w_9577),.q(n1858_1));
  bfr _b_4488(.a(_w_6390),.q(_w_6391));
  and_bb g522(.a(N18_15),.b(N460_5),.q(_w_12617));
  bfr _b_13411(.a(_w_15313),.q(_w_15314));
  bfr _b_10960(.a(_w_12862),.q(N86_7));
  bfr _b_9053(.a(_w_10955),.q(n1604));
  spl4L N307_s_0(.a(_w_15539),.q0(N307_0),.q1(N307_1),.q2(N307_2),.q3(N307_3));
  bfr _b_5499(.a(_w_7401),.q(_w_7402));
  bfr _b_3722(.a(_w_5624),.q(_w_5625));
  and_bb g146(.a(n109_1),.b(n145_0),.q(n146));
  bfr _b_8948(.a(_w_10850),.q(_w_10851));
  spl4L N86_s_3(.a(N86_2),.q0(N86_12),.q1(_w_12689),.q2(_w_12697),.q3(_w_12709));
  and_bi g1579(.a(n1578_0),.b(n1541_0),.q(n1579));
  bfr _b_4566(.a(_w_6468),.q(_w_6469));
  spl2 g1183_s_0(.a(n1183),.q0(n1183_0),.q1(n1183_1));
  and_bb g942(.a(N477_8),.b(N69_16),.q(n942));
  bfr _b_4643(.a(_w_6545),.q(N154_2));
  bfr _b_4803(.a(_w_6705),.q(N426_19));
  bfr _b_6313(.a(_w_8215),.q(n184));
  and_bi g953(.a(n875_1),.b(n878_1),.q(n953));
  and_bb g528(.a(N409_8),.b(N69_12),.q(n528));
  bfr _b_8612(.a(_w_10514),.q(_w_10515));
  bfr _b_9727(.a(_w_11629),.q(n203));
  or_bb g429(.a(n427_0),.b(n428),.q(n429));
  and_bi g1000(.a(n998_0),.b(n999),.q(n1000));
  spl2 g1406_s_0(.a(n1406),.q0(n1406_0),.q1(n1406_1));
  and_bi g529(.a(n490_1),.b(n493_1),.q(n529));
  and_bi g531(.a(n484_1),.b(n487_1),.q(n531));
  or_bb g483(.a(n481_0),.b(n482),.q(n483));
  bfr _b_4590(.a(_w_6492),.q(_w_6493));
  spl2 g1277_s_0(.a(n1277),.q0(n1277_0),.q1(n1277_1));
  bfr _b_12641(.a(_w_14543),.q(_w_14544));
  and_bi g1542(.a(n1497_1),.b(n1500_1),.q(n1542));
  bfr _b_9935(.a(_w_11837),.q(_w_11838));
  spl2 g573_s_0(.a(n573),.q0(n573_0),.q1(n573_1));
  or_bb g1015(.a(n1013_0),.b(n1014),.q(n1015));
  bfr _b_9984(.a(_w_11886),.q(_w_11887));
  spl2 g745_s_0(.a(n745),.q0(n745_0),.q1(n745_1));
  bfr _b_14248(.a(_w_16150),.q(_w_16151));
  and_bb g882(.a(n837_1),.b(n880_1),.q(_w_12729));
  and_bi g535(.a(n472_1),.b(n475_1),.q(n535));
  and_bi g284(.a(n234_1),.b(n282_1),.q(_w_12730));
  and_bb g536(.a(N137_8),.b(N341_12),.q(n536));
  bfr _b_8297(.a(_w_10199),.q(n1384));
  bfr _b_13131(.a(_w_15033),.q(_w_15034));
  bfr _b_9800(.a(_w_11702),.q(_w_11703));
  and_bi g1725(.a(n1724_0),.b(n1671_0),.q(n1725));
  bfr _b_3657(.a(_w_5559),.q(_w_5560));
  and_bi g549(.a(n548_0),.b(n540_0),.q(n549));
  and_bb g683(.a(n621_1),.b(n681_1),.q(_w_9243));
  bfr _b_4371(.a(_w_6273),.q(_w_6274));
  bfr _b_6435(.a(_w_8337),.q(_w_8338));
  bfr _b_8267(.a(_w_10169),.q(_w_10170));
  spl2 g1134_s_0(.a(n1134),.q0(n1134_0),.q1(n1134_1));
  bfr _b_3570(.a(_w_5472),.q(_w_5473));
  spl2 g612_s_0(.a(n612),.q0(n612_0),.q1(n612_1));
  and_bi g404(.a(n370_1),.b(n402_1),.q(_w_12732));
  bfr _b_12879(.a(_w_14781),.q(_w_14782));
  bfr _b_9405(.a(_w_11307),.q(N35_2));
  or_bb g552(.a(n539_0),.b(n551_0),.q(n552));
  or_bb g255(.a(n253_0),.b(n254),.q(n255));
  bfr _b_12688(.a(_w_14590),.q(_w_14591));
  and_bb g1828(.a(n1825_1),.b(n1826_1),.q(_w_12824));
  and_bi g903(.a(n830_1),.b(n901_1),.q(_w_12825));
  and_bb g876(.a(n839_1),.b(n874_1),.q(_w_12826));
  bfr _b_4430(.a(_w_6332),.q(_w_6333));
  bfr _b_6051(.a(_w_7953),.q(N188_6));
  bfr _b_12171(.a(_w_14073),.q(_w_14074));
  spl2 g725_s_0(.a(n725),.q0(n725_0),.q1(n725_1));
  bfr _b_5238(.a(_w_7140),.q(_w_7141));
  and_bb g1225(.a(n1174_1),.b(n1223_1),.q(_w_9134));
  and_bi g977(.a(n976_0),.b(n958_0),.q(n977));
  bfr _b_9903(.a(_w_11805),.q(n431));
  bfr _b_9066(.a(_w_10968),.q(_w_10969));
  bfr _b_10075(.a(_w_11977),.q(_w_11978));
  bfr _b_3912(.a(_w_5814),.q(N256_1));
  and_bi g560(.a(n558_0),.b(n559),.q(n560));
  spl4L N307_s_3(.a(N307_2),.q0(N307_12),.q1(N307_13),.q2(N307_14),.q3(N307_15));
  bfr _b_11765(.a(_w_13667),.q(_w_13668));
  bfr _b_9714(.a(_w_11616),.q(_w_11617));
  or_bb g501(.a(n499_0),.b(n500),.q(n501));
  or_bb g569(.a(n567_0),.b(n568),.q(n569));
  bfr _b_5015(.a(_w_6917),.q(_w_6918));
  bfr _b_11384(.a(_w_13286),.q(_w_13287));
  spl2 g1203_s_0(.a(n1203),.q0(n1203_0),.q1(n1203_1));
  and_bi g871(.a(n869_0),.b(n870),.q(n871));
  spl2 g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1));
  and_bi g1086(.a(n1085_0),.b(n1072_0),.q(n1086));
  bfr _b_14346(.a(_w_16248),.q(_w_16249));
  bfr _b_12237(.a(_w_14139),.q(_w_14140));
  bfr _b_7115(.a(_w_9017),.q(_w_9018));
  bfr _b_9635(.a(_w_11537),.q(_w_11538));
  bfr _b_5022(.a(_w_6924),.q(_w_6925));
  bfr _b_10022(.a(_w_11924),.q(_w_11925));
  or_bb g570(.a(n533_0),.b(n569_0),.q(n570));
  and_bb g1742(.a(n1739_1),.b(n1740_1),.q(_w_14234));
  bfr _b_3939(.a(_w_5841),.q(_w_5842));
  spl2 g1308_s_0(.a(n1308),.q0(n1308_0),.q1(n1308_1));
  or_bb g1623(.a(n1621_0),.b(n1622_0),.q(n1623));
  bfr _b_4127(.a(_w_6029),.q(_w_6030));
  bfr _b_6256(.a(_w_8158),.q(_w_8159));
  and_bb g714(.a(N18_17),.b(N494_5),.q(_w_12841));
  bfr _b_9415(.a(_w_11317),.q(_w_11318));
  bfr _b_7294(.a(_w_9196),.q(_w_9197));
  bfr _b_4098(.a(_w_6000),.q(_w_6001));
  bfr _b_4597(.a(_w_6499),.q(_w_6500));
  spl2 g384_s_0(.a(n384),.q0(n384_0),.q1(n384_1));
  spl2 g1496_s_0(.a(n1496),.q0(n1496_0),.q1(n1496_1));
  or_bb g1143(.a(n1053_0),.b(n1142_0),.q(n1143));
  bfr _b_13824(.a(_w_15726),.q(_w_15670));
  bfr _b_3482(.a(_w_5384),.q(_w_5385));
  and_bi g523(.a(n508_1),.b(n511_1),.q(n523));
  spl2 g57_s_0(.a(n57),.q0(n57_0),.q1(n57_1));
  bfr _b_11053(.a(_w_12955),.q(n1473_1));
  bfr _b_7560(.a(_w_9462),.q(_w_9463));
  and_bb g1144(.a(n1053_1),.b(n1142_1),.q(_w_12850));
  bfr _b_7787(.a(_w_9689),.q(_w_9690));
  bfr _b_3756(.a(_w_5658),.q(_w_5659));
  spl2 g1392_s_0(.a(n1392),.q0(n1392_0),.q1(_w_12851));
  bfr _b_6905(.a(_w_8807),.q(n113));
  bfr _b_6438(.a(_w_8340),.q(_w_8341));
  bfr _b_14295(.a(N52),.q(_w_16197));
  bfr _b_10633(.a(_w_12535),.q(_w_12536));
  bfr _b_4852(.a(_w_6754),.q(_w_6755));
  bfr _b_12185(.a(_w_14087),.q(_w_14088));
  bfr _b_4558(.a(_w_6460),.q(_w_6461));
  bfr _b_8664(.a(_w_10566),.q(n134));
  spl4L N477_s_4(.a(N477_3),.q0(N477_16),.q1(N477_17),.q2(N477_18),.q3(N477_19));
  bfr _b_13001(.a(_w_14903),.q(_w_14904));
  spl2 g1262_s_0(.a(n1262),.q0(n1262_0),.q1(n1262_1));
  and_bb g1150(.a(n1051_1),.b(n1148_1),.q(_w_12855));
  and_bi g189(.a(n150_1),.b(n153_1),.q(n189));
  bfr _b_13293(.a(_w_15195),.q(_w_15196));
  bfr _b_9322(.a(_w_11224),.q(_w_11225));
  spl2 g1217_s_0(.a(n1217),.q0(n1217_0),.q1(n1217_1));
  and_bi g1151(.a(n1149_0),.b(n1150),.q(n1151));
  bfr _b_3705(.a(_w_5607),.q(_w_5608));
  bfr _b_5037(.a(_w_6939),.q(_w_6940));
  bfr _b_11477(.a(_w_13379),.q(_w_13380));
  spl2 g618_s_0(.a(n618),.q0(n618_0),.q1(n618_1));
  bfr _b_5162(.a(_w_7064),.q(_w_7065));
  or_bb g1403(.a(n1401_0),.b(n1402),.q(n1403));
  bfr _b_5529(.a(_w_7431),.q(_w_7432));
  and_bb g1261(.a(n1162_1),.b(n1259_1),.q(_w_13039));
  bfr _b_4782(.a(_w_6684),.q(_w_6685));
  bfr _b_8951(.a(_w_10853),.q(_w_10854));
  and_bi g847(.a(n738_1),.b(N256_13),.q(n847));
  bfr _b_13190(.a(_w_15092),.q(n1327_1));
  bfr _b_10774(.a(_w_12676),.q(_w_12677));
  and_bb g1268(.a(N528_8),.b(N69_19),.q(_w_12864));
  bfr _b_3734(.a(_w_5636),.q(_w_5637));
  and_bi g1159(.a(n1046_2),.b(n1157_1),.q(_w_12888));
  bfr _b_4324(.a(_w_6226),.q(_w_6227));
  spl2 g252_s_0(.a(n252),.q0(n252_0),.q1(n252_1));
  bfr _b_11327(.a(_w_13229),.q(_w_13230));
  bfr _b_7635(.a(_w_9537),.q(_w_9538));
  bfr _b_4014(.a(_w_5916),.q(_w_5917));
  and_bi g149(.a(n148),.b(n146_0),.q(n149));
  bfr _b_9783(.a(_w_11685),.q(_w_11686));
  bfr _b_10230(.a(_w_12132),.q(_w_12133));
  bfr _b_14229(.a(_w_16131),.q(_w_16132));
  bfr _b_13764(.a(_w_15666),.q(_w_15667));
  and_bb g1163(.a(N52_19),.b(N528_7),.q(_w_12889));
  bfr _b_11425(.a(_w_13327),.q(_w_13328));
  bfr _b_3989(.a(_w_5891),.q(_w_5892));
  and_bb g1165(.a(N511_8),.b(N69_18),.q(_w_12914));
  and_bi g1166(.a(n1137_1),.b(n1140_1),.q(n1166));
  bfr _b_5324(.a(_w_7226),.q(_w_7227));
  and_bb g1169(.a(N103_16),.b(N477_10),.q(n1169));
  bfr _b_14314(.a(_w_16216),.q(_w_16217));
  bfr _b_9874(.a(_w_11776),.q(_w_11777));
  bfr _b_12637(.a(_w_14539),.q(n532));
  bfr _b_5048(.a(_w_6950),.q(_w_6951));
  and_bb g304(.a(N103_7),.b(N324_10),.q(_w_12938));
  bfr _b_5444(.a(_w_7346),.q(_w_7347));
  bfr _b_10642(.a(_w_12544),.q(_w_12545));
  and_bi g1172(.a(n1119_1),.b(n1122_1),.q(n1172));
  bfr _b_14258(.a(_w_16160),.q(_w_16161));
  bfr _b_5096(.a(_w_6998),.q(_w_6999));
  and_bb g1571(.a(n1544_1),.b(n1569_1),.q(_w_11628));
  bfr _b_6127(.a(_w_8029),.q(_w_8030));
  bfr _b_3581(.a(_w_5483),.q(_w_5484));
  and_bb g1175(.a(N154_13),.b(N426_13),.q(n1175));
  spl2 g1473_s_0(.a(n1473),.q0(n1473_0),.q1(_w_12952));
  bfr _b_8206(.a(_w_10108),.q(_w_10109));
  bfr _b_4766(.a(_w_6668),.q(_w_6669));
  bfr _b_4797(.a(_w_6699),.q(_w_6700));
  bfr _b_4609(.a(_w_6511),.q(_w_6512));
  bfr _b_12445(.a(_w_14347),.q(_w_14348));
  and_bi g133(.a(n132_0),.b(n100_0),.q(n133));
  bfr _b_7117(.a(_w_9019),.q(_w_9020));
  bfr _b_8427(.a(_w_10329),.q(_w_10330));
  bfr _b_5378(.a(_w_7280),.q(_w_7281));
  bfr _b_9625(.a(_w_11527),.q(_w_11528));
  bfr _b_5846(.a(_w_7748),.q(_w_7749));
  bfr _b_7579(.a(_w_9481),.q(_w_9482));
  bfr _b_4665(.a(_w_6567),.q(_w_6568));
  bfr _b_6924(.a(_w_8826),.q(_w_8827));
  bfr _b_6906(.a(_w_8808),.q(n1636));
  bfr _b_11808(.a(_w_13710),.q(_w_13711));
  bfr _b_8157(.a(_w_10059),.q(_w_10060));
  and_bb g1179(.a(N188_11),.b(N392_15),.q(n1179));
  bfr _b_10975(.a(_w_12877),.q(_w_12878));
  bfr _b_4309(.a(_w_6211),.q(n664_1));
  spl2 g895_s_0(.a(n895),.q0(n895_0),.q1(n895_1));
  spl2 g1744_s_0(.a(n1744),.q0(n1744_0),.q1(n1744_1));
  bfr _b_7687(.a(_w_9589),.q(_w_9590));
  bfr _b_10321(.a(_w_12223),.q(_w_12224));
  bfr _b_4161(.a(_w_6063),.q(_w_6064));
  and_bb g1183(.a(N222_15),.b(N358_17),.q(_w_12956));
  and_bb g1470(.a(N239_11),.b(N392_18),.q(n1470));
  bfr _b_5875(.a(_w_7777),.q(_w_7778));
  or_bb g1188(.a(n1186_0),.b(n1187_0),.q(n1188));
  bfr _b_7553(.a(_w_9455),.q(_w_9456));
  and_bb g1189(.a(n1186_1),.b(n1187_1),.q(_w_12979));
  or_bb g1193(.a(n1191_0),.b(n1192),.q(n1193));
  or_bb g411(.a(n409_0),.b(n410),.q(n411));
  bfr _b_9457(.a(_w_11359),.q(_w_11360));
  spl2 g96_s_0(.a(n96),.q0(n96_0),.q1(n96_1));
  bfr _b_11576(.a(_w_13478),.q(_w_13479));
  bfr _b_6863(.a(_w_8765),.q(_w_8766));
  bfr _b_6131(.a(_w_8033),.q(_w_8034));
  bfr _b_8111(.a(_w_10013),.q(_w_10014));
  spl2 g1614_s_0(.a(n1614),.q0(n1614_0),.q1(n1614_1));
  and_bi g1197(.a(n1196_0),.b(n1183_0),.q(n1197));
  bfr _b_5651(.a(_w_7553),.q(_w_7554));
  bfr _b_12090(.a(_w_13992),.q(_w_13993));
  bfr _b_4155(.a(_w_6057),.q(_w_6058));
  bfr _b_3822(.a(_w_5724),.q(_w_5725));
  or_bb g1199(.a(n1197_0),.b(n1198),.q(n1199));
  bfr _b_12783(.a(_w_14685),.q(n1856));
  bfr _b_11838(.a(_w_13740),.q(_w_13741));
  or_bb g1205(.a(n1203_0),.b(n1204),.q(n1205));
  and_bb g571(.a(n533_1),.b(n569_1),.q(_w_12840));
  spl2 g1863_s_0(.a(n1863),.q0(n1863_0),.q1(n1863_1));
  spl2 g838_s_0(.a(n838),.q0(n838_0),.q1(n838_1));
  and_bb g1201(.a(n1182_1),.b(n1199_1),.q(_w_13001));
  bfr _b_14035(.a(_w_15937),.q(_w_15938));
  and_bi g1210(.a(n1179_1),.b(n1208_1),.q(_w_13002));
  spl2 g1852_s_0(.a(n1852),.q0(n1852_0),.q1(n1852_1));
  bfr _b_5488(.a(_w_7390),.q(_w_7391));
  bfr _b_12356(.a(_w_14258),.q(_w_14259));
  bfr _b_8467(.a(_w_10369),.q(_w_10370));
  or_bb g1212(.a(n1178_0),.b(n1211_0),.q(n1212));
  bfr _b_12541(.a(_w_14443),.q(_w_14444));
  bfr _b_10688(.a(_w_12590),.q(_w_12591));
  bfr _b_5971(.a(_w_7873),.q(N222_1));
  bfr _b_9963(.a(_w_11865),.q(_w_11866));
  bfr _b_6166(.a(_w_8068),.q(_w_8069));
  bfr _b_5921(.a(_w_7823),.q(_w_7824));
  bfr _b_3436(.a(_w_5338),.q(_w_5339));
  spl2 g997_s_0(.a(n997),.q0(n997_0),.q1(n997_1));
  bfr _b_5938(.a(_w_7840),.q(_w_7841));
  and_bi g1214(.a(n1212_0),.b(n1213),.q(n1214));
  bfr _b_3467(.a(_w_5369),.q(_w_5370));
  bfr _b_4798(.a(_w_6700),.q(_w_6701));
  spl2 g603_s_0(.a(n603),.q0(n603_0),.q1(n603_1));
  bfr _b_9862(.a(_w_11764),.q(_w_11765));
  or_bb g1445(.a(n1443_0),.b(n1444),.q(n1445));
  and_bi g1829(.a(n1827_0),.b(n1828),.q(n1829));
  or_bb g231(.a(n229_0),.b(n230),.q(_w_9759));
  bfr _b_7727(.a(_w_9629),.q(_w_9630));
  or_bb g1022(.a(n1021_0),.b(n943_0),.q(n1022));
  bfr _b_4486(.a(_w_6388),.q(_w_6389));
  bfr _b_5475(.a(_w_7377),.q(_w_7378));
  bfr _b_13117(.a(_w_15019),.q(n1340));
  spl2 g605_s_0(.a(n605),.q0(n605_0),.q1(n605_1));
  bfr _b_4508(.a(_w_6410),.q(_w_6411));
  bfr _b_12705(.a(_w_14607),.q(_w_14608));
  bfr _b_5803(.a(_w_7705),.q(_w_7706));
  spl2 g1851_s_0(.a(n1851),.q0(n1851_0),.q1(n1851_1));
  bfr _b_11515(.a(_w_13417),.q(_w_13418));
  bfr _b_4737(.a(_w_6639),.q(_w_6640));
  bfr _b_9410(.a(_w_11312),.q(_w_11313));
  or_bb g1217(.a(n1215_0),.b(n1216),.q(n1217));
  bfr _b_4115(.a(_w_6017),.q(_w_6018));
  bfr _b_6679(.a(_w_8581),.q(_w_8582));
  bfr _b_6601(.a(_w_8503),.q(_w_8504));
  bfr _b_8306(.a(_w_10208),.q(_w_10209));
  and_bb g840(.a(N171_9),.b(N358_14),.q(_w_9965));
  spl2 g624_s_0(.a(n624),.q0(n624_0),.q1(n624_1));
  and_bb g1219(.a(n1176_1),.b(n1217_1),.q(_w_13004));
  bfr _b_5375(.a(_w_7277),.q(_w_7278));
  bfr _b_9092(.a(_w_10994),.q(_w_10995));
  or_bb g323(.a(n321_0),.b(n322),.q(n323));
  bfr _b_12632(.a(_w_14534),.q(_w_14535));
  bfr _b_9375(.a(_w_11277),.q(_w_11278));
  and_bi g1533(.a(n1527_1),.b(n1530_1),.q(n1533));
  bfr _b_4169(.a(_w_6071),.q(_w_6072));
  and_bb g193(.a(N120_5),.b(N273_11),.q(n193));
  bfr _b_5913(.a(_w_7815),.q(_w_7816));
  spl2 g339_s_0(.a(n339),.q0(n339_0),.q1(n339_1));
  bfr _b_6821(.a(_w_8723),.q(_w_8724));
  bfr _b_12466(.a(_w_14368),.q(n682_1));
  and_bi g643(.a(n642_0),.b(n634_0),.q(n643));
  and_bi g1222(.a(n1175_1),.b(n1220_1),.q(_w_13005));
  or_bb g400(.a(n371_0),.b(n399_0),.q(n400));
  bfr _b_3596(.a(_w_5498),.q(_w_5499));
  spl2 g1431_s_0(.a(n1431),.q0(n1431_0),.q1(n1431_1));
  bfr _b_7137(.a(_w_9039),.q(_w_9040));
  bfr _b_4239(.a(_w_6141),.q(_w_6142));
  and_bb g1547(.a(N222_11),.b(N426_17),.q(n1547));
  spl2 g881_s_0(.a(n881),.q0(n881_0),.q1(_w_13006));
  and_bi g1232(.a(n1230_0),.b(n1231),.q(n1232));
  spl3L g542_s_0(.a(n542),.q0(n542_0),.q1(_w_14829),.q2(_w_14831));
  bfr _b_14052(.a(_w_15954),.q(_w_15955));
  bfr _b_7268(.a(_w_9170),.q(_w_9171));
  bfr _b_8163(.a(_w_10065),.q(_w_10066));
  bfr _b_8488(.a(_w_10390),.q(_w_10391));
  bfr _b_10067(.a(_w_11969),.q(_w_11970));
  and_bb g956(.a(N188_9),.b(N358_15),.q(_w_12347));
  or_bb g161(.a(n159_0),.b(n160),.q(n161));
  spl2 g983_s_0(.a(n983),.q0(n983_0),.q1(n983_1));
  bfr _b_3578(.a(_w_5480),.q(_w_5481));
  and_bi g788(.a(n722_1),.b(n786_1),.q(_w_13011));
  bfr _b_10839(.a(_w_12741),.q(_w_12742));
  and_bi g1245(.a(n1244_0),.b(n1167_0),.q(n1245));
  and_bb g665(.a(n627_1),.b(n663_1),.q(_w_8730));
  bfr _b_3978(.a(_w_5880),.q(_w_5881));
  and_bi g1246(.a(n1167_1),.b(n1244_1),.q(_w_13012));
  bfr _b_5676(.a(_w_7578),.q(_w_7579));
  and_bi g1714(.a(n1675_1),.b(n1712_1),.q(_w_13013));
  bfr _b_3870(.a(_w_5772),.q(_w_5773));
  bfr _b_12350(.a(_w_14252),.q(_w_14253));
  spl2 g1146_s_0(.a(n1146),.q0(n1146_0),.q1(n1146_1));
  spl2 g1174_s_0(.a(n1174),.q0(n1174_0),.q1(n1174_1));
  and_bb g1249(.a(n1166_1),.b(n1247_1),.q(_w_13014));
  and_bi g1529(.a(n1527_0),.b(n1528),.q(_w_13016));
  bfr _b_11775(.a(_w_13677),.q(_w_13678));
  spl2 g691_s_0(.a(n691),.q0(n691_0),.q1(n691_1));
  and_bi g1251(.a(n1250_0),.b(n1165_0),.q(n1251));
  bfr _b_12430(.a(_w_14332),.q(_w_14333));
  bfr _b_11574(.a(_w_13476),.q(_w_13477));
  and_bi g1252(.a(n1165_1),.b(n1250_1),.q(_w_13032));
  bfr _b_3430(.a(_w_5332),.q(_w_5333));
  bfr _b_7805(.a(_w_9707),.q(_w_9708));
  bfr _b_5949(.a(_w_7851),.q(_w_7852));
  spl2 g1177_s_0(.a(n1177),.q0(n1177_0),.q1(n1177_1));
  bfr _b_5411(.a(_w_7313),.q(_w_7314));
  bfr _b_11295(.a(_w_13197),.q(N103_11));
  or_bb g1254(.a(n1164_0),.b(n1253_0),.q(n1254));
  bfr _b_3534(.a(_w_5436),.q(_w_5437));
  bfr _b_6565(.a(_w_8467),.q(_w_8468));
  bfr _b_13356(.a(_w_15258),.q(_w_15259));
  spl2 g1570_s_0(.a(n1570),.q0(n1570_0),.q1(_w_13033));
  spl2 g1872_s_0(.a(n1872),.q0(n1872_0),.q1(n1872_1));
  spl2 g751_s_0(.a(n751),.q0(n751_0),.q1(n751_1));
  bfr _b_5386(.a(_w_7288),.q(_w_7289));
  and_bi g1257(.a(n1256_0),.b(n1163_0),.q(n1257));
  bfr _b_6246(.a(_w_8148),.q(_w_8149));
  bfr _b_4128(.a(_w_6030),.q(_w_6031));
  bfr _b_3977(.a(_w_5879),.q(_w_5880));
  bfr _b_3483(.a(_w_5385),.q(_w_5386));
  bfr _b_8172(.a(_w_10074),.q(_w_10075));
  spl2 g760_s_0(.a(n760),.q0(n760_0),.q1(_w_13044));
  spl2 g626_s_0(.a(n626),.q0(n626_0),.q1(n626_1));
  and_bb g1280(.a(N171_13),.b(N426_14),.q(n1280));
  bfr _b_4879(.a(_w_6781),.q(_w_6782));
  bfr _b_3943(.a(_w_5845),.q(_w_5846));
  and_bi g1267(.a(n1254_1),.b(n1257_1),.q(n1267));
  spl2 g1342_s_0(.a(n1342),.q0(n1342_0),.q1(n1342_1));
  bfr _b_6091(.a(_w_7993),.q(_w_7994));
  bfr _b_7597(.a(_w_9499),.q(_w_9500));
  bfr _b_8923(.a(_w_10825),.q(_w_10826));
  bfr _b_9281(.a(_w_11183),.q(_w_11184));
  bfr _b_3942(.a(_w_5844),.q(n929_1));
  and_bb g244(.a(N103_6),.b(N307_10),.q(_w_13049));
  or_bb g1875(.a(n1873_0),.b(n1874),.q(_w_13055));
  and_bi g447(.a(n400_1),.b(n403_1),.q(n447));
  and_bi g1269(.a(n1248_1),.b(n1251_1),.q(n1269));
  and_bb g1310(.a(n1283_1),.b(n1308_1),.q(_w_12913));
  bfr _b_7998(.a(_w_9900),.q(_w_9901));
  bfr _b_4000(.a(_w_5902),.q(_w_5903));
  bfr _b_3805(.a(_w_5707),.q(_w_5708));
  bfr _b_8502(.a(_w_10404),.q(_w_10405));
  and_bb g1270(.a(N511_9),.b(N86_18),.q(_w_13063));
  bfr _b_3639(.a(_w_5541),.q(_w_5542));
  and_bi g1273(.a(n1236_1),.b(n1239_1),.q(n1273));
  bfr _b_4582(.a(_w_6484),.q(_w_6485));
  bfr _b_9258(.a(_w_11160),.q(_w_11161));
  bfr _b_3898(.a(_w_5800),.q(_w_5801));
  and_bi g1592(.a(n1537_1),.b(n1590_1),.q(_w_13091));
  bfr _b_6890(.a(_w_8792),.q(n324_1));
  spl2 g1068_s_0(.a(n1068),.q0(n1068_0),.q1(n1068_1));
  bfr _b_4144(.a(_w_6046),.q(_w_6047));
  and_bi g494(.a(n444_1),.b(n492_1),.q(_w_10779));
  spl2 g1546_s_0(.a(n1546),.q0(n1546_0),.q1(n1546_1));
  bfr _b_7886(.a(_w_9788),.q(_w_9789));
  bfr _b_13650(.a(_w_15552),.q(_w_15553));
  spl2 g1407_s_0(.a(n1407),.q0(n1407_0),.q1(n1407_1));
  spl2 g1741_s_0(.a(n1741),.q0(n1741_0),.q1(_w_13092));
  bfr _b_5684(.a(_w_7586),.q(_w_7587));
  and_bi g1277(.a(n1224_1),.b(n1227_1),.q(n1277));
  and_bi g1279(.a(n1218_1),.b(n1221_1),.q(n1279));
  bfr _b_4234(.a(_w_6136),.q(_w_6137));
  bfr _b_4880(.a(_w_6782),.q(_w_6783));
  bfr _b_10043(.a(_w_11945),.q(_w_11946));
  bfr _b_11210(.a(_w_13112),.q(_w_13113));
  or_bb g1812(.a(n1778_0),.b(n1811_0),.q(_w_13101));
  bfr _b_10669(.a(_w_12571),.q(_w_12572));
  spl2 g525_s_0(.a(n525),.q0(n525_0),.q1(n525_1));
  bfr _b_7100(.a(_w_9002),.q(_w_9003));
  bfr _b_9430(.a(_w_11332),.q(_w_11333));
  bfr _b_14302(.a(_w_16204),.q(_w_16205));
  or_bb g273(.a(n271_0),.b(n272),.q(n273));
  bfr _b_5739(.a(_w_7641),.q(_w_7642));
  bfr _b_5842(.a(_w_7744),.q(_w_7745));
  bfr _b_9062(.a(_w_10964),.q(_w_10965));
  and_bb g1789(.a(n1786_1),.b(n1787_1),.q(_w_13149));
  and_bb g1286(.a(N222_14),.b(N375_17),.q(_w_13150));
  bfr _b_4478(.a(_w_6380),.q(_w_6381));
  and_bi g1596(.a(n1594_0),.b(n1595),.q(n1596));
  bfr _b_13194(.a(_w_15096),.q(n1309_1));
  and_bb g618(.a(N443_7),.b(N52_14),.q(_w_13166));
  and_bb g1289(.a(N256_16),.b(N341_19),.q(_w_13170));
  spl4L N103_s_2(.a(N103_1),.q0(N103_8),.q1(N103_9),.q2(N103_10),.q3(_w_13174));
  and_bi g1290(.a(n1188_1),.b(n1191_1),.q(n1290));
  bfr _b_7380(.a(_w_9282),.q(_w_9283));
  and_bb g1292(.a(n1289_1),.b(n1290_1),.q(_w_13199));
  spl2 g472_s_0(.a(n472),.q0(n472_0),.q1(_w_13200));
  bfr _b_10601(.a(_w_12503),.q(_w_12504));
  or_bb g1296(.a(n1294_0),.b(n1295),.q(n1296));
  bfr _b_14170(.a(_w_16072),.q(_w_16073));
  bfr _b_4094(.a(_w_5996),.q(_w_5997));
  and_bi g1091(.a(n1089_0),.b(n1090),.q(n1091));
  or_bb g893(.a(n833_0),.b(n892_0),.q(n893));
  bfr _b_5395(.a(_w_7297),.q(_w_7298));
  and_bi g1457(.a(n1428_1),.b(n1431_1),.q(n1457));
  bfr _b_4365(.a(_w_6267),.q(N120_11));
  bfr _b_9370(.a(_w_11272),.q(_w_11273));
  bfr _b_10806(.a(_w_12708),.q(N86_14));
  and_bi g1300(.a(n1299_0),.b(n1286_0),.q(n1300));
  bfr _b_12923(.a(_w_14825),.q(_w_14826));
  bfr _b_8438(.a(_w_10340),.q(_w_10341));
  and_bi g1306(.a(n1305_0),.b(n1284_0),.q(n1306));
  bfr _b_8844(.a(_w_10746),.q(_w_10747));
  bfr _b_5606(.a(_w_7508),.q(_w_7509));
  bfr _b_10228(.a(_w_12130),.q(_w_12131));
  or_bb g1314(.a(n1312_0),.b(n1313),.q(n1314));
  bfr _b_5743(.a(_w_7645),.q(_w_7646));
  bfr _b_5332(.a(_w_7234),.q(N545));
  bfr _b_9113(.a(_w_11015),.q(n110));
  spl2 g444_s_0(.a(n444),.q0(n444_0),.q1(n444_1));
  spl2 g368_s_0(.a(n368),.q0(n368_0),.q1(n368_1));
  spl2 g1806_s_0(.a(n1806),.q0(n1806_0),.q1(_w_6296));
  and_bi g959(.a(n857_1),.b(n860_1),.q(n959));
  bfr _b_6111(.a(_w_8013),.q(_w_8014));
  spl2 g1540_s_0(.a(n1540),.q0(n1540_0),.q1(n1540_1));
  and_bi g1777(.a(n1771_1),.b(n1774_1),.q(n1777));
  spl2 g1248_s_0(.a(n1248),.q0(n1248_0),.q1(_w_15105));
  bfr _b_4907(.a(_w_6809),.q(_w_6810));
  bfr _b_3857(.a(_w_5759),.q(_w_5760));
  and_bi g1319(.a(n1280_1),.b(n1317_1),.q(_w_13346));
  spl4L N256_s_2(.a(N256_1),.q0(_w_13347),.q1(N256_9),.q2(N256_10),.q3(N256_11));
  or_bb g1320(.a(n1318_0),.b(n1319),.q(n1320));
  spl2 g268_s_0(.a(n268),.q0(n268_0),.q1(_w_13367));
  and_bb g828(.a(N460_8),.b(N69_15),.q(_w_8927));
  and_bi g212(.a(n186_1),.b(n210_1),.q(_w_13371));
  spl2 g1107_s_0(.a(n1107),.q0(n1107_0),.q1(_w_15007));
  and_bi g731(.a(n652_1),.b(n655_1),.q(n731));
  bfr _b_9489(.a(_w_11391),.q(_w_11392));
  bfr _b_4762(.a(_w_6664),.q(_w_6665));
  or_bb g557(.a(n555_0),.b(n556),.q(n557));
  or_bb g1321(.a(n1279_0),.b(n1320_0),.q(n1321));
  bfr _b_10047(.a(_w_11949),.q(_w_11950));
  spl2 g536_s_0(.a(n536),.q0(n536_0),.q1(n536_1));
  bfr _b_7174(.a(_w_9076),.q(_w_9077));
  bfr _b_7209(.a(_w_9111),.q(_w_9112));
  bfr _b_8225(.a(_w_10127),.q(_w_10128));
  spl2 g481_s_0(.a(n481),.q0(n481_0),.q1(n481_1));
  or_bb g1845(.a(n1819_0),.b(n1844_0),.q(_w_14573));
  and_bi g937(.a(n923_1),.b(n926_1),.q(n937));
  and_bi g1323(.a(n1321_0),.b(n1322),.q(n1323));
  bfr _b_8091(.a(_w_9993),.q(_w_9994));
  bfr _b_9921(.a(_w_11823),.q(_w_11824));
  and_bi g717(.a(n694_1),.b(n697_1),.q(n717));
  bfr _b_7138(.a(_w_9040),.q(N188_2));
  and_bi g853(.a(n852_0),.b(n847),.q(n853));
  spl2 g1781_s_0(.a(n1781),.q0(n1781_0),.q1(n1781_1));
  and_bi g122(.a(n104_1),.b(n120_1),.q(_w_11024));
  spl2 g1764_s_0(.a(n1764),.q0(n1764_0),.q1(n1764_1));
  bfr _b_5749(.a(_w_7651),.q(_w_7652));
  and_bi g1325(.a(n1278_1),.b(n1323_1),.q(_w_13372));
  spl4L N443_s_2(.a(N443_1),.q0(N443_8),.q1(N443_9),.q2(N443_10),.q3(N443_11));
  spl2 g1588_s_0(.a(n1588),.q0(n1588_0),.q1(_w_13373));
  and_bi g1370(.a(n1333_1),.b(n1336_1),.q(n1370));
  and_bi g1329(.a(n1327_0),.b(n1328),.q(n1329));
  spl2 g898_s_0(.a(n898),.q0(n898_0),.q1(n898_1));
  and_bi g1784(.a(n1747_1),.b(n1750_1),.q(n1784));
  and_bi g1335(.a(n1333_0),.b(n1334),.q(n1335));
  bfr _b_4066(.a(_w_5968),.q(_w_5969));
  bfr _b_6921(.a(_w_8823),.q(_w_8824));
  bfr _b_7488(.a(_w_9390),.q(_w_9391));
  spl2 g1227_s_0(.a(n1227),.q0(n1227_0),.q1(n1227_1));
  spl4L N86_s_0(.a(_w_16288),.q0(N86_0),.q1(_w_7295),.q2(_w_7319),.q3(_w_7375));
  or_bb g1339(.a(n1273_0),.b(n1338_0),.q(n1339));
  spl2 g484_s_0(.a(n484),.q0(n484_0),.q1(_w_13426));
  spl4L N307_s_1(.a(N307_0),.q0(N307_4),.q1(N307_5),.q2(N307_6),.q3(N307_7));
  or_bb g1532(.a(n1530_0),.b(n1531),.q(_w_12241));
  bfr _b_9621(.a(_w_11523),.q(_w_11524));
  bfr _b_4960(.a(_w_6862),.q(_w_6863));
  and_bi g1341(.a(n1339_0),.b(n1340),.q(n1341));
  bfr _b_8749(.a(_w_10651),.q(_w_10652));
  bfr _b_10871(.a(_w_12773),.q(_w_12774));
  and_bi g1348(.a(n1347_0),.b(n1270_0),.q(n1348));
  bfr _b_12306(.a(_w_14208),.q(_w_14209));
  spl2 g1461_s_0(.a(n1461),.q0(n1461_0),.q1(n1461_1));
  and_bi g984(.a(n956_1),.b(n982_1),.q(_w_13433));
  spl2 g558_s_0(.a(n558),.q0(n558_0),.q1(_w_9578));
  or_bb g1350(.a(n1348_0),.b(n1349),.q(n1350));
  bfr _b_3480(.a(_w_5382),.q(_w_5383));
  bfr _b_3788(.a(_w_5690),.q(_w_5691));
  bfr _b_4448(.a(_w_6350),.q(_w_6351));
  bfr _b_5870(.a(_w_7772),.q(_w_7773));
  bfr _b_5910(.a(_w_7812),.q(_w_7813));
  or_bb g1351(.a(n1269_0),.b(n1350_0),.q(n1351));
  and_bb g1352(.a(n1269_1),.b(n1350_1),.q(_w_13434));
  and_bi g1353(.a(n1351_0),.b(n1352),.q(n1353));
  and_bi g1354(.a(n1353_0),.b(n1268_0),.q(n1354));
  bfr _b_10614(.a(_w_12516),.q(n497));
  bfr _b_9154(.a(_w_11056),.q(_w_11057));
  spl4L N375_s_2(.a(N375_1),.q0(N375_8),.q1(N375_9),.q2(N375_10),.q3(N375_11));
  or_bb g808(.a(n715_0),.b(n807_0),.q(n808));
  bfr _b_9863(.a(_w_11765),.q(_w_11766));
  bfr _b_4525(.a(_w_6427),.q(N137_6));
  and_bi g1843(.a(n1820_1),.b(n1841_1),.q(_w_13437));
  bfr _b_4008(.a(_w_5910),.q(N239_6));
  and_bb g1358(.a(n1267_1),.b(n1356_1),.q(_w_13438));
  and_bi g1359(.a(n1357_0),.b(n1358),.q(n1359));
  bfr _b_12644(.a(_w_14546),.q(_w_14547));
  bfr _b_9532(.a(_w_11434),.q(_w_11435));
  bfr _b_3434(.a(_w_5336),.q(_w_5337));
  and_bi g1043(.a(n1042_0),.b(n936_0),.q(n1043));
  or_bb g1362(.a(n1360_0),.b(n1361),.q(_w_13448));
  bfr _b_8998(.a(_w_10900),.q(_w_10901));
  bfr _b_3618(.a(_w_5520),.q(_w_5521));
  bfr _b_8372(.a(_w_10274),.q(_w_10275));
  bfr _b_10048(.a(_w_11950),.q(_w_11951));
  bfr _b_10953(.a(_w_12855),.q(n1150));
  bfr _b_9669(.a(_w_11571),.q(_w_11572));
  bfr _b_7868(.a(_w_9770),.q(_w_9771));
  and_bi g1891(.a(n1876_1),.b(n1889_1),.q(_w_13512));
  bfr _b_8000(.a(_w_9902),.q(_w_9903));
  bfr _b_9885(.a(_w_11787),.q(_w_11788));
  bfr _b_4772(.a(_w_6674),.q(_w_6675));
  and_bi g1368(.a(n1339_1),.b(n1342_1),.q(n1368));
  bfr _b_9348(.a(_w_11250),.q(_w_11251));
  and_bb g1126(.a(n1059_1),.b(n1124_1),.q(_w_10821));
  or_bb g353(.a(n351_0),.b(n352),.q(n353));
  bfr _b_9024(.a(_w_10926),.q(_w_10927));
  bfr _b_9840(.a(_w_11742),.q(_w_11743));
  and_bb g1369(.a(N120_17),.b(N494_11),.q(_w_13513));
  bfr _b_13581(.a(_w_15483),.q(_w_15484));
  bfr _b_4413(.a(_w_6315),.q(_w_6316));
  bfr _b_6046(.a(_w_7948),.q(_w_7949));
  bfr _b_3894(.a(_w_5796),.q(_w_5797));
  and_bi g907(.a(n905_0),.b(n906),.q(n907));
  bfr _b_8289(.a(_w_10191),.q(_w_10192));
  spl2 g412_s_0(.a(n412),.q0(n412_0),.q1(_w_13521));
  bfr _b_11792(.a(_w_13694),.q(_w_13695));
  and_bi g432(.a(n430_0),.b(n431),.q(n432));
  spl2 g1787_s_0(.a(n1787),.q0(n1787_0),.q1(n1787_1));
  bfr _b_13892(.a(_w_15794),.q(_w_15795));
  spl2 g645_s_0(.a(n645),.q0(n645_0),.q1(n645_1));
  spl2 g1547_s_0(.a(n1547),.q0(n1547_0),.q1(n1547_1));
  bfr _b_4754(.a(_w_6656),.q(_w_6657));
  and_bi g704(.a(n614_1),.b(n702_1),.q(_w_13038));
  bfr _b_7168(.a(_w_9070),.q(_w_9071));
  spl2 g560_s_0(.a(n560),.q0(n560_0),.q1(n560_1));
  bfr _b_8828(.a(_w_10730),.q(_w_10731));
  and_bb g1373(.a(N154_15),.b(N460_13),.q(_w_13525));
  spl2 g646_s_0(.a(n646),.q0(n646_0),.q1(_w_11602));
  bfr _b_6674(.a(_w_8576),.q(_w_8577));
  and_bi g1374(.a(n1321_1),.b(n1324_1),.q(n1374));
  bfr _b_6728(.a(_w_8630),.q(_w_8631));
  bfr _b_13775(.a(_w_15677),.q(_w_15678));
  spl3L g737_s_0(.a(n737),.q0(n737_0),.q1(_w_13537),.q2(n737_2));
  and_bb g1377(.a(N188_13),.b(N426_15),.q(n1377));
  and_bi g1380(.a(n1303_1),.b(n1306_1),.q(n1380));
  bfr _b_4136(.a(_w_6038),.q(_w_6039));
  bfr _b_8788(.a(_w_10690),.q(_w_10691));
  bfr _b_5033(.a(_w_6935),.q(_w_6936));
  bfr _b_9420(.a(_w_11322),.q(_w_11323));
  or_bb g1858(.a(n1856_0),.b(n1857_0),.q(n1858));
  and_bb g1381(.a(N222_4),.b(N392_17),.q(n1381));
  bfr _b_4906(.a(_w_6808),.q(_w_6809));
  bfr _b_7509(.a(_w_9411),.q(_w_9412));
  spl2 g1163_s_0(.a(n1163),.q0(n1163_0),.q1(n1163_1));
  bfr _b_10944(.a(_w_12846),.q(_w_12847));
  bfr _b_4146(.a(_w_6048),.q(_w_6049));
  spl2 g1499_s_0(.a(n1499),.q0(n1499_0),.q1(n1499_1));
  or_bb g1386(.a(n1384_0),.b(n1385_0),.q(n1386));
  and_bi g1388(.a(n1386_0),.b(n1387),.q(n1388));
  bfr _b_7232(.a(_w_9134),.q(n1225));
  bfr _b_3852(.a(_w_5754),.q(_w_5755));
  bfr _b_4649(.a(_w_6551),.q(_w_6552));
  spl2 g1400_s_0(.a(n1400),.q0(n1400_0),.q1(n1400_1));
  bfr _b_7673(.a(_w_9575),.q(_w_9576));
  and_bi g1809(.a(n1808_0),.b(n1779_0),.q(n1809));
  bfr _b_12104(.a(_w_14006),.q(_w_14007));
  bfr _b_10504(.a(_w_12406),.q(_w_12407));
  bfr _b_5088(.a(_w_6990),.q(_w_6991));
  bfr _b_5716(.a(_w_7618),.q(_w_7619));
  bfr _b_5399(.a(_w_7301),.q(_w_7302));
  spl2 g522_s_0(.a(n522),.q0(n522_0),.q1(n522_1));
  bfr _b_8552(.a(_w_10454),.q(_w_10455));
  spl2 g694_s_0(.a(n694),.q0(n694_0),.q1(_w_6192));
  bfr _b_5075(.a(_w_6977),.q(_w_6978));
  bfr _b_4125(.a(_w_6027),.q(_w_6028));
  bfr _b_7054(.a(_w_8956),.q(_w_8957));
  spl2 g1200_s_0(.a(n1200),.q0(n1200_0),.q1(_w_13566));
  and_bb g1393(.a(n1382_1),.b(n1391_1),.q(_w_13570));
  or_bb g1397(.a(n1395_0),.b(n1396),.q(n1397));
  bfr _b_7753(.a(_w_9655),.q(_w_9656));
  bfr _b_11201(.a(_w_13103),.q(_w_13104));
  bfr _b_8539(.a(_w_10441),.q(n918));
  and_bi g243(.a(n196_1),.b(n199_1),.q(n243));
  bfr _b_3428(.a(_w_5330),.q(_w_5331));
  and_bi g1701(.a(n1700_0),.b(n1679_0),.q(n1701));
  bfr _b_6400(.a(_w_8302),.q(_w_8303));
  bfr _b_10825(.a(_w_12727),.q(_w_12728));
  or_bb g1409(.a(n1407_0),.b(n1408),.q(n1409));
  bfr _b_12927(.a(_w_14829),.q(_w_14830));
  and_bb g577(.a(n531_1),.b(n575_1),.q(_w_13578));
  bfr _b_6062(.a(_w_7964),.q(_w_7965));
  and_bi g1412(.a(n1410_0),.b(n1411),.q(n1412));
  spl2 g1112_s_0(.a(n1112),.q0(n1112_0),.q1(n1112_1));
  or_bb g1416(.a(n1374_0),.b(n1415_0),.q(n1416));
  bfr _b_14018(.a(_w_15920),.q(_w_15921));
  spl2 g1299_s_0(.a(n1299),.q0(n1299_0),.q1(n1299_1));
  spl4L N358_s_4(.a(N358_3),.q0(N358_16),.q1(N358_17),.q2(N358_18),.q3(N358_19));
  bfr _b_9156(.a(_w_11058),.q(_w_11059));
  and_bi g1418(.a(n1416_0),.b(n1417),.q(n1418));
  bfr _b_11140(.a(_w_13042),.q(_w_13043));
  and_bi g1420(.a(n1373_1),.b(n1418_1),.q(_w_13581));
  and_bi g121(.a(n120_0),.b(n104_0),.q(n121));
  bfr _b_4312(.a(_w_6214),.q(_w_6215));
  or_bb g1421(.a(n1419_0),.b(n1420),.q(n1421));
  or_bb g82(.a(n56_1),.b(n81_0),.q(n82));
  bfr _b_13387(.a(_w_15289),.q(_w_15290));
  bfr _b_7186(.a(_w_9088),.q(_w_9089));
  bfr _b_8530(.a(_w_10432),.q(_w_10433));
  and_bb g1693(.a(n1682_1),.b(n1691_1),.q(_w_14114));
  bfr _b_9626(.a(_w_11528),.q(_w_11529));
  bfr _b_10515(.a(_w_12417),.q(_w_12418));
  bfr _b_7903(.a(_w_9805),.q(_w_9806));
  spl2 g1710_s_0(.a(n1710),.q0(n1710_0),.q1(_w_9253));
  bfr _b_4052(.a(_w_5954),.q(_w_5955));
  and_bi g1755(.a(n1753_0),.b(n1754),.q(n1755));
  spl2 g68_s_0(.a(n68),.q0(n68_0),.q1(n68_1));
  and_bi g1424(.a(n1422_0),.b(n1423),.q(n1424));
  and_bi g270(.a(n268_0),.b(n269),.q(n270));
  bfr _b_3551(.a(_w_5453),.q(_w_5454));
  bfr _b_13768(.a(N409),.q(_w_15671));
  bfr _b_6321(.a(_w_8223),.q(n1077_1));
  or_bb g1427(.a(n1425_0),.b(n1426),.q(n1427));
  bfr _b_9013(.a(_w_10915),.q(_w_10916));
  or_bb g563(.a(n561_0),.b(n562),.q(n563));
  bfr _b_8780(.a(_w_10682),.q(_w_10683));
  bfr _b_13427(.a(_w_15329),.q(_w_15330));
  and_bb g138(.a(N18_9),.b(N358_5),.q(_w_11109));
  and_bi g1176(.a(n1107_1),.b(n1110_1),.q(n1176));
  bfr _b_13179(.a(_w_15081),.q(_w_15082));
  or_bb g1148(.a(n1146_0),.b(n1147),.q(n1148));
  bfr _b_9162(.a(_w_11064),.q(_w_11065));
  or_bb g1428(.a(n1370_0),.b(n1427_0),.q(n1428));
  and_bi g1430(.a(n1428_0),.b(n1429),.q(n1430));
  bfr _b_12477(.a(_w_14379),.q(_w_14380));
  spl2 g466_s_0(.a(n466),.q0(n466_0),.q1(_w_13746));
  bfr _b_9355(.a(_w_11257),.q(_w_11258));
  bfr _b_3413(.a(_w_5315),.q(_w_5316));
  bfr _b_5879(.a(_w_7781),.q(_w_7782));
  bfr _b_4207(.a(_w_6109),.q(_w_6110));
  and_bi g1437(.a(n1436_0),.b(n1367_0),.q(n1437));
  bfr _b_4351(.a(_w_6253),.q(_w_6254));
  spl2 g418_s_0(.a(n418),.q0(n418_0),.q1(_w_13752));
  bfr _b_4547(.a(_w_6449),.q(N154_14));
  bfr _b_5862(.a(_w_7764),.q(_w_7765));
  bfr _b_6665(.a(_w_8567),.q(_w_8568));
  bfr _b_12179(.a(_w_14081),.q(_w_14082));
  bfr _b_8913(.a(_w_10815),.q(_w_10816));
  bfr _b_13023(.a(_w_14925),.q(_w_14926));
  and_bi g1448(.a(n1446_0),.b(n1447),.q(_w_13757));
  bfr _b_6865(.a(_w_8767),.q(_w_8768));
  bfr _b_8662(.a(_w_10564),.q(n1089_1));
  bfr _b_14338(.a(_w_16240),.q(_w_16241));
  bfr _b_10814(.a(_w_12716),.q(_w_12717));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(n140_1));
  spl2 g947_s_0(.a(n947),.q0(n947_0),.q1(n947_1));
  bfr _b_12438(.a(_w_14340),.q(n1775));
  spl4L N103_s_3(.a(N103_2),.q0(N103_12),.q1(_w_13770),.q2(_w_13778),.q3(_w_13790));
  or_bb g1697(.a(n1695_0),.b(n1696),.q(n1697));
  and_bb g1454(.a(N103_19),.b(N528_10),.q(_w_13802));
  spl2 g362_s_0(.a(n362),.q0(n362_0),.q1(n362_1));
  bfr _b_7284(.a(_w_9186),.q(_w_9187));
  bfr _b_9404(.a(_w_11306),.q(_w_11307));
  and_bi g1455(.a(n1434_1),.b(n1437_1),.q(n1455));
  bfr _b_4729(.a(_w_6631),.q(_w_6632));
  and_bi g295(.a(n280_1),.b(n283_1),.q(n295));
  spl2 g1284_s_0(.a(n1284),.q0(n1284_0),.q1(n1284_1));
  bfr _b_6049(.a(_w_7951),.q(N188_11));
  and_bb g1316(.a(n1281_1),.b(n1314_1),.q(_w_12076));
  and_bb g1458(.a(N137_17),.b(N494_12),.q(_w_13826));
  spl2 g1273_s_0(.a(n1273),.q0(n1273_0),.q1(n1273_1));
  spl2 g1713_s_0(.a(n1713),.q0(n1713_0),.q1(n1713_1));
  bfr _b_5595(.a(_w_7497),.q(_w_7498));
  spl2 g1718_s_0(.a(n1718),.q0(n1718_0),.q1(n1718_1));
  and_bb g553(.a(n539_1),.b(n551_1),.q(_w_10880));
  and_bb g1781(.a(N205_18),.b(N511_16),.q(_w_13834));
  bfr _b_9055(.a(_w_10957),.q(_w_10958));
  and_bi g1459(.a(n1422_1),.b(n1425_1),.q(n1459));
  bfr _b_13608(.a(_w_15510),.q(_w_15511));
  bfr _b_9591(.a(_w_11493),.q(_w_11494));
  spl2 g537_s_0(.a(n537),.q0(n537_0),.q1(n537_1));
  spl2 N256_s_5(.a(N256_19),.q0(N256_20),.q1(N256_21));
  bfr _b_10034(.a(_w_11936),.q(_w_11937));
  bfr _b_7010(.a(_w_8912),.q(_w_8913));
  bfr _b_12625(.a(_w_14527),.q(_w_14528));
  or_bb g220(.a(n183_0),.b(n219_0),.q(n220));
  spl2 g1893_s_0(.a(n1893),.q0(n1893_0),.q1(n1893_1));
  bfr _b_4727(.a(_w_6629),.q(_w_6630));
  bfr _b_4779(.a(_w_6681),.q(_w_6682));
  bfr _b_10835(.a(_w_12737),.q(_w_12738));
  spl2 g451_s_0(.a(n451),.q0(n451_0),.q1(n451_1));
  bfr _b_9471(.a(_w_11373),.q(_w_11374));
  bfr _b_7720(.a(_w_9622),.q(n592));
  and_bi g1463(.a(n1410_1),.b(n1413_1),.q(n1463));
  bfr _b_3720(.a(_w_5622),.q(_w_5623));
  bfr _b_7052(.a(_w_8954),.q(n1230_1));
  bfr _b_13834(.a(_w_15736),.q(_w_15737));
  bfr _b_10031(.a(_w_11933),.q(_w_11934));
  spl2 g1072_s_0(.a(n1072),.q0(n1072_0),.q1(n1072_1));
  bfr _b_4666(.a(_w_6568),.q(_w_6569));
  bfr _b_3815(.a(_w_5717),.q(_w_5718));
  bfr _b_6210(.a(_w_8112),.q(_w_8113));
  bfr _b_13918(.a(_w_15820),.q(_w_15821));
  bfr _b_9597(.a(_w_11499),.q(_w_11500));
  and_bi g770(.a(n728_1),.b(n768_1),.q(_w_9131));
  and_bi g781(.a(n780_0),.b(n724_0),.q(n781));
  and_bi g1597(.a(n1596_0),.b(n1535_0),.q(n1597));
  bfr _b_8344(.a(_w_10246),.q(_w_10247));
  bfr _b_8350(.a(_w_10252),.q(_w_10253));
  bfr _b_3485(.a(_w_5387),.q(_w_5388));
  bfr _b_4040(.a(_w_5942),.q(_w_5943));
  bfr _b_4222(.a(_w_6124),.q(N171_15));
  and_bi g1472(.a(n1386_1),.b(n1389_1),.q(n1472));
  bfr _b_3881(.a(_w_5783),.q(_w_5784));
  spl2 g1561_s_0(.a(n1561),.q0(n1561_0),.q1(n1561_1));
  spl2 g1898_s_0(.a(n1898),.q0(n1898_0),.q1(n1898_1));
  bfr _b_11505(.a(_w_13407),.q(_w_13408));
  bfr _b_5206(.a(_w_7108),.q(_w_7109));
  and_bi g224(.a(n182_1),.b(n222_1),.q(_w_13854));
  bfr _b_11581(.a(_w_13483),.q(_w_13484));
  and_bi g988(.a(n986_0),.b(n987),.q(n988));
  bfr _b_9687(.a(_w_11589),.q(_w_11590));
  and_bb g1480(.a(n1469_1),.b(n1478_1),.q(_w_13855));
  bfr _b_9629(.a(_w_11531),.q(_w_11532));
  bfr _b_13283(.a(_w_15185),.q(_w_15186));
  spl2 g1314_s_0(.a(n1314),.q0(n1314_0),.q1(n1314_1));
  and_bi g1202(.a(n1200_0),.b(n1201),.q(n1202));
  and_bi g1637(.a(n1635_0),.b(n1636),.q(n1637));
  bfr _b_8171(.a(_w_10073),.q(_w_10074));
  or_bb g1485(.a(n1467_0),.b(n1484_0),.q(n1485));
  spl2 g1455_s_0(.a(n1455),.q0(n1455_0),.q1(n1455_1));
  spl2 g155_s_0(.a(n155),.q0(n155_0),.q1(n155_1));
  or_bb g1040(.a(n1039_0),.b(n937_0),.q(n1040));
  or_bb g87(.a(n85_0),.b(n86),.q(n87));
  bfr _b_9483(.a(_w_11385),.q(_w_11386));
  bfr _b_13821(.a(_w_15723),.q(_w_15724));
  spl2 g1208_s_0(.a(n1208),.q0(n1208_0),.q1(n1208_1));
  spl2 g1616_s_0(.a(n1616),.q0(n1616_0),.q1(n1616_1));
  bfr _b_8607(.a(_w_10509),.q(_w_10510));
  and_bi g602(.a(n600_0),.b(n601),.q(n602));
  bfr _b_10063(.a(_w_11965),.q(_w_11966));
  or_bb g1491(.a(n1465_0),.b(n1490_0),.q(n1491));
  bfr _b_6121(.a(_w_8023),.q(N205_7));
  bfr _b_9241(.a(_w_11143),.q(_w_11144));
  bfr _b_9353(.a(_w_11255),.q(_w_11256));
  bfr _b_3746(.a(_w_5648),.q(_w_5649));
  spl2 g1457_s_0(.a(n1457),.q0(n1457_0),.q1(n1457_1));
  and_bi g1494(.a(n1493_0),.b(n1464_0),.q(n1494));
  and_bb g1498(.a(n1463_1),.b(n1496_1),.q(_w_13862));
  spl4L N239_s_4(.a(N239_3),.q0(N239_16),.q1(N239_17),.q2(N239_18),.q3(N239_19));
  and_bi g1499(.a(n1497_0),.b(n1498),.q(n1499));
  bfr _b_10941(.a(_w_12843),.q(_w_12844));
  bfr _b_5390(.a(_w_7292),.q(_w_7293));
  or_bb g1502(.a(n1500_0),.b(n1501),.q(n1502));
  bfr _b_13322(.a(_w_15224),.q(_w_15225));
  and_bb g1365(.a(N528_9),.b(N86_19),.q(_w_9892));
  and_bi g1506(.a(n1505_0),.b(n1460_0),.q(n1506));
  bfr _b_6598(.a(_w_8500),.q(_w_8501));
  and_bb g1673(.a(N154_19),.b(N528_13),.q(_w_9660));
  or_bb g207(.a(n205_0),.b(n206),.q(n207));
  spl2 g301_s_0(.a(n301),.q0(n301_0),.q1(n301_1));
  spl4L N375_s_3(.a(N375_2),.q0(N375_12),.q1(N375_13),.q2(N375_14),.q3(N375_15));
  and_bi g1507(.a(n1460_1),.b(n1505_1),.q(_w_13863));
  bfr _b_5363(.a(_w_7265),.q(_w_7266));
  or_bb g1509(.a(n1459_0),.b(n1508_0),.q(n1509));
  bfr _b_3738(.a(_w_5640),.q(_w_5641));
  spl4L N307_s_4(.a(N307_3),.q0(N307_16),.q1(N307_17),.q2(N307_18),.q3(N307_19));
  bfr _b_7069(.a(_w_8971),.q(_w_8972));
  spl2 g1524_s_0(.a(n1524),.q0(n1524_0),.q1(n1524_1));
  bfr _b_12841(.a(_w_14743),.q(_w_14744));
  bfr _b_11963(.a(_w_13865),.q(_w_13866));
  bfr _b_7177(.a(_w_9079),.q(_w_9080));
  bfr _b_6072(.a(_w_7974),.q(_w_7975));
  bfr _b_12274(.a(_w_14176),.q(n1853));
  bfr _b_4904(.a(_w_6806),.q(_w_6807));
  bfr _b_10271(.a(_w_12173),.q(_w_12174));
  bfr _b_9994(.a(_w_11896),.q(_w_11897));
  and_bi g1719(.a(n1718_0),.b(n1673_0),.q(n1719));
  bfr _b_4189(.a(_w_6091),.q(_w_6092));
  and_bi g1511(.a(n1509_0),.b(n1510),.q(n1511));
  or_bb g1758(.a(n1756_0),.b(n1757),.q(n1758));
  and_bi g1512(.a(n1511_0),.b(n1458_0),.q(n1512));
  bfr _b_13063(.a(_w_14965),.q(_w_14966));
  bfr _b_11008(.a(_w_12910),.q(_w_12911));
  bfr _b_6129(.a(_w_8031),.q(n1022_1));
  bfr _b_4979(.a(_w_6881),.q(n1653_1));
  bfr _b_14126(.a(_w_16028),.q(_w_16029));
  bfr _b_4404(.a(_w_6306),.q(_w_6307));
  spl2 g1074_s_0(.a(n1074),.q0(n1074_0),.q1(n1074_1));
  bfr _b_12556(.a(_w_14458),.q(_w_14459));
  and_bi g1342(.a(n1341_0),.b(n1272_0),.q(n1342));
  bfr _b_8896(.a(_w_10798),.q(_w_10799));
  bfr _b_13458(.a(_w_15360),.q(_w_15361));
  spl2 g1001_s_0(.a(n1001),.q0(n1001_0),.q1(n1001_1));
  or_bb g405(.a(n403_0),.b(n404),.q(n405));
  spl4L N69_s_4(.a(N69_3),.q0(N69_16),.q1(N69_17),.q2(N69_18),.q3(N69_19));
  spl2 g189_s_0(.a(n189),.q0(n189_0),.q1(n189_1));
  and_bi g1378(.a(n1309_1),.b(n1312_1),.q(n1378));
  bfr _b_11184(.a(_w_13086),.q(n1272));
  bfr _b_7021(.a(_w_8923),.q(_w_8924));
  bfr _b_10438(.a(_w_12340),.q(_w_12341));
  bfr _b_8792(.a(_w_10694),.q(_w_10695));
  bfr _b_7627(.a(_w_9529),.q(_w_9530));
  and_bb g1522(.a(n1455_1),.b(n1520_1),.q(_w_13873));
  bfr _b_6795(.a(_w_8697),.q(_w_8698));
  bfr _b_4188(.a(_w_6090),.q(_w_6091));
  bfr _b_3603(.a(_w_5505),.q(_w_5506));
  bfr _b_3662(.a(_w_5564),.q(n1040_1));
  bfr _b_5116(.a(_w_7018),.q(_w_7019));
  bfr _b_13547(.a(_w_15449),.q(_w_15450));
  bfr _b_13315(.a(_w_15217),.q(_w_15218));
  bfr _b_11094(.a(_w_12996),.q(_w_12997));
  spl2 g120_s_0(.a(n120),.q0(n120_0),.q1(n120_1));
  bfr _b_4935(.a(_w_6837),.q(_w_6838));
  bfr _b_3715(.a(_w_5617),.q(_w_5618));
  spl2 g946_s_0(.a(n946),.q0(n946_0),.q1(n946_1));
  bfr _b_4524(.a(_w_6426),.q(_w_6427));
  and_bi g1695(.a(n1694_0),.b(n1681_0),.q(n1695));
  bfr _b_5276(.a(_w_7178),.q(_w_7179));
  or_bb g1527(.a(n1453_0),.b(n1526_0),.q(n1527));
  bfr _b_6364(.a(_w_8266),.q(_w_8267));
  and_bb g1528(.a(n1453_1),.b(n1526_1),.q(_w_13886));
  bfr _b_3711(.a(_w_5613),.q(_w_5614));
  or_bb g148(.a(n107_1),.b(n147_0),.q(_w_11599));
  bfr _b_8264(.a(_w_10166),.q(_w_10167));
  bfr _b_9592(.a(_w_11494),.q(_w_11495));
  bfr _b_5562(.a(_w_7464),.q(_w_7465));
  bfr _b_14087(.a(_w_15989),.q(_w_15990));
  bfr _b_11363(.a(_w_13265),.q(_w_13266));
  and_bi g398(.a(n372_1),.b(n396_1),.q(_w_13901));
  and_bi g1536(.a(n1515_1),.b(n1518_1),.q(n1536));
  bfr _b_11202(.a(_w_13104),.q(_w_13105));
  bfr _b_6268(.a(_w_8170),.q(_w_8171));
  spl2 g1712_s_0(.a(n1712),.q0(n1712_0),.q1(n1712_1));
  bfr _b_3988(.a(_w_5890),.q(_w_5891));
  and_bi g1014(.a(n946_1),.b(n1012_1),.q(_w_13906));
  bfr _b_8987(.a(_w_10889),.q(_w_10890));
  and_bi g617(.a(n594_1),.b(n597_1),.q(n617));
  or_bb g1659(.a(n1609_0),.b(n1658_0),.q(n1659));
  spl2 g357_s_0(.a(n357),.q0(n357_0),.q1(n357_1));
  bfr _b_5898(.a(_w_7800),.q(_w_7801));
  and_bb g1545(.a(N205_14),.b(N443_16),.q(_w_13923));
  and_bi g1488(.a(n1487_0),.b(n1466_0),.q(n1488));
  bfr _b_6546(.a(_w_8448),.q(_w_8449));
  and_bi g1548(.a(n1479_1),.b(n1482_1),.q(n1548));
  bfr _b_10124(.a(_w_12026),.q(n380));
  bfr _b_11358(.a(_w_13260),.q(_w_13261));
  and_bb g1553(.a(n1550_1),.b(n1551_1),.q(_w_13927));
  and_bi g902(.a(n901_0),.b(n830_0),.q(n902));
  bfr _b_5624(.a(_w_7526),.q(_w_7527));
  bfr _b_10657(.a(_w_12559),.q(_w_12560));
  bfr _b_6167(.a(_w_8069),.q(_w_8070));
  bfr _b_6218(.a(_w_8120),.q(_w_8121));
  or_bb g651(.a(n649_0),.b(n650),.q(n651));
  and_bi g1562(.a(n1547_1),.b(n1560_1),.q(_w_13933));
  bfr _b_12928(.a(_w_14830),.q(n542_1));
  spl2 g1136_s_0(.a(n1136),.q0(n1136_0),.q1(n1136_1));
  bfr _b_9861(.a(_w_11763),.q(_w_11764));
  or_bb g1563(.a(n1561_0),.b(n1562),.q(n1563));
  bfr _b_10343(.a(_w_12245),.q(_w_12246));
  or_bb g472(.a(n451_0),.b(n471_0),.q(n472));
  or_bb g1564(.a(n1546_0),.b(n1563_0),.q(n1564));
  and_bb g1565(.a(n1546_1),.b(n1563_1),.q(_w_13938));
  bfr _b_3584(.a(_w_5486),.q(_w_5487));
  spl2 g528_s_0(.a(n528),.q0(n528_0),.q1(n528_1));
  and_bi g1566(.a(n1564_0),.b(n1565),.q(n1566));
  bfr _b_4872(.a(_w_6774),.q(_w_6775));
  bfr _b_10065(.a(_w_11967),.q(_w_11968));
  and_bb g457(.a(N188_5),.b(N273_15),.q(n457));
  and_bi g1712(.a(n1710_0),.b(n1711),.q(n1712));
  bfr _b_8752(.a(_w_10654),.q(_w_10655));
  bfr _b_5343(.a(_w_7245),.q(_w_7246));
  and_bi g644(.a(n634_1),.b(n642_1),.q(_w_13939));
  spl2 g1157_s_0(.a(n1157),.q0(n1157_0),.q1(n1157_1));
  bfr _b_4537(.a(_w_6439),.q(_w_6440));
  and_bi g1567(.a(n1566_0),.b(n1545_0),.q(n1567));
  bfr _b_7485(.a(_w_9387),.q(_w_9388));
  spl2 g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1));
  or_bb g1570(.a(n1544_0),.b(n1569_0),.q(n1570));
  spl2 g596_s_0(.a(n596),.q0(n596_0),.q1(n596_1));
  and_bi g1574(.a(n1543_1),.b(n1572_1),.q(_w_13941));
  bfr _b_13889(.a(_w_15791),.q(_w_15727));
  bfr _b_6965(.a(_w_8867),.q(_w_8868));
  bfr _b_9599(.a(_w_11501),.q(_w_11502));
  bfr _b_4963(.a(_w_6865),.q(_w_6866));
  bfr _b_11866(.a(_w_13768),.q(n1448));
  bfr _b_11048(.a(_w_12950),.q(_w_12951));
  bfr _b_3645(.a(_w_5547),.q(_w_5548));
  and_bi g516(.a(n514_0),.b(n515),.q(n516));
  or_bb g1576(.a(n1542_0),.b(n1575_0),.q(n1576));
  bfr _b_4675(.a(_w_6577),.q(_w_6578));
  bfr _b_5463(.a(_w_7365),.q(_w_7366));
  and_bb g1577(.a(n1542_1),.b(n1575_1),.q(_w_13942));
  bfr _b_5454(.a(_w_7356),.q(_w_7357));
  and_bi g1580(.a(n1541_1),.b(n1578_1),.q(_w_13943));
  bfr _b_9285(.a(_w_11187),.q(_w_11188));
  spl2 g992_s_0(.a(n992),.q0(n992_0),.q1(_w_13944));
  or_bb g600(.a(n523_0),.b(n599_0),.q(n600));
  spl4L N18_s_4(.a(N18_3),.q0(N18_16),.q1(N18_17),.q2(N18_18),.q3(N18_19));
  bfr _b_11518(.a(_w_13420),.q(_w_13421));
  bfr _b_7352(.a(_w_9254),.q(_w_9255));
  bfr _b_13981(.a(_w_15883),.q(_w_15884));
  spl2 g619_s_0(.a(n619),.q0(n619_0),.q1(n619_1));
  bfr _b_5874(.a(_w_7776),.q(_w_7777));
  bfr _b_7416(.a(_w_9318),.q(_w_9319));
  and_bb g43(.a(N273_6),.b(N35_5),.q(n43));
  bfr _b_5115(.a(_w_7017),.q(_w_7018));
  and_bb g1583(.a(n1540_1),.b(n1581_1),.q(_w_13949));
  spl2 g845_s_0(.a(n845),.q0(n845_0),.q1(n845_1));
  bfr _b_8465(.a(_w_10367),.q(_w_10368));
  bfr _b_13827(.a(_w_15729),.q(_w_15730));
  spl2 g1755_s_0(.a(n1755),.q0(n1755_0),.q1(n1755_1));
  or_bb g1587(.a(n1585_0),.b(n1586),.q(n1587));
  and_bb g1186(.a(N256_17),.b(N324_19),.q(_w_12964));
  bfr _b_10246(.a(_w_12148),.q(_w_12149));
  or_bb g1588(.a(n1538_0),.b(n1587_0),.q(n1588));
  bfr _b_4908(.a(_w_6810),.q(_w_6811));
  and_bi g259(.a(n258_0),.b(n242_0),.q(n259));
  bfr _b_5833(.a(_w_7735),.q(_w_7736));
  spl2 g74_s_0(.a(n74),.q0(n74_0),.q1(n74_1));
  bfr _b_8293(.a(_w_10195),.q(_w_10196));
  and_bb g975(.a(n959_1),.b(n973_1),.q(_w_13951));
  bfr _b_14024(.a(_w_15926),.q(_w_15927));
  bfr _b_4120(.a(_w_6022),.q(_w_6023));
  bfr _b_4092(.a(_w_5994),.q(_w_5995));
  and_bi g1180(.a(n1095_1),.b(n1098_1),.q(n1180));
  and_bi g1598(.a(n1535_1),.b(n1596_1),.q(_w_13957));
  bfr _b_7880(.a(_w_9782),.q(_w_9783));
  and_bi g1603(.a(n1602_0),.b(n1533_0),.q(n1603));
  bfr _b_4785(.a(_w_6687),.q(_w_6688));
  bfr _b_4701(.a(_w_6603),.q(_w_6604));
  bfr _b_8711(.a(_w_10613),.q(_w_10614));
  bfr _b_4270(.a(_w_6172),.q(n911_1));
  bfr _b_9894(.a(_w_11796),.q(_w_11797));
  and_bi g1453(.a(n1440_1),.b(n1443_1),.q(n1453));
  and_bi g1609(.a(n1588_1),.b(n1591_1),.q(n1609));
  bfr _b_14169(.a(_w_16071),.q(_w_16072));
  bfr _b_3965(.a(_w_5867),.q(_w_5868));
  bfr _b_6525(.a(_w_8427),.q(_w_8428));
  bfr _b_14253(.a(_w_16155),.q(_w_16156));
  spl2 g73_s_0(.a(n73),.q0(n73_0),.q1(n73_1));
  bfr _b_5945(.a(_w_7847),.q(_w_7848));
  bfr _b_11300(.a(_w_13202),.q(_w_13203));
  bfr _b_3604(.a(_w_5506),.q(_w_5507));
  bfr _b_7081(.a(_w_8983),.q(_w_8984));
  bfr _b_12597(.a(_w_14499),.q(_w_14500));
  bfr _b_9939(.a(_w_11841),.q(n1044));
  bfr _b_10000(.a(_w_11902),.q(_w_11903));
  bfr _b_5820(.a(_w_7722),.q(_w_7723));
  and_bi g1622(.a(n1552_1),.b(n1555_1),.q(n1622));
  bfr _b_6206(.a(_w_8108),.q(_w_8109));
  bfr _b_12087(.a(_w_13989),.q(_w_13990));
  and_bb g1624(.a(n1621_1),.b(n1622_1),.q(_w_13970));
  and_bi g171(.a(n170_0),.b(n138_0),.q(n171));
  spl2 g766_s_0(.a(n766),.q0(n766_0),.q1(_w_13971));
  or_bb g544(.a(n455_1),.b(n543_0),.q(_w_13975));
  spl2 g133_s_0(.a(n133),.q0(n133_0),.q1(n133_1));
  and_bi g1625(.a(n1623_0),.b(n1624),.q(n1625));
  bfr _b_4515(.a(_w_6417),.q(_w_6418));
  bfr _b_3679(.a(_w_5581),.q(_w_5582));
  bfr _b_11019(.a(_w_12921),.q(_w_12922));
  spl2 g1410_s_0(.a(n1410),.q0(n1410_0),.q1(_w_14226));
  bfr _b_8211(.a(_w_10113),.q(_w_10114));
  spl2 g856_s_0(.a(n856),.q0(n856_0),.q1(n856_1));
  or_bb g1582(.a(n1540_0),.b(n1581_0),.q(n1582));
  spl2 g1854_s_0(.a(n1854),.q0(n1854_0),.q1(n1854_1));
  spl2 g1482_s_0(.a(n1482),.q0(n1482_0),.q1(n1482_1));
  and_bb g547(.a(n456_2),.b(n545_1),.q(_w_13948));
  bfr _b_7394(.a(_w_9296),.q(_w_9297));
  and_bi g1826(.a(n1788_1),.b(n1791_1),.q(n1826));
  bfr _b_3638(.a(_w_5540),.q(_w_5541));
  spl2 g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1));
  spl2 g811_s_0(.a(n811),.q0(n811_0),.q1(n811_1));
  or_bb g1635(.a(n1617_0),.b(n1634_0),.q(n1635));
  and_bi g1481(.a(n1479_0),.b(n1480),.q(n1481));
  bfr _b_8031(.a(_w_9933),.q(_w_9934));
  bfr _b_5239(.a(_w_7141),.q(_w_7142));
  spl4L N69_s_3(.a(N69_2),.q0(N69_12),.q1(_w_7479),.q2(_w_7487),.q3(_w_7499));
  or_bb g1640(.a(n1638_0),.b(n1639),.q(n1640));
  bfr _b_14107(.a(_w_16009),.q(_w_16010));
  bfr _b_5111(.a(_w_7013),.q(_w_7014));
  spl4L N324_s_1(.a(N324_0),.q0(N324_4),.q1(N324_5),.q2(N324_6),.q3(N324_7));
  bfr _b_9257(.a(_w_11159),.q(_w_11160));
  and_bi g177(.a(n176_0),.b(n136_0),.q(n177));
  or_bb g1641(.a(n1615_0),.b(n1640_0),.q(n1641));
  spl2 g405_s_0(.a(n405),.q0(n405_0),.q1(n405_1));
  bfr _b_7500(.a(_w_9402),.q(_w_9403));
  and_bb g1642(.a(n1615_1),.b(n1640_1),.q(_w_13977));
  and_bi g1644(.a(n1643_0),.b(n1614_0),.q(n1644));
  bfr _b_4402(.a(_w_6304),.q(n635_1));
  bfr _b_4101(.a(_w_6003),.q(_w_6004));
  bfr _b_5413(.a(_w_7315),.q(_w_7316));
  bfr _b_10192(.a(_w_12094),.q(n355));
  spl4L N1_s_1(.a(N1_0),.q0(N1_4),.q1(N1_5),.q2(N1_6),.q3(N1_7));
  bfr _b_7057(.a(_w_8959),.q(n830));
  bfr _b_3838(.a(_w_5740),.q(_w_5741));
  or_bb g1646(.a(n1644_0),.b(n1645),.q(n1646));
  or_bb g1647(.a(n1613_0),.b(n1646_0),.q(n1647));
  bfr _b_8859(.a(_w_10761),.q(_w_10762));
  spl2 g288_s_0(.a(n288),.q0(n288_0),.q1(n288_1));
  and_bb g791(.a(n721_1),.b(n789_1),.q(_w_13978));
  bfr _b_11077(.a(_w_12979),.q(n1189));
  spl2 g261_s_0(.a(n261),.q0(n261_0),.q1(n261_1));
  and_bi g1649(.a(n1647_0),.b(n1648),.q(n1649));
  and_bb g826(.a(N477_7),.b(N52_16),.q(n826));
  bfr _b_5735(.a(_w_7637),.q(_w_7638));
  spl2 g490_s_0(.a(n490),.q0(n490_0),.q1(_w_12406));
  or_bb g1652(.a(n1650_0),.b(n1651),.q(n1652));
  or_bb g1653(.a(n1611_0),.b(n1652_0),.q(n1653));
  bfr _b_6973(.a(_w_8875),.q(_w_8876));
  bfr _b_7448(.a(_w_9350),.q(_w_9351));
  and_bi g1663(.a(n1608_1),.b(n1661_1),.q(_w_13985));
  or_bb g1664(.a(n1662_0),.b(n1663),.q(n1664));
  bfr _b_10071(.a(_w_11973),.q(_w_11974));
  spl2 g557_s_0(.a(n557),.q0(n557_0),.q1(n557_1));
  bfr _b_10776(.a(_w_12678),.q(_w_12679));
  bfr _b_10005(.a(_w_11907),.q(_w_11908));
  or_bb g1665(.a(n1607_0),.b(n1664_0),.q(_w_13986));
  bfr _b_5983(.a(_w_7885),.q(_w_7886));
  bfr _b_8953(.a(_w_10855),.q(_w_10856));
  bfr _b_8280(.a(_w_10182),.q(n172));
  and_bb g163(.a(n141_1),.b(n161_1),.q(_w_10560));
  and_bi g1668(.a(n1667_0),.b(n1606_0),.q(n1668));
  spl2 g1880_s_0(.a(n1880),.q0(n1880_0),.q1(n1880_1));
  bfr _b_12353(.a(_w_14255),.q(_w_14256));
  bfr _b_3997(.a(_w_5899),.q(_w_5900));
  bfr _b_9049(.a(_w_10951),.q(_w_10952));
  spl2 g754_s_0(.a(n754),.q0(n754_0),.q1(_w_14038));
  bfr _b_13629(.a(N188),.q(_w_15531));
  and_bb g1675(.a(N171_18),.b(N511_14),.q(_w_14042));
  bfr _b_11847(.a(_w_13749),.q(n466_1));
  and_bi g1676(.a(n1647_1),.b(n1650_1),.q(n1676));
  or_bb g558(.a(n537_0),.b(n557_0),.q(n558));
  spl2 g1752_s_0(.a(n1752),.q0(n1752_0),.q1(n1752_1));
  and_bb g281(.a(n235_1),.b(n279_1),.q(_w_14078));
  bfr _b_7823(.a(_w_9725),.q(_w_9726));
  and_bb g1677(.a(N188_17),.b(N494_15),.q(_w_14079));
  and_bb g1879(.a(N256_6),.b(N511_19),.q(_w_14087));
  and_bi g945(.a(n899_1),.b(n902_1),.q(n945));
  and_bi g1791(.a(n1790_0),.b(n1785_0),.q(n1791));
  and_bi g879(.a(n838_1),.b(n877_1),.q(_w_14107));
  bfr _b_8956(.a(_w_10858),.q(n1456));
  and_bi g1680(.a(n1635_1),.b(n1638_1),.q(n1680));
  bfr _b_12602(.a(_w_14504),.q(_w_14505));
  bfr _b_11830(.a(_w_13732),.q(_w_13733));
  and_bi g315(.a(n314_0),.b(n306_0),.q(n315));
  bfr _b_7972(.a(_w_9874),.q(_w_9875));
  bfr _b_7681(.a(_w_9583),.q(n310));
  bfr _b_7751(.a(_w_9653),.q(_w_9654));
  bfr _b_13828(.a(_w_15730),.q(_w_15731));
  bfr _b_5156(.a(_w_7058),.q(_w_7059));
  and_bi g1682(.a(n1629_1),.b(n1632_1),.q(n1682));
  bfr _b_6376(.a(_w_8278),.q(_w_8279));
  bfr _b_9104(.a(_w_11006),.q(_w_11007));
  and_bi g1889(.a(n1887_0),.b(n1888),.q(n1889));
  bfr _b_9557(.a(_w_11459),.q(_w_11460));
  bfr _b_4920(.a(_w_6822),.q(_w_6823));
  bfr _b_10788(.a(_w_12690),.q(_w_12691));
  and_bb g1466(.a(N205_13),.b(N426_16),.q(n1466));
  bfr _b_9237(.a(_w_11139),.q(_w_11140));
  and_bi g966(.a(n964_1),.b(n963_1),.q(_w_14108));
  bfr _b_12129(.a(_w_14031),.q(_w_14032));
  spl2 g1827_s_0(.a(n1827),.q0(n1827_0),.q1(_w_14230));
  and_bi g1688(.a(n1686_0),.b(n1687),.q(n1688));
  spl4L N205_s_3(.a(N205_2),.q0(N205_12),.q1(_w_7964),.q2(_w_7972),.q3(_w_7984));
  bfr _b_7952(.a(_w_9854),.q(_w_9855));
  bfr _b_7071(.a(_w_8973),.q(_w_8974));
  bfr _b_3769(.a(_w_5671),.q(_w_5672));
  bfr _b_5061(.a(_w_6963),.q(_w_6964));
  spl2 g1488_s_0(.a(n1488),.q0(n1488_0),.q1(n1488_1));
  bfr _b_4099(.a(_w_6001),.q(_w_6002));
  spl2 g772_s_0(.a(n772),.q0(n772_0),.q1(_w_14109));
  and_bi g1690(.a(n1683_1),.b(n1688_1),.q(_w_14113));
  and_bi g1774(.a(n1773_0),.b(n1728_0),.q(n1774));
  bfr _b_5730(.a(_w_7632),.q(_w_7633));
  bfr _b_4645(.a(_w_6547),.q(_w_6548));
  bfr _b_4569(.a(_w_6471),.q(_w_6472));
  or_bb g1692(.a(n1682_0),.b(n1691_0),.q(n1692));
  bfr _b_4071(.a(_w_5973),.q(_w_5974));
  and_bi g1299(.a(n1297_0),.b(n1298),.q(n1299));
  bfr _b_5932(.a(_w_7834),.q(_w_7835));
  bfr _b_12096(.a(_w_13998),.q(_w_13999));
  and_bi g1633(.a(n1618_1),.b(n1631_1),.q(_w_13976));
  spl2 g837_s_0(.a(n837),.q0(n837_0),.q1(n837_1));
  bfr _b_3970(.a(_w_5872),.q(N239_14));
  bfr _b_3713(.a(_w_5615),.q(_w_5616));
  bfr _b_9647(.a(_w_11549),.q(_w_11550));
  bfr _b_13285(.a(_w_15187),.q(_w_15188));
  spl2 g1823_s_0(.a(n1823),.q0(n1823_0),.q1(n1823_1));
  bfr _b_9231(.a(_w_11133),.q(n1849));
  bfr _b_10317(.a(_w_12219),.q(_w_12220));
  spl2 g989_s_0(.a(n989),.q0(n989_0),.q1(n989_1));
  and_bi g165(.a(n164_0),.b(n140_0),.q(n165));
  bfr _b_8721(.a(_w_10623),.q(n166));
  spl2 g253_s_0(.a(n253),.q0(n253_0),.q1(n253_1));
  bfr _b_8947(.a(_w_10849),.q(_w_10850));
  spl2 g1582_s_0(.a(n1582),.q0(n1582_0),.q1(_w_14118));
  bfr _b_13408(.a(_w_15310),.q(n263));
  or_bb g1709(.a(n1707_0),.b(n1708),.q(n1709));
  bfr _b_4909(.a(_w_6811),.q(_w_6812));
  bfr _b_10040(.a(_w_11942),.q(_w_11943));
  and_bi g878(.a(n877_0),.b(n838_0),.q(n878));
  or_bb g1710(.a(n1676_0),.b(n1709_0),.q(n1710));
  bfr _b_9081(.a(_w_10983),.q(_w_10984));
  bfr _b_3878(.a(_w_5780),.q(_w_5781));
  and_bi g1713(.a(n1712_0),.b(n1675_0),.q(n1713));
  bfr _b_12281(.a(_w_14183),.q(_w_14184));
  bfr _b_4781(.a(_w_6683),.q(_w_6684));
  bfr _b_9493(.a(_w_11395),.q(N35_3));
  or_bb g1715(.a(n1713_0),.b(n1714),.q(n1715));
  or_bb g1716(.a(n1674_0),.b(n1715_0),.q(n1716));
  bfr _b_12193(.a(_w_14095),.q(_w_14096));
  bfr _b_10386(.a(_w_12288),.q(_w_12289));
  and_bi g1720(.a(n1673_1),.b(n1718_1),.q(_w_14122));
  and_bb g1723(.a(n1672_1),.b(n1721_1),.q(_w_14151));
  bfr _b_8242(.a(_w_10144),.q(_w_10145));
  spl2 g1830_s_0(.a(n1830),.q0(n1830_0),.q1(n1830_1));
  bfr _b_10304(.a(_w_12206),.q(n1213));
  bfr _b_3605(.a(_w_5507),.q(_w_5508));
  and_bi g1726(.a(n1671_1),.b(n1724_1),.q(_w_14152));
  spl2 g33_s_0(.a(n33),.q0(_w_5559),.q1(n33_1));
  and_bb g1853(.a(N222_5),.b(N528_17),.q(_w_14153));
  and_bb g1730(.a(N171_19),.b(N528_14),.q(_w_14177));
  bfr _b_9938(.a(_w_11840),.q(n94_1));
  or_bb g324(.a(n303_0),.b(n323_0),.q(n324));
  spl2 g1841_s_0(.a(n1841),.q0(n1841_0),.q1(n1841_1));
  bfr _b_3766(.a(_w_5668),.q(_w_5669));
  and_bi g1024(.a(n1022_0),.b(n1023),.q(n1024));
  bfr _b_8564(.a(_w_10466),.q(_w_10467));
  spl4L N409_s_4(.a(N409_3),.q0(N409_16),.q1(N409_17),.q2(N409_18),.q3(N409_19));
  and_bi g568(.a(n534_1),.b(n566_1),.q(_w_14217));
  bfr _b_4867(.a(_w_6769),.q(_w_6770));
  or_bb g1691(.a(n1689_0),.b(n1690),.q(n1691));
  bfr _b_3919(.a(_w_5821),.q(_w_5822));
  bfr _b_10653(.a(_w_12555),.q(_w_12556));
  bfr _b_10641(.a(_w_12543),.q(_w_12544));
  and_bb g1736(.a(N222_8),.b(N477_17),.q(n1736));
  spl2 g540_s_0(.a(n540),.q0(n540_0),.q1(n540_1));
  bfr _b_10780(.a(_w_12682),.q(_w_12683));
  spl2 g1866_s_0(.a(n1866),.q0(n1866_0),.q1(n1866_1));
  or_bb g1741(.a(n1739_0),.b(n1740_0),.q(n1741));
  bfr _b_8834(.a(_w_10736),.q(_w_10737));
  and_bb g1846(.a(n1819_1),.b(n1844_1),.q(_w_14235));
  bfr _b_3542(.a(_w_5444),.q(_w_5445));
  bfr _b_7167(.a(_w_9069),.q(_w_9070));
  and_bi g1203(.a(n1202_0),.b(n1181_0),.q(n1203));
  and_bi g1745(.a(n1738_1),.b(n1743_1),.q(_w_14276));
  or_bb g1747(.a(n1737_0),.b(n1746_0),.q(n1747));
  bfr _b_6353(.a(_w_8255),.q(_w_8256));
  and_bb g95(.a(n73_1),.b(n93_1),.q(_w_12517));
  bfr _b_3530(.a(_w_5432),.q(_w_5433));
  bfr _b_14011(.a(_w_15913),.q(_w_15914));
  spl2 g438_s_0(.a(n438),.q0(n438_0),.q1(n438_1));
  bfr _b_3820(.a(_w_5722),.q(_w_5723));
  and_bi g1790(.a(n1788_0),.b(n1789),.q(n1790));
  spl2 g1303_s_0(.a(n1303),.q0(n1303_0),.q1(_w_6706));
  bfr _b_7626(.a(_w_9528),.q(_w_9529));
  and_bi g1876(.a(n1870_1),.b(n1873_1),.q(n1876));
  bfr _b_10726(.a(_w_12628),.q(n522));
  bfr _b_4915(.a(_w_6817),.q(_w_6818));
  bfr _b_6660(.a(_w_8562),.q(_w_8563));
  or_bb g1753(.a(n1735_0),.b(n1752_0),.q(n1753));
  bfr _b_9199(.a(_w_11101),.q(_w_11102));
  spl2 g1133_s_0(.a(n1133),.q0(n1133_0),.q1(n1133_1));
  bfr _b_12457(.a(_w_14359),.q(_w_14360));
  bfr _b_11514(.a(_w_13416),.q(_w_13417));
  bfr _b_9441(.a(_w_11343),.q(_w_11344));
  and_bi g1756(.a(n1755_0),.b(n1734_0),.q(n1756));
  bfr _b_8436(.a(_w_10338),.q(_w_10339));
  bfr _b_11624(.a(_w_13526),.q(_w_13527));
  spl2 g493_s_0(.a(n493),.q0(n493_0),.q1(n493_1));
  bfr _b_8521(.a(_w_10423),.q(_w_10424));
  bfr _b_13588(.a(_w_15490),.q(_w_15491));
  and_bi g1757(.a(n1734_1),.b(n1755_1),.q(_w_14291));
  bfr _b_13186(.a(_w_15088),.q(n1339_1));
  bfr _b_4296(.a(_w_6198),.q(_w_6199));
  bfr _b_5292(.a(_w_7194),.q(_w_7195));
  bfr _b_3449(.a(_w_5351),.q(_w_5352));
  spl2 g1416_s_0(.a(n1416),.q0(n1416_0),.q1(_w_15062));
  bfr _b_3625(.a(_w_5527),.q(_w_5528));
  bfr _b_10137(.a(_w_12039),.q(_w_12040));
  bfr _b_8086(.a(_w_9988),.q(_w_9989));
  bfr _b_8364(.a(_w_10266),.q(_w_10267));
  bfr _b_11039(.a(_w_12941),.q(_w_12942));
  bfr _b_8429(.a(_w_10331),.q(_w_10332));
  bfr _b_13586(.a(_w_15488),.q(N18_7));
  and_bi g1762(.a(n1761_0),.b(n1732_0),.q(n1762));
  bfr _b_4287(.a(_w_6189),.q(_w_6190));
  bfr _b_7179(.a(_w_9081),.q(_w_9082));
  bfr _b_5234(.a(_w_7136),.q(_w_7137));
  bfr _b_14095(.a(_w_15997),.q(_w_15998));
  bfr _b_9954(.a(_w_11856),.q(_w_11857));
  and_bi g1763(.a(n1732_1),.b(n1761_1),.q(_w_14306));
  bfr _b_6968(.a(_w_8870),.q(_w_8871));
  spl2 g687_s_0(.a(n687),.q0(n687_0),.q1(n687_1));
  and_bb g1766(.a(n1731_1),.b(n1764_1),.q(_w_14307));
  bfr _b_9689(.a(_w_11591),.q(_w_11592));
  and_bi g1768(.a(n1767_0),.b(n1730_0),.q(n1768));
  bfr _b_7164(.a(_w_9066),.q(_w_9067));
  spl4L N341_s_4(.a(N341_3),.q0(N341_16),.q1(N341_17),.q2(N341_18),.q3(N341_19));
  bfr _b_8423(.a(_w_10325),.q(_w_10326));
  and_bi g1775(.a(n1728_1),.b(n1773_1),.q(_w_14340));
  bfr _b_4897(.a(_w_6799),.q(_w_6800));
  and_bb g1783(.a(N222_7),.b(N494_17),.q(_w_14341));
  and_bi g1787(.a(n1741_1),.b(n1744_1),.q(n1787));
  spl2 g682_s_0(.a(n682),.q0(n682_0),.q1(_w_14365));
  bfr _b_6557(.a(_w_8459),.q(_w_8460));
  spl2 g874_s_0(.a(n874),.q0(n874_0),.q1(n874_1));
  and_bi g943(.a(n905_1),.b(n908_1),.q(n943));
  and_bb g234(.a(N18_11),.b(N392_5),.q(n234));
  spl2 g829_s_0(.a(n829),.q0(n829_0),.q1(n829_1));
  and_bi g1872(.a(n1870_0),.b(n1871),.q(n1872));
  bfr _b_9160(.a(_w_11062),.q(n1717));
  and_bb g538(.a(N154_7),.b(N324_13),.q(_w_13887));
  or_bb g1793(.a(n1791_0),.b(n1792),.q(n1793));
  spl4L N69_s_1(.a(N69_0),.q0(N69_4),.q1(N69_5),.q2(_w_14370),.q3(_w_14372));
  or_bb g99(.a(n97_0),.b(n98),.q(_w_14374));
  bfr _b_6698(.a(_w_8600),.q(_w_8601));
  and_bi g357(.a(n356_0),.b(n292_0),.q(n357));
  bfr _b_4360(.a(_w_6262),.q(_w_6263));
  spl2 g1606_s_0(.a(n1606),.q0(n1606_0),.q1(n1606_1));
  bfr _b_7150(.a(_w_9052),.q(_w_9053));
  bfr _b_10187(.a(_w_12089),.q(_w_12090));
  bfr _b_3937(.a(_w_5839),.q(_w_5840));
  and_bi g1643(.a(n1641_0),.b(n1642),.q(n1643));
  and_bi g1796(.a(n1794_0),.b(n1795),.q(n1796));
  bfr _b_8493(.a(_w_10395),.q(_w_10396));
  and_bi g1797(.a(n1796_0),.b(n1783_0),.q(n1797));
  bfr _b_9548(.a(_w_11450),.q(_w_11451));
  and_bi g1835(.a(n1833_0),.b(n1834),.q(n1835));
  bfr _b_8895(.a(_w_10797),.q(_w_10798));
  and_bb g1801(.a(n1782_1),.b(n1799_1),.q(_w_14523));
  spl2 g1305_s_0(.a(n1305),.q0(n1305_0),.q1(n1305_1));
  bfr _b_7996(.a(_w_9898),.q(_w_9899));
  bfr _b_14051(.a(_w_15953),.q(_w_15954));
  bfr _b_6307(.a(_w_8209),.q(_w_8210));
  and_bi g1802(.a(n1800_0),.b(n1801),.q(n1802));
  bfr _b_4272(.a(_w_6174),.q(_w_6175));
  bfr _b_11804(.a(_w_13706),.q(_w_13707));
  bfr _b_3612(.a(_w_5514),.q(_w_5515));
  bfr _b_8290(.a(_w_10192),.q(_w_10193));
  and_bb g734(.a(N188_7),.b(N324_15),.q(_w_9163));
  and_bi g1501(.a(n1462_1),.b(n1499_1),.q(_w_12857));
  and_bb g1772(.a(n1729_1),.b(n1770_1),.q(_w_13436));
  bfr _b_4495(.a(_w_6397),.q(_w_6398));
  and_bi g1815(.a(n1814_0),.b(n1777_0),.q(n1815));
  bfr _b_12623(.a(_w_14525),.q(_w_14526));
  and_bi g1818(.a(n1812_1),.b(n1815_1),.q(n1818));
  spl2 g1267_s_0(.a(n1267),.q0(n1267_0),.q1(n1267_1));
  bfr _b_6327(.a(_w_8229),.q(_w_8230));
  bfr _b_12067(.a(_w_13969),.q(n1618));
  and_bb g1824(.a(N239_17),.b(N494_18),.q(_w_14557));
  and_bb g1825(.a(N256_8),.b(N477_19),.q(_w_14565));
  and_bb g467(.a(n453_1),.b(n465_1),.q(_w_14569));
  spl2 g561_s_0(.a(n561),.q0(n561_0),.q1(n561_1));
  bfr _b_7323(.a(_w_9225),.q(n1278));
  or_bb g1838(.a(n1836_0),.b(n1837),.q(n1838));
  bfr _b_7355(.a(_w_9257),.q(_w_9258));
  bfr _b_7486(.a(_w_9388),.q(_w_9389));
  and_bi g1836(.a(n1835_0),.b(n1822_0),.q(n1836));
  and_bb g1732(.a(N188_18),.b(N511_15),.q(_w_14201));
  spl2 g730_s_0(.a(n730),.q0(n730_0),.q1(n730_1));
  spl2 g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1));
  spl2 g1877_s_0(.a(n1877),.q0(n1877_0),.q1(n1877_1));
  bfr _b_10766(.a(_w_12668),.q(_w_12669));
  bfr _b_5590(.a(_w_7492),.q(_w_7493));
  spl2 g1154_s_0(.a(n1154),.q0(n1154_0),.q1(n1154_1));
  bfr _b_7077(.a(_w_8979),.q(_w_8980));
  and_bi g684(.a(n682_0),.b(n683),.q(n684));
  bfr _b_8101(.a(_w_10003),.q(_w_10004));
  bfr _b_3982(.a(_w_5884),.q(N239_15));
  bfr _b_7070(.a(_w_8972),.q(_w_8973));
  bfr _b_14333(.a(_w_16235),.q(_w_16236));
  bfr _b_7141(.a(_w_9043),.q(_w_9044));
  or_bb g261(.a(n259_0),.b(n260),.q(n261));
  and_bb g1859(.a(n1856_1),.b(n1857_1),.q(_w_14686));
  and_bi g1861(.a(n1860_0),.b(n1855_0),.q(n1861));
  bfr _b_3663(.a(_w_5565),.q(_w_5566));
  and_bi g1868(.a(n1853_1),.b(n1866_1),.q(_w_14687));
  bfr _b_9215(.a(_w_11117),.q(_w_11118));
  spl2 g1590_s_0(.a(n1590),.q0(n1590_0),.q1(n1590_1));
  bfr _b_5419(.a(_w_7321),.q(_w_7322));
  bfr _b_8586(.a(_w_10488),.q(_w_10489));
  bfr _b_10768(.a(_w_12670),.q(_w_12671));
  bfr _b_3509(.a(_w_5411),.q(_w_5412));
  spl2 g1811_s_0(.a(n1811),.q0(n1811_0),.q1(n1811_1));
  bfr _b_8473(.a(_w_10375),.q(_w_10376));
  bfr _b_13809(.a(_w_15711),.q(_w_15712));
  bfr _b_4416(.a(_w_6318),.q(_w_6319));
  and_bi g1874(.a(n1851_1),.b(n1872_1),.q(_w_14688));
  bfr _b_11284(.a(_w_13186),.q(_w_13187));
  and_bi g1877(.a(n1864_1),.b(n1867_1),.q(_w_14689));
  bfr _b_5573(.a(_w_7475),.q(_w_7476));
  spl2 g314_s_0(.a(n314),.q0(n314_0),.q1(n314_1));
  bfr _b_7287(.a(_w_9189),.q(_w_9190));
  bfr _b_7802(.a(_w_9704),.q(_w_9705));
  bfr _b_4190(.a(_w_6092),.q(n802_1));
  spl2 g391_s_0(.a(n391),.q0(n391_0),.q1(n391_1));
  and_bi g1880(.a(n1858_1),.b(n1861_1),.q(n1880));
  bfr _b_11403(.a(_w_13305),.q(_w_13306));
  bfr _b_9351(.a(_w_11253),.q(_w_11254));
  bfr _b_4513(.a(_w_6415),.q(_w_6416));
  bfr _b_11375(.a(_w_13277),.q(_w_13278));
  spl2 g1709_s_0(.a(n1709),.q0(n1709_0),.q1(n1709_1));
  or_bb g382(.a(n308_1),.b(n381_0),.q(n382));
  or_bb g1881(.a(n1879_0),.b(n1880_0),.q(n1881));
  bfr _b_11353(.a(_w_13255),.q(_w_13256));
  spl2 g1576_s_0(.a(n1576),.q0(n1576_0),.q1(_w_14765));
  bfr _b_6577(.a(_w_8479),.q(_w_8480));
  bfr _b_6388(.a(_w_8290),.q(_w_8291));
  and_bi g1884(.a(n1883_0),.b(n1878_0),.q(n1884));
  bfr _b_10129(.a(_w_12031),.q(n278));
  bfr _b_3526(.a(_w_5428),.q(_w_5429));
  bfr _b_3519(.a(_w_5421),.q(_w_5422));
  and_bi g1885(.a(n1878_1),.b(n1883_1),.q(_w_14770));
  and_bb g215(.a(n185_1),.b(n213_1),.q(_w_9956));
  bfr _b_7308(.a(_w_9210),.q(n710));
  and_bb g438(.a(N18_14),.b(N443_5),.q(_w_14819));
  bfr _b_7030(.a(_w_8932),.q(_w_8933));
  and_bb g1888(.a(n1877_1),.b(n1886_1),.q(_w_14823));
  bfr _b_4831(.a(_w_6733),.q(N137_1));
  bfr _b_11888(.a(_w_13790),.q(_w_13791));
  bfr _b_10362(.a(_w_12264),.q(_w_12265));
  bfr _b_3929(.a(_w_5831),.q(_w_5832));
  bfr _b_5317(.a(_w_7219),.q(_w_7220));
  spl2 g1805_s_0(.a(n1805),.q0(n1805_0),.q1(n1805_1));
  bfr _b_13671(.a(_w_15573),.q(_w_15574));
  and_bi g1890(.a(n1889_0),.b(n1876_0),.q(n1890));
  bfr _b_12000(.a(_w_13902),.q(_w_13903));
  bfr _b_7091(.a(_w_8993),.q(_w_8994));
  bfr _b_5284(.a(_w_7186),.q(_w_7187));
  spl2 g1761_s_0(.a(n1761),.q0(n1761_0),.q1(n1761_1));
  or_bb g1895(.a(n1893_0),.b(n1894_0),.q(_w_14833));
  bfr _b_6950(.a(_w_8852),.q(_w_8853));
  bfr _b_13132(.a(_w_15034),.q(_w_15035));
  bfr _b_4921(.a(_w_6823),.q(_w_6824));
  bfr _b_9988(.a(_w_11890),.q(_w_11891));
  and_bb g1897(.a(n1893_1),.b(n1894_1),.q(_w_14885));
  bfr _b_7422(.a(_w_9324),.q(_w_9325));
  bfr _b_8255(.a(_w_10157),.q(_w_10158));
  and_bi g1899(.a(n1898_0),.b(n1896_0),.q(n1899));
  bfr _b_8054(.a(_w_9956),.q(n215));
  and_bi g1750(.a(n1749_0),.b(n1736_0),.q(n1750));
  spl2 g1015_s_0(.a(n1015),.q0(n1015_0),.q1(n1015_1));
  bfr _b_3871(.a(_w_5773),.q(_w_5774));
  bfr _b_9108(.a(_w_11010),.q(n1672));
  or_bb g1902(.a(n1899_1),.b(n1901),.q(N6288));
  bfr _b_8685(.a(_w_10587),.q(_w_10588));
  spl2 g1585_s_0(.a(n1585),.q0(n1585_0),.q1(n1585_1));
  bfr _b_6386(.a(_w_8288),.q(_w_8289));
  spl2 g1894_s_0(.a(n1894),.q0(n1894_0),.q1(n1894_1));
  bfr _b_12378(.a(_w_14280),.q(n60_1));
  bfr _b_4585(.a(_w_6487),.q(_w_6488));
  bfr _b_11898(.a(_w_13800),.q(_w_13801));
  bfr _b_6935(.a(_w_8837),.q(_w_8838));
  spl2 g351_s_0(.a(n351),.q0(n351_0),.q1(n351_1));
  spl2 g1881_s_0(.a(n1881),.q0(n1881_0),.q1(_w_14947));
  bfr _b_5321(.a(_w_7223),.q(_w_7224));
  spl2 g1372_s_0(.a(n1372),.q0(n1372_0),.q1(n1372_1));
  bfr _b_8945(.a(_w_10847),.q(_w_10848));
  bfr _b_6054(.a(_w_7956),.q(_w_7957));
  spl2 g1826_s_0(.a(n1826),.q0(n1826_0),.q1(n1826_1));
  and_bb g1074(.a(N239_7),.b(N324_18),.q(_w_13874));
  bfr _b_6590(.a(_w_8492),.q(_w_8493));
  bfr _b_5018(.a(_w_6920),.q(_w_6921));
  and_bb g1041(.a(n1039_1),.b(n937_1),.q(_w_10183));
  and_bi g1740(.a(n1686_1),.b(n1689_1),.q(n1740));
  bfr _b_13598(.a(_w_15500),.q(_w_15501));
  bfr _b_3597(.a(_w_5499),.q(_w_5500));
  bfr _b_11917(.a(_w_13819),.q(_w_13820));
  bfr _b_7082(.a(_w_8984),.q(N188_1));
  bfr _b_9087(.a(_w_10989),.q(_w_10990));
  bfr _b_9293(.a(_w_11195),.q(_w_11196));
  bfr _b_3716(.a(_w_5618),.q(_w_5619));
  and_bi g1104(.a(n1103_0),.b(n1066_0),.q(n1104));
  and_bb g1589(.a(n1538_1),.b(n1587_1),.q(_w_14951));
  spl2 g442_s_0(.a(n442),.q0(n442_0),.q1(n442_1));
  and_bi g971(.a(n970_0),.b(n960_0),.q(n971));
  spl2 g1791_s_0(.a(n1791),.q0(n1791_0),.q1(n1791_1));
  bfr _b_11966(.a(_w_13868),.q(n1510));
  bfr _b_3946(.a(_w_5848),.q(n220_1));
  spl2 g1786_s_0(.a(n1786),.q0(n1786_0),.q1(n1786_1));
  spl2 g1181_s_0(.a(n1181),.q0(n1181_0),.q1(n1181_1));
  bfr _b_13424(.a(_w_15326),.q(_w_15327));
  spl2 g1778_s_0(.a(n1778),.q0(n1778_0),.q1(n1778_1));
  spl2 g1771_s_0(.a(n1771),.q0(n1771_0),.q1(_w_14956));
  or_bb g1357(.a(n1267_0),.b(n1356_0),.q(_w_14960));
  bfr _b_10581(.a(_w_12483),.q(_w_12484));
  bfr _b_5814(.a(_w_7716),.q(_w_7717));
  bfr _b_7617(.a(_w_9519),.q(_w_9520));
  bfr _b_6657(.a(_w_8559),.q(n1099));
  bfr _b_3729(.a(_w_5631),.q(_w_5632));
  bfr _b_5709(.a(_w_7611),.q(_w_7612));
  spl2 g1770_s_0(.a(n1770),.q0(n1770_0),.q1(n1770_1));
  spl2 g1768_s_0(.a(n1768),.q0(n1768_0),.q1(n1768_1));
  spl2 g1765_s_0(.a(n1765),.q0(n1765_0),.q1(_w_14969));
  bfr _b_7997(.a(_w_9899),.q(_w_9900));
  or_bb g588(.a(n527_0),.b(n587_0),.q(n588));
  spl2 g1753_s_0(.a(n1753),.q0(n1753_0),.q1(_w_14973));
  spl2 g1672_s_0(.a(n1672),.q0(n1672_0),.q1(n1672_1));
  bfr _b_13331(.a(_w_15233),.q(_w_15234));
  bfr _b_5223(.a(_w_7125),.q(_w_7126));
  spl2 g247_s_0(.a(n247),.q0(n247_0),.q1(n247_1));
  spl2 g1544_s_0(.a(n1544),.q0(n1544_0),.q1(n1544_1));
  spl2 g705_s_0(.a(n705),.q0(n705_0),.q1(n705_1));
  spl2 g1733_s_0(.a(n1733),.q0(n1733_0),.q1(n1733_1));
  spl2 g1822_s_0(.a(n1822),.q0(n1822_0),.q1(n1822_1));
  bfr _b_13297(.a(_w_15199),.q(_w_15200));
  bfr _b_7478(.a(_w_9380),.q(_w_9381));
  bfr _b_3692(.a(_w_5594),.q(_w_5595));
  bfr _b_12172(.a(_w_14074),.q(_w_14075));
  bfr _b_8667(.a(_w_10569),.q(_w_10570));
  bfr _b_10068(.a(_w_11970),.q(_w_11971));
  bfr _b_8787(.a(_w_10689),.q(_w_10690));
  and_bi g919(.a(n917_0),.b(n918),.q(n919));
  spl2 g1706_s_0(.a(n1706),.q0(n1706_0),.q1(n1706_1));
  bfr _b_7665(.a(_w_9567),.q(n160));
  spl2 g220_s_0(.a(n220),.q0(n220_0),.q1(_w_5845));
  spl2 g1521_s_0(.a(n1521),.q0(n1521_0),.q1(_w_15097));
  and_bi g861(.a(n844_1),.b(n859_1),.q(_w_8780));
  bfr _b_3723(.a(_w_5625),.q(_w_5626));
  spl2 g1205_s_0(.a(n1205),.q0(n1205_0),.q1(n1205_1));
  and_bb g1539(.a(N154_17),.b(N494_13),.q(_w_14981));
  and_bb g436(.a(N1_15),.b(N460_4),.q(_w_14989));
  spl2 g1689_s_0(.a(n1689),.q0(n1689_0),.q1(n1689_1));
  bfr _b_13684(.a(_w_15586),.q(_w_15587));
  bfr _b_9101(.a(_w_11003),.q(_w_11004));
  bfr _b_5004(.a(_w_6906),.q(_w_6907));
  and_bi g1444(.a(n1365_1),.b(n1442_1),.q(_w_15001));
  spl2 g1688_s_0(.a(n1688),.q0(n1688_0),.q1(n1688_1));
  bfr _b_5542(.a(_w_7444),.q(_w_7445));
  spl2 g1685_s_0(.a(n1685),.q0(n1685_0),.q1(n1685_1));
  and_bi g1174(.a(n1113_1),.b(n1116_1),.q(n1174));
  spl2 g1683_s_0(.a(n1683),.q0(n1683_0),.q1(n1683_1));
  bfr _b_9527(.a(_w_11429),.q(_w_11430));
  spl2 g1607_s_0(.a(n1607),.q0(n1607_0),.q1(n1607_1));
  spl2 g1682_s_0(.a(n1682),.q0(n1682_0),.q1(n1682_1));
  spl2 g1363_s_0(.a(n1363),.q0(n1363_0),.q1(n1363_1));
  spl2 g1676_s_0(.a(n1676),.q0(n1676_0),.q1(n1676_1));
  spl2 g1658_s_0(.a(n1658),.q0(n1658_0),.q1(n1658_1));
  bfr _b_6695(.a(_w_8597),.q(_w_8598));
  bfr _b_4229(.a(_w_6131),.q(_w_6132));
  spl2 g623_s_0(.a(n623),.q0(n623_0),.q1(n623_1));
  bfr _b_7042(.a(_w_8944),.q(_w_8945));
  bfr _b_7271(.a(_w_9173),.q(_w_9174));
  bfr _b_9124(.a(_w_11026),.q(n325));
  bfr _b_14138(.a(_w_16040),.q(_w_16041));
  or_bb g1236(.a(n1170_0),.b(n1235_0),.q(n1236));
  spl2 g1656_s_0(.a(n1656),.q0(n1656_0),.q1(n1656_1));
  and_bb g485(.a(n447_1),.b(n483_1),.q(_w_15006));
  bfr _b_3470(.a(_w_5372),.q(_w_5373));
  spl2 g1649_s_0(.a(n1649),.q0(n1649_0),.q1(n1649_1));
  and_bi g1901(.a(n1896_1),.b(n1898_1),.q(_w_14938));
  bfr _b_10134(.a(_w_12036),.q(_w_12037));
  spl4L N290_s_2(.a(N290_1),.q0(N290_8),.q1(N290_9),.q2(N290_10),.q3(N290_11));
  spl2 g1737_s_0(.a(n1737),.q0(n1737_0),.q1(n1737_1));
  spl2 g1644_s_0(.a(n1644),.q0(n1644_0),.q1(n1644_1));
  spl2 g1638_s_0(.a(n1638),.q0(n1638_0),.q1(n1638_1));
  or_bb g1101(.a(n1067_0),.b(n1100_0),.q(n1101));
  spl2 g1632_s_0(.a(n1632),.q0(n1632_0),.q1(n1632_1));
  bfr _b_12473(.a(_w_14375),.q(_w_14376));
  bfr _b_10502(.a(_w_12404),.q(n508_1));
  bfr _b_4633(.a(_w_6535),.q(_w_6536));
  spl2 g1631_s_0(.a(n1631),.q0(n1631_0),.q1(n1631_1));
  bfr _b_9196(.a(_w_11098),.q(_w_11099));
  spl2 g226_s_0(.a(n226),.q0(n226_0),.q1(_w_15011));
  bfr _b_8176(.a(_w_10078),.q(_w_10079));
  spl2 g1626_s_0(.a(n1626),.q0(n1626_0),.q1(n1626_1));
  bfr _b_4725(.a(_w_6627),.q(_w_6628));
  bfr _b_7804(.a(_w_9706),.q(_w_9707));
  spl2 g1722_s_0(.a(n1722),.q0(n1722_0),.q1(_w_15015));
  or_bb g564(.a(n535_0),.b(n563_0),.q(n564));
  spl2 g1503_s_0(.a(n1503),.q0(n1503_0),.q1(_w_15020));
  bfr _b_4425(.a(_w_6327),.q(_w_6328));
  bfr _b_3622(.a(_w_5524),.q(_w_5525));
  spl2 g1615_s_0(.a(n1615),.q0(n1615_0),.q1(n1615_1));
  bfr _b_3636(.a(_w_5538),.q(N52_3));
  spl2 g1603_s_0(.a(n1603),.q0(n1603_0),.q1(n1603_1));
  spl2 g1520_s_0(.a(n1520),.q0(n1520_0),.q1(n1520_1));
  bfr _b_8446(.a(_w_10348),.q(_w_10349));
  spl2 g1593_s_0(.a(n1593),.q0(n1593_0),.q1(n1593_1));
  bfr _b_11108(.a(_w_13010),.q(n1234));
  and_bb g236(.a(N35_10),.b(N375_6),.q(_w_15024));
  bfr _b_11221(.a(_w_13123),.q(_w_13124));
  spl2 g1378_s_0(.a(n1378),.q0(n1378_0),.q1(n1378_1));
  bfr _b_10136(.a(_w_12038),.q(_w_12039));
  spl2 g1655_s_0(.a(n1655),.q0(n1655_0),.q1(n1655_1));
  bfr _b_9858(.a(_w_11760),.q(_w_11761));
  spl2 g1643_s_0(.a(n1643),.q0(n1643_0),.q1(n1643_1));
  spl2 g1551_s_0(.a(n1551),.q0(n1551_0),.q1(n1551_1));
  bfr _b_8125(.a(_w_10027),.q(_w_10028));
  bfr _b_4090(.a(_w_5992),.q(N239_2));
  spl2 g1545_s_0(.a(n1545),.q0(n1545_0),.q1(n1545_1));
  spl2 g1071_s_0(.a(n1071),.q0(n1071_0),.q1(n1071_1));
  bfr _b_4703(.a(_w_6605),.q(_w_6606));
  bfr _b_10189(.a(_w_12091),.q(n1260));
  bfr _b_11745(.a(_w_13647),.q(_w_13648));
  spl2 g1329_s_0(.a(n1329),.q0(n1329_0),.q1(n1329_1));
  bfr _b_11097(.a(_w_12999),.q(n1600));
  spl2 g1537_s_0(.a(n1537),.q0(n1537_0),.q1(n1537_1));
  bfr _b_5110(.a(_w_7012),.q(_w_7013));
  bfr _b_7269(.a(_w_9171),.q(_w_9172));
  bfr _b_13632(.a(N256),.q(_w_15535));
  bfr _b_13320(.a(_w_15222),.q(_w_15223));
  spl2 g584_s_0(.a(n584),.q0(n584_0),.q1(n584_1));
  bfr _b_12852(.a(_w_14754),.q(_w_14755));
  bfr _b_3497(.a(_w_5399),.q(_w_5400));
  and_bb g1620(.a(N239_13),.b(N426_18),.q(n1620));
  bfr _b_13374(.a(_w_15276),.q(_w_15277));
  bfr _b_5119(.a(_w_7021),.q(_w_7022));
  spl2 g211_s_0(.a(n211),.q0(n211_0),.q1(n211_1));
  or_bb g1345(.a(n1271_0),.b(n1344_0),.q(n1345));
  spl2 g1515_s_0(.a(n1515),.q0(n1515_0),.q1(_w_15044));
  spl2 g1297_s_0(.a(n1297),.q0(n1297_0),.q1(_w_13562));
  spl2 g1502_s_0(.a(n1502),.q0(n1502_0),.q1(n1502_1));
  spl2 g1667_s_0(.a(n1667),.q0(n1667_0),.q1(n1667_1));
  spl2 g305_s_0(.a(n305),.q0(n305_0),.q1(n305_1));
  bfr _b_10234(.a(_w_12136),.q(_w_12137));
  spl2 g1493_s_0(.a(n1493),.q0(n1493_0),.q1(n1493_1));
  bfr _b_8543(.a(_w_10445),.q(_w_10446));
  bfr _b_3755(.a(_w_5657),.q(_w_5658));
  bfr _b_8240(.a(_w_10142),.q(_w_10143));
  bfr _b_9332(.a(_w_11234),.q(_w_11235));
  bfr _b_4389(.a(_w_6291),.q(n588_1));
  bfr _b_3415(.a(_w_5317),.q(_w_5318));
  spl2 g1464_s_0(.a(n1464),.q0(n1464_0),.q1(n1464_1));
  bfr _b_4543(.a(_w_6445),.q(_w_6446));
  bfr _b_4141(.a(_w_6043),.q(_w_6044));
  spl4L N273_s_0(.a(_w_15537),.q0(N273_0),.q1(N273_1),.q2(N273_2),.q3(N273_3));
  spl2 g1462_s_0(.a(n1462),.q0(n1462_0),.q1(n1462_1));
  spl2 g628_s_0(.a(n628),.q0(n628_0),.q1(n628_1));
  spl2 g1458_s_0(.a(n1458),.q0(n1458_0),.q1(n1458_1));
  and_bi g745(.a(n744_0),.b(n736_0),.q(n745));
  spl2 g449_s_0(.a(n449),.q0(n449_0),.q1(n449_1));
  bfr _b_4233(.a(_w_6135),.q(_w_6136));
  bfr _b_4130(.a(_w_6032),.q(_w_6033));
  bfr _b_7956(.a(_w_9858),.q(_w_9859));
  bfr _b_8638(.a(_w_10540),.q(_w_10541));
  spl2 g534_s_0(.a(n534),.q0(n534_0),.q1(n534_1));
  spl2 g1445_s_0(.a(n1445),.q0(n1445_0),.q1(n1445_1));
  spl2 g1506_s_0(.a(n1506),.q0(n1506_0),.q1(n1506_1));
  or_bb g196(.a(n146_1),.b(n195_0),.q(n196));
  bfr _b_9958(.a(_w_11860),.q(_w_11861));
  spl2 g579_s_0(.a(n579),.q0(n579_0),.q1(n579_1));
  bfr _b_4383(.a(_w_6285),.q(_w_6286));
  spl2 g1428_s_0(.a(n1428),.q0(n1428_0),.q1(_w_15053));
  and_bi g1198(.a(n1183_1),.b(n1196_1),.q(_w_15057));
  bfr _b_11824(.a(_w_13726),.q(_w_13727));
  bfr _b_5570(.a(_w_7472),.q(_w_7473));
  spl2 g1427_s_0(.a(n1427),.q0(n1427_0),.q1(n1427_1));
  spl2 g1422_s_0(.a(n1422),.q0(n1422_0),.q1(_w_15058));
  spl2 g1785_s_0(.a(n1785),.q0(n1785_0),.q1(n1785_1));
  bfr _b_4570(.a(_w_6472),.q(_w_6473));
  bfr _b_7184(.a(_w_9086),.q(_w_9087));
  bfr _b_6391(.a(_w_8293),.q(_w_8294));
  bfr _b_9536(.a(_w_11438),.q(_w_11439));
  bfr _b_4088(.a(_w_5990),.q(_w_5991));
  spl2 g1460_s_0(.a(n1460),.q0(n1460_0),.q1(n1460_1));
  spl2 g1857_s_0(.a(n1857),.q0(n1857_0),.q1(n1857_1));
  spl2 g1652_s_0(.a(n1652),.q0(n1652_0),.q1(n1652_1));
  bfr _b_9952(.a(_w_11854),.q(_w_11855));
  bfr _b_4996(.a(_w_6898),.q(_w_6899));
  and_bi g476(.a(n450_1),.b(n474_1),.q(_w_15066));
  bfr _b_12107(.a(_w_14009),.q(n1665));
  spl2 g1386_s_0(.a(n1386),.q0(n1386_0),.q1(_w_15067));
  bfr _b_12210(.a(_w_14112),.q(n772_1));
  spl2 g1382_s_0(.a(n1382),.q0(n1382_0),.q1(n1382_1));
  bfr _b_9763(.a(_w_11665),.q(_w_11666));
  and_bi g1170(.a(n1125_1),.b(n1128_1),.q(n1170));
  and_bi g218(.a(n184_1),.b(n216_1),.q(_w_15071));
  bfr _b_12187(.a(_w_14089),.q(_w_14090));
  spl2 g1155_s_0(.a(n1155),.q0(n1155_0),.q1(_w_15072));
  spl2 g1374_s_0(.a(n1374),.q0(n1374_0),.q1(n1374_1));
  spl2 g1788_s_0(.a(n1788),.q0(n1788_0),.q1(_w_15076));
  bfr _b_11154(.a(_w_13056),.q(_w_13057));
  and_bi g92(.a(n74_1),.b(n90_1),.q(_w_15080));
  bfr _b_11985(.a(_w_13887),.q(_w_13888));
  bfr _b_4758(.a(_w_6660),.q(_w_6661));
  spl2 g1739_s_0(.a(n1739),.q0(n1739_0),.q1(n1739_1));
  bfr _b_5172(.a(_w_7074),.q(_w_7075));
  spl2 g1359_s_0(.a(n1359),.q0(n1359_0),.q1(n1359_1));
  and_bi g1140(.a(n1139_0),.b(n1054_0),.q(n1140));
  bfr _b_10025(.a(_w_11927),.q(_w_11928));
  bfr _b_8016(.a(_w_9918),.q(_w_9919));
  spl2 g1345_s_0(.a(n1345),.q0(n1345_0),.q1(_w_15081));
  bfr _b_6251(.a(_w_8153),.q(n1669));
  spl2 g1339_s_0(.a(n1339),.q0(n1339_0),.q1(_w_15085));
  bfr _b_6992(.a(_w_8894),.q(_w_8895));
  bfr _b_14232(.a(_w_16134),.q(_w_16135));
  and_bi g518(.a(n436_1),.b(n516_1),.q(_w_12523));
  spl2 g1327_s_0(.a(n1327),.q0(n1327_0),.q1(_w_15089));
  bfr _b_5021(.a(_w_6923),.q(_w_6924));
  or_bb g280(.a(n235_0),.b(n279_0),.q(n280));
  spl2 g1142_s_0(.a(n1142),.q0(n1142_0),.q1(n1142_1));
  bfr _b_3492(.a(_w_5394),.q(N52_1));
  bfr _b_10028(.a(_w_11930),.q(_w_11931));
  spl2 g1326_s_0(.a(n1326),.q0(n1326_0),.q1(n1326_1));
  spl2 g1317_s_0(.a(n1317),.q0(n1317_0),.q1(n1317_1));
  bfr _b_5672(.a(_w_7574),.q(n1016_1));
  spl2 g1094_s_0(.a(n1094),.q0(n1094_0),.q1(n1094_1));
  and_bi g1551(.a(n1473_1),.b(n1476_1),.q(n1551));
  and_bi g787(.a(n786_0),.b(n722_0),.q(n787));
  bfr _b_7657(.a(_w_9559),.q(_w_9560));
  bfr _b_8401(.a(_w_10303),.q(_w_10304));
  bfr _b_10200(.a(_w_12102),.q(_w_12103));
  spl2 g1369_s_0(.a(n1369),.q0(n1369_0),.q1(n1369_1));
  spl2 g805_s_0(.a(n805),.q0(n805_0),.q1(n805_1));
  bfr _b_9598(.a(_w_11500),.q(_w_11501));
  bfr _b_12114(.a(_w_14016),.q(_w_14017));
  bfr _b_10324(.a(_w_12226),.q(_w_12227));
  spl2 g1538_s_0(.a(n1538),.q0(n1538_0),.q1(n1538_1));
  bfr _b_10097(.a(_w_11999),.q(_w_12000));
  bfr _b_4739(.a(_w_6641),.q(N1_13));
  spl2 g1288_s_0(.a(n1288),.q0(n1288_0),.q1(n1288_1));
  spl2 g1715_s_0(.a(n1715),.q0(n1715_0),.q1(n1715_1));
  bfr _b_4571(.a(_w_6473),.q(_w_6474));
  or_bb g1490(.a(n1488_0),.b(n1489),.q(n1490));
  bfr _b_10173(.a(_w_12075),.q(n413));
  spl2 g1454_s_0(.a(n1454),.q0(n1454_0),.q1(n1454_1));
  bfr _b_12183(.a(_w_14085),.q(_w_14086));
  spl2 g1266_s_0(.a(n1266),.q0(n1266_0),.q1(n1266_1));
  spl2 g457_s_0(.a(n457),.q0(n457_0),.q1(n457_1));
  bfr _b_10583(.a(_w_12485),.q(n824));
  or_bb g88(.a(n75_0),.b(n87_0),.q(n88));
  bfr _b_5388(.a(_w_7290),.q(_w_7291));
  and_bi g603(.a(n602_0),.b(n522_0),.q(n603));
  bfr _b_7631(.a(_w_9533),.q(_w_9534));
  spl2 g1260_s_0(.a(n1260),.q0(n1260_0),.q1(_w_15101));
  bfr _b_14206(.a(N511),.q(_w_16109));
  spl2 g1256_s_0(.a(n1256),.q0(n1256_0),.q1(n1256_1));
  bfr _b_6149(.a(_w_8051),.q(_w_8052));
  spl2 g1253_s_0(.a(n1253),.q0(n1253_0),.q1(n1253_1));
  bfr _b_3851(.a(_w_5753),.q(_w_5754));
  bfr _b_5186(.a(_w_7088),.q(_w_7089));
  spl2 g1381_s_0(.a(n1381),.q0(n1381_0),.q1(n1381_1));
  bfr _b_3740(.a(_w_5642),.q(_w_5643));
  bfr _b_7889(.a(_w_9791),.q(_w_9792));
  spl2 g771_s_0(.a(n771),.q0(n771_0),.q1(n771_1));
  spl2 g1245_s_0(.a(n1245),.q0(n1245_0),.q1(n1245_1));
  or_bb g1218(.a(n1176_0),.b(n1217_0),.q(n1218));
  spl2 g747_s_0(.a(n747),.q0(n747_0),.q1(n747_1));
  bfr _b_4998(.a(_w_6900),.q(_w_6901));
  and_bi g537(.a(n466_1),.b(n469_1),.q(n537));
  bfr _b_6802(.a(_w_8704),.q(_w_8705));
  bfr _b_7468(.a(_w_9370),.q(_w_9371));
  spl2 g1238_s_0(.a(n1238),.q0(n1238_0),.q1(n1238_1));
  bfr _b_12370(.a(_w_14272),.q(_w_14273));
  spl4L N188_s_2(.a(N188_1),.q0(N188_8),.q1(N188_9),.q2(N188_10),.q3(_w_7928));
  spl2 g1232_s_0(.a(n1232),.q0(n1232_0),.q1(n1232_1));
  bfr _b_4646(.a(_w_6548),.q(_w_6549));
  bfr _b_4230(.a(_w_6132),.q(_w_6133));
  and_bb g1284(.a(N205_11),.b(N392_16),.q(n1284));
  bfr _b_9176(.a(_w_11078),.q(_w_11079));
  bfr _b_4713(.a(_w_6615),.q(_w_6616));
  spl2 g1581_s_0(.a(n1581),.q0(n1581_0),.q1(n1581_1));
  bfr _b_5682(.a(_w_7584),.q(_w_7585));
  bfr _b_4163(.a(_w_6065),.q(_w_6066));
  spl2 g1578_s_0(.a(n1578),.q0(n1578_0),.q1(n1578_1));
  spl2 g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1));
  bfr _b_7799(.a(_w_9701),.q(_w_9702));
  spl2 g1212_s_0(.a(n1212),.q0(n1212_0),.q1(_w_15110));
  spl2 g1190_s_0(.a(n1190),.q0(n1190_0),.q1(n1190_1));
  bfr _b_3683(.a(_w_5585),.q(_w_5586));
  bfr _b_6765(.a(_w_8667),.q(_w_8668));
  and_bi g90(.a(n88_0),.b(n89),.q(n90));
  spl2 g1608_s_0(.a(n1608),.q0(n1608_0),.q1(n1608_1));
  spl2 g810_s_0(.a(n810),.q0(n810_0),.q1(n810_1));
  and_bb g313(.a(n246_2),.b(n311_1),.q(_w_15114));
  spl2 g1818_s_0(.a(n1818),.q0(n1818_0),.q1(n1818_1));
  bfr _b_14194(.a(_w_16096),.q(_w_16097));
  bfr _b_4414(.a(_w_6316),.q(n778_1));
  spl2 g1182_s_0(.a(n1182),.q0(n1182_0),.q1(n1182_1));
  spl2 g1861_s_0(.a(n1861),.q0(n1861_0),.q1(n1861_1));
  bfr _b_9675(.a(_w_11577),.q(n1147));
  bfr _b_3719(.a(_w_5621),.q(_w_5622));
  bfr _b_5050(.a(_w_6952),.q(_w_6953));
  bfr _b_8508(.a(_w_10410),.q(_w_10411));
  spl2 g1151_s_0(.a(n1151),.q0(n1151_0),.q1(n1151_1));
  bfr _b_6430(.a(_w_8332),.q(_w_8333));
  spl2 g1018_s_0(.a(n1018),.q0(n1018_0),.q1(n1018_1));
  bfr _b_14091(.a(_w_15993),.q(_w_15994));
  bfr _b_3992(.a(_w_5894),.q(_w_5895));
  bfr _b_5521(.a(_w_7423),.q(_w_7424));
  bfr _b_4503(.a(_w_6405),.q(_w_6406));
  spl2 g1180_s_0(.a(n1180),.q0(n1180_0),.q1(n1180_1));
  bfr _b_7598(.a(_w_9500),.q(_w_9501));
  bfr _b_13226(.a(_w_15128),.q(_w_15129));
  bfr _b_8425(.a(_w_10327),.q(_w_10328));
  spl2 g808_s_0(.a(n808),.q0(n808_0),.q1(_w_15115));
  bfr _b_6024(.a(_w_7926),.q(_w_7927));
  bfr _b_10276(.a(_w_12178),.q(_w_12179));
  spl2 g652_s_0(.a(n652),.q0(n652_0),.q1(_w_15119));
  bfr _b_5163(.a(_w_7065),.q(_w_7066));
  bfr _b_11612(.a(_w_13514),.q(_w_13515));
  spl2 g1152_s_0(.a(n1152),.q0(n1152_0),.q1(n1152_1));
  bfr _b_3750(.a(_w_5652),.q(_w_5653));
  bfr _b_12835(.a(_w_14737),.q(_w_14738));
  bfr _b_12021(.a(_w_13923),.q(_w_13924));
  spl4L N69_s_0(.a(_w_16287),.q0(N69_0),.q1(_w_15123),.q2(_w_15147),.q3(_w_15203));
  spl2 g1148_s_0(.a(n1148),.q0(n1148_0),.q1(n1148_1));
  bfr _b_11899(.a(_w_13801),.q(N103_15));
  bfr _b_7275(.a(_w_9177),.q(_w_9178));
  bfr _b_9638(.a(_w_11540),.q(_w_11541));
  bfr _b_4653(.a(_w_6555),.q(_w_6556));
  bfr _b_9408(.a(_w_11310),.q(_w_11311));
  and_bi g1146(.a(n1145_0),.b(n1052_0),.q(n1146));
  or_bb g1526(.a(n1524_0),.b(n1525),.q(n1526));
  bfr _b_11613(.a(_w_13515),.q(_w_13516));
  bfr _b_9509(.a(_w_11411),.q(_w_11412));
  spl2 g1055_s_0(.a(n1055),.q0(n1055_0),.q1(n1055_1));
  bfr _b_10850(.a(_w_12752),.q(_w_12753));
  bfr _b_7144(.a(_w_9046),.q(_w_9047));
  and_bb g331(.a(n301_1),.b(n329_1),.q(_w_15295));
  spl2 g1106_s_0(.a(n1106),.q0(n1106_0),.q1(n1106_1));
  bfr _b_5506(.a(_w_7408),.q(_w_7409));
  bfr _b_4526(.a(_w_6428),.q(_w_6429));
  bfr _b_6358(.a(_w_8260),.q(_w_8261));
  bfr _b_12613(.a(_w_14515),.q(_w_14516));
  spl2 g1104_s_0(.a(n1104),.q0(n1104_0),.q1(n1104_1));
  bfr _b_5577(.a(_w_7479),.q(_w_7480));
  and_bi g627(.a(n564_1),.b(n567_1),.q(n627));
  spl2 g1290_s_0(.a(n1290),.q0(n1290_0),.q1(n1290_1));
  bfr _b_3481(.a(_w_5383),.q(_w_5384));
  and_bb g407(.a(n369_1),.b(n405_1),.q(_w_8206));
  spl2 g292_s_0(.a(n292),.q0(n292_0),.q1(n292_1));
  bfr _b_12948(.a(_w_14850),.q(_w_14851));
  spl2 g1555_s_0(.a(n1555),.q0(n1555_0),.q1(n1555_1));
  bfr _b_7207(.a(_w_9109),.q(_w_9110));
  spl2 g507_s_0(.a(n507),.q0(n507_0),.q1(n507_1));
  bfr _b_9275(.a(_w_11177),.q(_w_11178));
  bfr _b_8005(.a(_w_9907),.q(_w_9908));
  spl3L g56_s_0(.a(n56),.q0(n56_0),.q1(_w_15296),.q2(_w_15298));
  bfr _b_8623(.a(_w_10525),.q(_w_10526));
  bfr _b_4243(.a(_w_6145),.q(_w_6146));
  bfr _b_9256(.a(_w_11158),.q(_w_11159));
  and_bi g1076(.a(n962_1),.b(n965_1),.q(n1076));
  spl2 g1853_s_0(.a(n1853),.q0(n1853_0),.q1(n1853_1));
  bfr _b_8882(.a(_w_10784),.q(N52_7));
  bfr _b_6238(.a(_w_8140),.q(_w_8141));
  bfr _b_6483(.a(_w_8385),.q(_w_8386));
  bfr _b_9646(.a(_w_11548),.q(_w_11549));
  bfr _b_10896(.a(_w_12798),.q(_w_12799));
  and_bi g1382(.a(n1297_1),.b(n1300_1),.q(n1382));
  and_bi g170(.a(n168_0),.b(n169),.q(n170));
  bfr _b_6789(.a(_w_8691),.q(_w_8692));
  bfr _b_9194(.a(_w_11096),.q(_w_11097));
  spl2 g468_s_0(.a(n468),.q0(n468_0),.q1(n468_1));
  and_bb g1684(.a(N256_11),.b(N426_19),.q(n1684));
  and_bi g1419(.a(n1418_0),.b(n1373_0),.q(n1419));
  bfr _b_5063(.a(_w_6965),.q(N103_2));
  bfr _b_6403(.a(_w_8305),.q(_w_8306));
  bfr _b_4848(.a(_w_6750),.q(_w_6751));
  bfr _b_3859(.a(_w_5761),.q(_w_5762));
  bfr _b_5089(.a(_w_6991),.q(_w_6992));
  bfr _b_4964(.a(_w_6866),.q(_w_6867));
  bfr _b_3936(.a(_w_5838),.q(n78_1));
  and_bi g1461(.a(n1416_1),.b(n1419_1),.q(n1461));
  spl2 g914_s_0(.a(n914),.q0(n914_0),.q1(n914_1));
  spl2 g1057_s_0(.a(n1057),.q0(n1057_0),.q1(n1057_1));
  bfr _b_3435(.a(_w_5337),.q(_w_5338));
  bfr _b_5805(.a(_w_7707),.q(_w_7708));
  bfr _b_5158(.a(_w_7060),.q(_w_7061));
  and_bb g47(.a(n35_2),.b(n45_1),.q(_w_10838));
  bfr _b_4042(.a(_w_5944),.q(_w_5945));
  bfr _b_4084(.a(_w_5986),.q(_w_5987));
  and_bb g263(.a(n241_1),.b(n261_1),.q(_w_15310));
  bfr _b_9260(.a(_w_11162),.q(_w_11163));
  bfr _b_8759(.a(_w_10661),.q(n993));
  and_bi g373(.a(n318_1),.b(n321_1),.q(n373));
  bfr _b_4060(.a(_w_5962),.q(_w_5963));
  bfr _b_3682(.a(_w_5584),.q(_w_5585));
  or_bb g502(.a(n441_0),.b(n501_0),.q(n502));
  bfr _b_7290(.a(_w_9192),.q(_w_9193));
  spl2 g450_s_0(.a(n450),.q0(n450_0),.q1(n450_1));
  bfr _b_3626(.a(_w_5528),.q(_w_5529));
  and_bi g1285(.a(n1200_1),.b(n1203_1),.q(n1285));
  spl2 g486_s_0(.a(n486),.q0(n486_0),.q1(n486_1));
  and_bi g556(.a(n538_1),.b(n554_1),.q(_w_15311));
  bfr _b_3553(.a(_w_5455),.q(_w_5456));
  spl2 g1467_s_0(.a(n1467),.q0(n1467_0),.q1(n1467_1));
  bfr _b_13203(.a(_w_15105),.q(_w_15106));
  bfr _b_7995(.a(_w_9897),.q(_w_9898));
  spl2 g402_s_0(.a(n402),.q0(n402_0),.q1(n402_1));
  spl2 g1145_s_0(.a(n1145),.q0(n1145_0),.q1(n1145_1));
  bfr _b_3414(.a(_w_5316),.q(_w_5317));
  spl2 g474_s_0(.a(n474),.q0(n474_0),.q1(n474_1));
  bfr _b_5349(.a(_w_7251),.q(_w_7252));
  spl2 g901_s_0(.a(n901),.q0(n901_0),.q1(n901_1));
  spl2 g970_s_0(.a(n970),.q0(n970_0),.q1(n970_1));
  bfr _b_3904(.a(_w_5806),.q(_w_5807));
  and_bi g258(.a(n256_0),.b(n257),.q(n258));
  bfr _b_7227(.a(_w_9129),.q(n776));
  bfr _b_11273(.a(_w_13175),.q(_w_13176));
  spl4L N375_s_0(.a(_w_15596),.q0(N375_0),.q1(N375_1),.q2(N375_2),.q3(N375_3));
  spl2 g1505_s_0(.a(n1505),.q0(n1505_0),.q1(n1505_1));
  bfr _b_3826(.a(_w_5728),.q(_w_5729));
  bfr _b_4692(.a(_w_6594),.q(_w_6595));
  bfr _b_5797(.a(_w_7699),.q(_w_7700));
  and_bb g1834(.a(n1823_1),.b(n1832_1),.q(_w_15316));
  bfr _b_5755(.a(_w_7657),.q(_w_7658));
  bfr _b_6369(.a(_w_8271),.q(_w_8272));
  bfr _b_9708(.a(_w_11610),.q(_w_11611));
  bfr _b_3847(.a(_w_5749),.q(_w_5750));
  spl4L N375_s_1(.a(N375_0),.q0(N375_4),.q1(N375_5),.q2(N375_6),.q3(N375_7));
  bfr _b_10115(.a(_w_12017),.q(_w_12018));
  bfr _b_5068(.a(_w_6970),.q(_w_6971));
  bfr _b_4709(.a(_w_6611),.q(_w_6612));
  or_bb g51(.a(n49_0),.b(n50),.q(_w_11847));
  bfr _b_9656(.a(_w_11558),.q(_w_11559));
  spl2 g1774_s_0(.a(n1774),.q0(n1774_0),.q1(n1774_1));
  or_bb g1788(.a(n1786_0),.b(n1787_0),.q(n1788));
  spl2 g1876_s_0(.a(n1876),.q0(n1876_0),.q1(n1876_1));
  bfr _b_13475(.a(_w_15377),.q(_w_15378));
  spl2 g437_s_0(.a(n437),.q0(n437_0),.q1(n437_1));
  bfr _b_12435(.a(_w_14337),.q(_w_14338));
  spl2 g399_s_0(.a(n399),.q0(n399_0),.q1(n399_1));
  and_bi g1032(.a(n940_1),.b(n1030_1),.q(_w_9162));
  bfr _b_4647(.a(_w_6549),.q(_w_6550));
  spl2 g1646_s_0(.a(n1646),.q0(n1646_0),.q1(n1646_1));
  bfr _b_6632(.a(_w_8534),.q(_w_8535));
  spl2 g1819_s_0(.a(n1819),.q0(n1819_0),.q1(n1819_1));
  and_bi g326(.a(n324_0),.b(n325),.q(n326));
  bfr _b_4308(.a(_w_6210),.q(_w_6211));
  bfr _b_11580(.a(_w_13482),.q(_w_13483));
  or_bb g880(.a(n878_0),.b(n879),.q(n880));
  spl4L N18_s_0(.a(_w_15530),.q0(N18_0),.q1(_w_15317),.q2(_w_15341),.q3(_w_15397));
  spl2 g394_s_0(.a(n394),.q0(n394_0),.q1(_w_7267));
  spl2 g1280_s_0(.a(n1280),.q0(n1280_0),.q1(n1280_1));
  bfr _b_9204(.a(_w_11106),.q(n1608));
  spl2 g1560_s_0(.a(n1560),.q0(n1560_0),.q1(n1560_1));
  bfr _b_5038(.a(_w_6940),.q(_w_6941));
  bfr _b_6084(.a(_w_7986),.q(_w_7987));
  bfr _b_6734(.a(_w_8636),.q(_w_8637));
  bfr _b_4283(.a(_w_6185),.q(_w_6186));
  bfr _b_9376(.a(_w_11278),.q(_w_11279));
  spl2 g865_s_0(.a(n865),.q0(n865_0),.q1(n865_1));
  bfr _b_3589(.a(_w_5491),.q(_w_5492));
  and_bb g779(.a(n725_1),.b(n777_1),.q(_w_15521));
  bfr _b_8980(.a(_w_10882),.q(_w_10883));
  or_bb g687(.a(n685_0),.b(n686),.q(n687));
  and_bb g1705(.a(n1678_1),.b(n1703_1),.q(_w_14117));
  spl2 g1091_s_0(.a(n1091),.q0(n1091_0),.q1(n1091_1));
  spl2 g1103_s_0(.a(n1103),.q0(n1103_0),.q1(n1103_1));
  and_bb g620(.a(N426_8),.b(N69_13),.q(n620));
  bfr _b_6507(.a(_w_8409),.q(_w_8410));
  spl2 g295_s_0(.a(n295),.q0(n295_0),.q1(n295_1));
  and_bi g62(.a(n60_0),.b(n61),.q(n62));
  spl2 g376_s_0(.a(n376),.q0(n376_0),.q1(n376_1));
  bfr _b_5087(.a(_w_6989),.q(_w_6990));
  bfr _b_5085(.a(_w_6987),.q(_w_6988));
  bfr _b_5090(.a(_w_6992),.q(_w_6993));
  bfr _b_5091(.a(_w_6993),.q(_w_6994));
  and_bb g1492(.a(n1465_1),.b(n1490_1),.q(_w_13857));
  bfr _b_5094(.a(_w_6996),.q(_w_6997));
  bfr _b_7641(.a(_w_9543),.q(_w_9544));
  spl2 g1836_s_0(.a(n1836),.q0(n1836_0),.q1(n1836_1));
  bfr _b_5095(.a(_w_6997),.q(_w_6998));
  bfr _b_7899(.a(_w_9801),.q(_w_9802));
  bfr _b_5098(.a(_w_7000),.q(_w_7001));
  bfr _b_4057(.a(_w_5959),.q(_w_5960));
  or_bb g1479(.a(n1469_0),.b(n1478_0),.q(n1479));
  bfr _b_8147(.a(_w_10049),.q(_w_10050));
  bfr _b_13349(.a(_w_15251),.q(_w_15252));
  bfr _b_5099(.a(_w_7001),.q(_w_7002));
  bfr _b_5100(.a(_w_7002),.q(_w_7003));
  bfr _b_5101(.a(_w_7003),.q(_w_7004));
  bfr _b_5503(.a(_w_7405),.q(_w_7406));
  bfr _b_5103(.a(_w_7005),.q(_w_7006));
  bfr _b_3653(.a(_w_5555),.q(_w_5556));
  bfr _b_5104(.a(_w_7006),.q(_w_7007));
  bfr _b_7937(.a(_w_9839),.q(_w_9840));
  bfr _b_5105(.a(_w_7007),.q(_w_7008));
  or_bb g1415(.a(n1413_0),.b(n1414),.q(n1415));
  bfr _b_5615(.a(_w_7517),.q(_w_7518));
  bfr _b_5106(.a(_w_7008),.q(_w_7009));
  bfr _b_6276(.a(_w_8178),.q(N6230));
  bfr _b_5109(.a(_w_7011),.q(_w_7012));
  bfr _b_5113(.a(_w_7015),.q(_w_7016));
  or_bb g777(.a(n775_0),.b(n776),.q(n777));
  bfr _b_5114(.a(_w_7016),.q(_w_7017));
  bfr _b_3743(.a(_w_5645),.q(_w_5646));
  bfr _b_5117(.a(_w_7019),.q(_w_7020));
  bfr _b_5118(.a(_w_7020),.q(_w_7021));
  bfr _b_5120(.a(_w_7022),.q(_w_7023));
  bfr _b_5121(.a(_w_7023),.q(_w_7024));
  bfr _b_5398(.a(_w_7300),.q(_w_7301));
  bfr _b_13042(.a(_w_14944),.q(_w_14945));
  bfr _b_5122(.a(_w_7024),.q(_w_7025));
  bfr _b_4459(.a(_w_6361),.q(n150_1));
  bfr _b_7558(.a(_w_9460),.q(_w_9461));
  bfr _b_9844(.a(_w_11746),.q(_w_11747));
  bfr _b_8391(.a(_w_10293),.q(_w_10294));
  spl2 g965_s_0(.a(n965),.q0(n965_0),.q1(n965_1));
  bfr _b_5123(.a(_w_7025),.q(_w_7026));
  bfr _b_5124(.a(_w_7026),.q(_w_7027));
  bfr _b_5125(.a(_w_7027),.q(_w_7028));
  bfr _b_5126(.a(_w_7028),.q(_w_7029));
  bfr _b_5127(.a(_w_7029),.q(_w_7030));
  bfr _b_5128(.a(_w_7030),.q(_w_7031));
  bfr _b_13336(.a(_w_15238),.q(_w_15239));
  bfr _b_5131(.a(_w_7033),.q(_w_7034));
  bfr _b_5134(.a(_w_7036),.q(_w_7037));
  and_bb g1760(.a(n1733_1),.b(n1758_1),.q(_w_14570));
  bfr _b_5135(.a(_w_7037),.q(_w_7038));
  spl2 g1621_s_0(.a(n1621),.q0(n1621_0),.q1(n1621_1));
  bfr _b_5878(.a(_w_7780),.q(_w_7781));
  bfr _b_13435(.a(_w_15337),.q(_w_15338));
  bfr _b_13075(.a(_w_14977),.q(_w_14978));
  bfr _b_5138(.a(_w_7040),.q(_w_7041));
  bfr _b_6117(.a(_w_8019),.q(N205_11));
  bfr _b_5844(.a(_w_7746),.q(_w_7747));
  bfr _b_5956(.a(_w_7858),.q(_w_7859));
  bfr _b_11491(.a(_w_13393),.q(_w_13394));
  bfr _b_5140(.a(_w_7042),.q(_w_7043));
  bfr _b_5141(.a(_w_7043),.q(_w_7044));
  bfr _b_13469(.a(_w_15371),.q(_w_15372));
  bfr _b_11057(.a(_w_12959),.q(_w_12960));
  and_bi g843(.a(n748_1),.b(n751_1),.q(n843));
  and_bi g1018(.a(n1016_0),.b(n1017),.q(n1018));
  bfr _b_5142(.a(_w_7044),.q(_w_7045));
  and_bb g1435(.a(n1368_1),.b(n1433_1),.q(_w_13750));
  bfr _b_5143(.a(_w_7045),.q(_w_7046));
  bfr _b_5145(.a(_w_7047),.q(_w_7048));
  bfr _b_5146(.a(_w_7048),.q(_w_7049));
  bfr _b_5148(.a(_w_7050),.q(_w_7051));
  bfr _b_9717(.a(_w_11619),.q(n428));
  bfr _b_5149(.a(_w_7051),.q(_w_7052));
  bfr _b_11092(.a(_w_12994),.q(_w_12995));
  bfr _b_5152(.a(_w_7054),.q(_w_7055));
  bfr _b_3976(.a(_w_5878),.q(_w_5879));
  bfr _b_5153(.a(_w_7055),.q(_w_7056));
  bfr _b_5155(.a(_w_7057),.q(n208_1));
  bfr _b_5161(.a(_w_7063),.q(_w_7064));
  bfr _b_5165(.a(_w_7067),.q(_w_7068));
  bfr _b_5166(.a(_w_7068),.q(_w_7069));
  and_bi g696(.a(n694_0),.b(n695),.q(n696));
  bfr _b_5167(.a(_w_7069),.q(_w_7070));
  bfr _b_5168(.a(_w_7070),.q(_w_7071));
  bfr _b_8262(.a(_w_10164),.q(_w_10165));
  bfr _b_5171(.a(_w_7073),.q(_w_7074));
  bfr _b_7870(.a(_w_9772),.q(_w_9773));
  or_bb g394(.a(n373_0),.b(n393_0),.q(n394));
  bfr _b_5174(.a(_w_7076),.q(_w_7077));
  bfr _b_3751(.a(_w_5653),.q(_w_5654));
  bfr _b_7570(.a(_w_9472),.q(_w_9473));
  bfr _b_5175(.a(_w_7077),.q(_w_7078));
  bfr _b_10450(.a(_w_12352),.q(_w_12353));
  bfr _b_8045(.a(_w_9947),.q(n1871));
  spl2 g436_s_0(.a(n436),.q0(n436_0),.q1(n436_1));
  bfr _b_5176(.a(_w_7078),.q(_w_7079));
  bfr _b_5179(.a(_w_7081),.q(_w_7082));
  bfr _b_5180(.a(_w_7082),.q(_w_7083));
  bfr _b_5183(.a(_w_7085),.q(_w_7086));
  bfr _b_5184(.a(_w_7086),.q(_w_7087));
  bfr _b_10119(.a(_w_12021),.q(_w_12022));
  bfr _b_8269(.a(_w_10171),.q(_w_10172));
  and_bi g1275(.a(n1230_1),.b(n1233_1),.q(n1275));
  bfr _b_5891(.a(_w_7793),.q(_w_7794));
  bfr _b_5188(.a(_w_7090),.q(_w_7091));
  bfr _b_11453(.a(_w_13355),.q(_w_13356));
  bfr _b_5190(.a(_w_7092),.q(_w_7093));
  bfr _b_6668(.a(_w_8570),.q(_w_8571));
  bfr _b_5192(.a(_w_7094),.q(_w_7095));
  bfr _b_5194(.a(_w_7096),.q(_w_7097));
  bfr _b_10143(.a(_w_12045),.q(_w_12046));
  bfr _b_5196(.a(_w_7098),.q(_w_7099));
  bfr _b_9834(.a(_w_11736),.q(_w_11737));
  bfr _b_5198(.a(_w_7100),.q(_w_7101));
  bfr _b_5199(.a(_w_7101),.q(_w_7102));
  bfr _b_5200(.a(_w_7102),.q(_w_7103));
  and_bi g1854(.a(n1833_1),.b(n1836_1),.q(n1854));
  and_bi g445(.a(n406_1),.b(n409_1),.q(n445));
  bfr _b_5201(.a(_w_7103),.q(_w_7104));
  bfr _b_9180(.a(_w_11082),.q(n900));
  bfr _b_5203(.a(_w_7105),.q(_w_7106));
  bfr _b_5204(.a(_w_7106),.q(_w_7107));
  bfr _b_4923(.a(_w_6825),.q(_w_6826));
  bfr _b_5205(.a(_w_7107),.q(_w_7108));
  bfr _b_5207(.a(_w_7109),.q(_w_7110));
  bfr _b_5209(.a(_w_7111),.q(_w_7112));
  bfr _b_5211(.a(_w_7113),.q(_w_7114));
  bfr _b_6475(.a(_w_8377),.q(_w_8378));
  bfr _b_8538(.a(_w_10440),.q(n175));
  bfr _b_8674(.a(_w_10576),.q(_w_10577));
  bfr _b_8527(.a(_w_10429),.q(_w_10430));
  bfr _b_3472(.a(_w_5374),.q(_w_5375));
  and_bi g127(.a(n126_0),.b(n102_0),.q(n127));
  bfr _b_7984(.a(_w_9886),.q(_w_9887));
  bfr _b_5214(.a(_w_7116),.q(_w_7117));
  bfr _b_5215(.a(_w_7117),.q(_w_7118));
  bfr _b_13860(.a(_w_15762),.q(_w_15763));
  bfr _b_10900(.a(_w_12802),.q(_w_12803));
  bfr _b_8534(.a(_w_10436),.q(_w_10437));
  bfr _b_11119(.a(_w_13021),.q(_w_13022));
  bfr _b_4452(.a(_w_6354),.q(_w_6355));
  bfr _b_8950(.a(_w_10852),.q(_w_10853));
  bfr _b_8982(.a(_w_10884),.q(n500));
  bfr _b_5216(.a(_w_7118),.q(_w_7119));
  bfr _b_5219(.a(_w_7121),.q(_w_7122));
  or_bb g611(.a(n609_0),.b(n610),.q(_w_12736));
  bfr _b_5220(.a(_w_7122),.q(_w_7123));
  bfr _b_5224(.a(_w_7126),.q(_w_7127));
  bfr _b_12877(.a(_w_14779),.q(_w_14780));
  bfr _b_5225(.a(_w_7127),.q(_w_7128));
  bfr _b_9753(.a(_w_11655),.q(_w_11656));
  bfr _b_6886(.a(_w_8788),.q(n88_1));
  bfr _b_5229(.a(_w_7131),.q(_w_7132));
  bfr _b_6365(.a(_w_8267),.q(_w_8268));
  bfr _b_7773(.a(_w_9675),.q(_w_9676));
  bfr _b_6904(.a(_w_8806),.q(n844));
  bfr _b_5231(.a(_w_7133),.q(_w_7134));
  bfr _b_5232(.a(_w_7134),.q(_w_7135));
  bfr _b_7023(.a(_w_8925),.q(n1243));
  bfr _b_5233(.a(_w_7135),.q(_w_7136));
  bfr _b_5235(.a(_w_7137),.q(_w_7138));
  and_bi g1544(.a(n1491_1),.b(n1494_1),.q(n1544));
  bfr _b_5240(.a(_w_7142),.q(_w_7143));
  bfr _b_6028(.a(_w_7930),.q(_w_7931));
  bfr _b_3926(.a(_w_5828),.q(_w_5829));
  bfr _b_7193(.a(_w_9095),.q(_w_9096));
  bfr _b_5243(.a(_w_7145),.q(_w_7146));
  bfr _b_5992(.a(_w_7894),.q(_w_7895));
  spl2 g123_s_0(.a(n123),.q0(n123_0),.q1(n123_1));
  bfr _b_9941(.a(_w_11843),.q(_w_11844));
  bfr _b_13693(.a(_w_15595),.q(_w_15571));
  and_bi g1831(.a(n1824_1),.b(n1829_1),.q(_w_14571));
  bfr _b_5246(.a(_w_7148),.q(_w_7149));
  bfr _b_5282(.a(_w_7184),.q(_w_7185));
  and_bi g441(.a(n418_1),.b(n421_1),.q(n441));
  bfr _b_5247(.a(_w_7149),.q(_w_7150));
  or_bb g1297(.a(n1287_0),.b(n1296_0),.q(n1297));
  bfr _b_10142(.a(_w_12044),.q(_w_12045));
  bfr _b_5353(.a(_w_7255),.q(_w_7256));
  or_bb g911(.a(n827_0),.b(n910_0),.q(n911));
  bfr _b_7666(.a(_w_9568),.q(_w_9569));
  bfr _b_4105(.a(_w_6007),.q(_w_6008));
  bfr _b_5249(.a(_w_7151),.q(_w_7152));
  and_bb g820(.a(N1_19),.b(N528_4),.q(_w_8809));
  and_bb g1173(.a(N137_14),.b(N443_12),.q(_w_12080));
  bfr _b_5250(.a(_w_7152),.q(_w_7153));
  and_bb g442(.a(N409_7),.b(N52_12),.q(n442));
  bfr _b_5251(.a(_w_7153),.q(_w_7154));
  bfr _b_7120(.a(_w_9022),.q(_w_9023));
  bfr _b_5252(.a(_w_7154),.q(_w_7155));
  bfr _b_14001(.a(_w_15903),.q(_w_15904));
  bfr _b_10135(.a(_w_12037),.q(_w_12038));
  bfr _b_7342(.a(_w_9244),.q(n194));
  bfr _b_5253(.a(_w_7155),.q(_w_7156));
  bfr _b_12530(.a(_w_14432),.q(_w_14433));
  bfr _b_8020(.a(_w_9922),.q(_w_9923));
  bfr _b_5254(.a(_w_7156),.q(_w_7157));
  bfr _b_9484(.a(_w_11386),.q(_w_11387));
  bfr _b_10813(.a(_w_12715),.q(_w_12716));
  bfr _b_5256(.a(_w_7158),.q(_w_7159));
  bfr _b_5257(.a(_w_7159),.q(_w_7160));
  bfr _b_11116(.a(_w_13018),.q(_w_13019));
  bfr _b_8628(.a(_w_10530),.q(_w_10531));
  bfr _b_5259(.a(_w_7161),.q(_w_7162));
  bfr _b_5260(.a(_w_7162),.q(_w_7163));
  bfr _b_12714(.a(_w_14616),.q(_w_14617));
  bfr _b_5262(.a(_w_7164),.q(_w_7165));
  bfr _b_8399(.a(_w_10301),.q(_w_10302));
  bfr _b_6095(.a(_w_7997),.q(_w_7998));
  and_bb g269(.a(n239_1),.b(n267_1),.q(_w_12856));
  bfr _b_5264(.a(_w_7166),.q(_w_7167));
  bfr _b_5265(.a(_w_7167),.q(_w_7168));
  spl2 g1698_s_0(.a(n1698),.q0(n1698_0),.q1(_w_5539));
  bfr _b_7310(.a(_w_9212),.q(_w_9213));
  spl2 g1283_s_0(.a(n1283),.q0(n1283_0),.q1(n1283_1));
  bfr _b_5266(.a(_w_7168),.q(_w_7169));
  bfr _b_4214(.a(_w_6116),.q(_w_6117));
  bfr _b_5267(.a(_w_7169),.q(_w_7170));
  bfr _b_5268(.a(_w_7170),.q(_w_7171));
  bfr _b_8434(.a(_w_10336),.q(_w_10337));
  bfr _b_5269(.a(_w_7171),.q(_w_7172));
  bfr _b_5270(.a(_w_7172),.q(_w_7173));
  bfr _b_6168(.a(_w_8070),.q(_w_8071));
  and_bi g1443(.a(n1442_0),.b(n1365_0),.q(n1443));
  bfr _b_5271(.a(_w_7173),.q(_w_7174));
  bfr _b_5272(.a(_w_7174),.q(_w_7175));
  bfr _b_6684(.a(_w_8586),.q(_w_8587));
  bfr _b_8094(.a(_w_9996),.q(_w_9997));
  bfr _b_8166(.a(_w_10068),.q(_w_10069));
  bfr _b_8194(.a(_w_10096),.q(_w_10097));
  bfr _b_5277(.a(_w_7179),.q(_w_7180));
  bfr _b_5280(.a(_w_7182),.q(_w_7183));
  bfr _b_6050(.a(_w_7952),.q(_w_7953));
  bfr _b_5281(.a(_w_7183),.q(_w_7184));
  bfr _b_5283(.a(_w_7185),.q(_w_7186));
  bfr _b_8876(.a(_w_10778),.q(n169));
  bfr _b_5285(.a(_w_7187),.q(_w_7188));
  bfr _b_5286(.a(_w_7188),.q(_w_7189));
  bfr _b_7208(.a(_w_9110),.q(_w_9111));
  bfr _b_5288(.a(_w_7190),.q(_w_7191));
  bfr _b_5290(.a(_w_7192),.q(_w_7193));
  bfr _b_6213(.a(_w_8115),.q(_w_8116));
  bfr _b_5291(.a(_w_7193),.q(_w_7194));
  bfr _b_5293(.a(_w_7195),.q(_w_7196));
  bfr _b_8681(.a(_w_10583),.q(_w_10584));
  bfr _b_5295(.a(_w_7197),.q(_w_7198));
  bfr _b_5296(.a(_w_7198),.q(_w_7199));
  bfr _b_11110(.a(_w_13012),.q(n1246));
  bfr _b_5173(.a(_w_7075),.q(_w_7076));
  bfr _b_5298(.a(_w_7200),.q(_w_7201));
  bfr _b_5299(.a(_w_7201),.q(_w_7202));
  bfr _b_5302(.a(_w_7204),.q(_w_7205));
  bfr _b_5304(.a(_w_7206),.q(_w_7207));
  bfr _b_7602(.a(_w_9504),.q(_w_9505));
  bfr _b_3830(.a(_w_5732),.q(_w_5733));
  bfr _b_5305(.a(_w_7207),.q(_w_7208));
  spl2 g344_s_0(.a(n344),.q0(n344_0),.q1(n344_1));
  bfr _b_5309(.a(_w_7211),.q(_w_7212));
  bfr _b_8346(.a(_w_10248),.q(_w_10249));
  bfr _b_9363(.a(_w_11265),.q(_w_11266));
  bfr _b_5311(.a(_w_7213),.q(_w_7214));
  and_bi g1426(.a(n1371_1),.b(n1424_1),.q(_w_13583));
  bfr _b_5314(.a(_w_7216),.q(_w_7217));
  bfr _b_5315(.a(_w_7217),.q(_w_7218));
  bfr _b_5318(.a(_w_7220),.q(_w_7221));
  bfr _b_12082(.a(_w_13984),.q(n1657));
  bfr _b_5319(.a(_w_7221),.q(_w_7222));
  bfr _b_13740(.a(_w_15642),.q(_w_15643));
  bfr _b_13575(.a(_w_15477),.q(_w_15478));
  bfr _b_3608(.a(_w_5510),.q(_w_5511));
  bfr _b_8506(.a(_w_10408),.q(_w_10409));
  bfr _b_7922(.a(_w_9824),.q(_w_9825));
  bfr _b_11427(.a(_w_13329),.q(_w_13330));
  bfr _b_5323(.a(_w_7225),.q(_w_7226));
  bfr _b_8748(.a(_w_10650),.q(_w_10651));
  bfr _b_5327(.a(_w_7229),.q(_w_7230));
  bfr _b_5329(.a(_w_7231),.q(_w_7232));
  bfr _b_5092(.a(_w_6994),.q(_w_6995));
  bfr _b_5330(.a(_w_7232),.q(_w_7233));
  bfr _b_4361(.a(_w_6263),.q(_w_6264));
  bfr _b_5333(.a(_w_7235),.q(_w_7236));
  bfr _b_13790(.a(_w_15692),.q(_w_15693));
  bfr _b_5334(.a(_w_7236),.q(_w_7237));
  bfr _b_11943(.a(_w_13845),.q(_w_13846));
  bfr _b_9960(.a(_w_11862),.q(_w_11863));
  bfr _b_5336(.a(_w_7238),.q(_w_7239));
  bfr _b_5337(.a(_w_7239),.q(_w_7240));
  bfr _b_9035(.a(_w_10937),.q(_w_10938));
  bfr _b_8097(.a(_w_9999),.q(_w_10000));
  bfr _b_5338(.a(_w_7240),.q(_w_7241));
  bfr _b_6976(.a(_w_8878),.q(_w_8879));
  bfr _b_8070(.a(_w_9972),.q(n840));
  bfr _b_10193(.a(_w_12095),.q(n178));
  bfr _b_7685(.a(_w_9587),.q(n962_1));
  bfr _b_5339(.a(_w_7241),.q(_w_7242));
  bfr _b_5340(.a(_w_7242),.q(_w_7243));
  bfr _b_5341(.a(_w_7243),.q(_w_7244));
  bfr _b_7363(.a(_w_9265),.q(_w_9266));
  bfr _b_9350(.a(_w_11252),.q(_w_11253));
  bfr _b_5346(.a(_w_7248),.q(_w_7249));
  bfr _b_5863(.a(_w_7765),.q(_w_7766));
  bfr _b_8585(.a(_w_10487),.q(_w_10488));
  bfr _b_5348(.a(_w_7250),.q(_w_7251));
  bfr _b_8431(.a(_w_10333),.q(_w_10334));
  or_bb g759(.a(n757_0),.b(n758),.q(n759));
  bfr _b_7879(.a(_w_9781),.q(_w_9782));
  bfr _b_8825(.a(_w_10727),.q(_w_10728));
  bfr _b_6362(.a(_w_8264),.q(_w_8265));
  bfr _b_5352(.a(_w_7254),.q(_w_7255));
  bfr _b_5354(.a(_w_7256),.q(_w_7257));
  bfr _b_13130(.a(_w_15032),.q(_w_15033));
  spl4L N494_s_3(.a(N494_2),.q0(N494_12),.q1(N494_13),.q2(N494_14),.q3(N494_15));
  bfr _b_5136(.a(_w_7038),.q(_w_7039));
  bfr _b_5356(.a(_w_7258),.q(N35_11));
  bfr _b_5191(.a(_w_7093),.q(_w_7094));
  bfr _b_5357(.a(_w_7259),.q(_w_7260));
  bfr _b_5358(.a(_w_7260),.q(N35_6));
  bfr _b_7270(.a(_w_9172),.q(_w_9173));
  bfr _b_5359(.a(_w_7261),.q(_w_7262));
  bfr _b_5360(.a(_w_7262),.q(N35_7));
  bfr _b_5361(.a(_w_7263),.q(_w_7264));
  bfr _b_9185(.a(_w_11087),.q(_w_11088));
  bfr _b_5362(.a(_w_7264),.q(_w_7265));
  bfr _b_5738(.a(_w_7640),.q(_w_7641));
  and_bb g1371(.a(N137_16),.b(N477_12),.q(n1371));
  bfr _b_5364(.a(_w_7266),.q(n1759_1));
  bfr _b_3801(.a(_w_5703),.q(_w_5704));
  bfr _b_5365(.a(_w_7267),.q(_w_7268));
  bfr _b_11246(.a(_w_13148),.q(n1681));
  bfr _b_7427(.a(_w_9329),.q(_w_9330));
  bfr _b_5366(.a(_w_7268),.q(_w_7269));
  bfr _b_10198(.a(_w_12100),.q(_w_12101));
  bfr _b_5368(.a(_w_7270),.q(n394_1));
  bfr _b_5369(.a(_w_7271),.q(_w_7272));
  bfr _b_7788(.a(_w_9690),.q(_w_9691));
  bfr _b_5370(.a(_w_7272),.q(_w_7273));
  bfr _b_12386(.a(_w_14288),.q(n940));
  bfr _b_5372(.a(_w_7274),.q(_w_7275));
  bfr _b_5927(.a(_w_7829),.q(_w_7830));
  and_bi g1617(.a(n1564_1),.b(n1567_1),.q(n1617));
  bfr _b_5376(.a(_w_7278),.q(_w_7279));
  bfr _b_9724(.a(_w_11626),.q(_w_11627));
  bfr _b_5377(.a(_w_7279),.q(_w_7280));
  bfr _b_7353(.a(_w_9255),.q(_w_9256));
  bfr _b_5384(.a(_w_7286),.q(_w_7287));
  and_bb g785(.a(n723_1),.b(n783_1),.q(_w_10451));
  and_bi g235(.a(n220_1),.b(n223_1),.q(n235));
  bfr _b_8420(.a(_w_10322),.q(_w_10323));
  bfr _b_5385(.a(_w_7287),.q(_w_7288));
  bfr _b_6467(.a(_w_8369),.q(n1207));
  bfr _b_5387(.a(_w_7289),.q(_w_7290));
  bfr _b_5389(.a(_w_7291),.q(_w_7292));
  bfr _b_5391(.a(_w_7293),.q(_w_7294));
  bfr _b_7655(.a(_w_9557),.q(_w_9558));
  bfr _b_9925(.a(_w_11827),.q(_w_11828));
  bfr _b_5392(.a(_w_7294),.q(N86_11));
  bfr _b_10580(.a(_w_12482),.q(_w_12483));
  bfr _b_9936(.a(_w_11838),.q(_w_11839));
  bfr _b_5393(.a(_w_7295),.q(_w_7296));
  bfr _b_5396(.a(_w_7298),.q(_w_7299));
  bfr _b_5397(.a(_w_7299),.q(_w_7300));
  bfr _b_8213(.a(_w_10115),.q(_w_10116));
  bfr _b_4536(.a(_w_6438),.q(_w_6439));
  bfr _b_4373(.a(_w_6275),.q(n640_1));
  bfr _b_7482(.a(_w_9384),.q(_w_9385));
  bfr _b_5400(.a(_w_7302),.q(_w_7303));
  and_bi g662(.a(n628_1),.b(n660_1),.q(_w_9247));
  bfr _b_5342(.a(_w_7244),.q(_w_7245));
  bfr _b_5401(.a(_w_7303),.q(_w_7304));
  bfr _b_5404(.a(_w_7306),.q(_w_7307));
  bfr _b_5405(.a(_w_7307),.q(_w_7308));
  bfr _b_5406(.a(_w_7308),.q(_w_7309));
  bfr _b_7651(.a(_w_9553),.q(_w_9554));
  bfr _b_7780(.a(_w_9682),.q(_w_9683));
  bfr _b_5409(.a(_w_7311),.q(_w_7312));
  bfr _b_6173(.a(_w_8075),.q(_w_8076));
  bfr _b_11276(.a(_w_13178),.q(_w_13179));
  bfr _b_5410(.a(_w_7312),.q(_w_7313));
  bfr _b_6077(.a(_w_7979),.q(_w_7980));
  bfr _b_5414(.a(_w_7316),.q(_w_7317));
  bfr _b_5417(.a(_w_7319),.q(_w_7320));
  bfr _b_6292(.a(_w_8194),.q(_w_8195));
  bfr _b_5418(.a(_w_7320),.q(_w_7321));
  bfr _b_5421(.a(_w_7323),.q(_w_7324));
  bfr _b_5422(.a(_w_7324),.q(_w_7325));
  bfr _b_4426(.a(_w_6328),.q(n600_1));
  bfr _b_5425(.a(_w_7327),.q(_w_7328));
  bfr _b_5426(.a(_w_7328),.q(_w_7329));
  bfr _b_9706(.a(_w_11608),.q(_w_11609));
  bfr _b_5430(.a(_w_7332),.q(_w_7333));
  bfr _b_5431(.a(_w_7333),.q(_w_7334));
  bfr _b_4937(.a(_w_6839),.q(_w_6840));
  bfr _b_3464(.a(_w_5366),.q(_w_5367));
  bfr _b_8724(.a(_w_10626),.q(n1038));
  bfr _b_12832(.a(_w_14734),.q(_w_14735));
  bfr _b_3725(.a(_w_5627),.q(_w_5628));
  bfr _b_5434(.a(_w_7336),.q(_w_7337));
  bfr _b_11428(.a(_w_13330),.q(_w_13331));
  or_bb g458(.a(n377_1),.b(n457_0),.q(_w_12486));
  bfr _b_6287(.a(_w_8189),.q(_w_8190));
  bfr _b_7008(.a(_w_8910),.q(_w_8911));
  bfr _b_3775(.a(_w_5677),.q(_w_5678));
  bfr _b_5435(.a(_w_7337),.q(_w_7338));
  bfr _b_12219(.a(_w_14121),.q(n1582_1));
  or_bb g1315(.a(n1281_0),.b(n1314_0),.q(n1315));
  bfr _b_5436(.a(_w_7338),.q(_w_7339));
  bfr _b_5438(.a(_w_7340),.q(_w_7341));
  bfr _b_5440(.a(_w_7342),.q(_w_7343));
  bfr _b_5441(.a(_w_7343),.q(_w_7344));
  bfr _b_4802(.a(_w_6704),.q(_w_6705));
  bfr _b_5217(.a(_w_7119),.q(_w_7120));
  bfr _b_5442(.a(_w_7344),.q(_w_7345));
  bfr _b_5443(.a(_w_7345),.q(_w_7346));
  bfr _b_4640(.a(_w_6542),.q(_w_6543));
  bfr _b_5445(.a(_w_7347),.q(_w_7348));
  bfr _b_7354(.a(_w_9256),.q(n1710_1));
  and_bi g517(.a(n516_0),.b(n436_0),.q(n517));
  spl2 g951_s_0(.a(n951),.q0(n951_0),.q1(n951_1));
  bfr _b_8134(.a(_w_10036),.q(_w_10037));
  bfr _b_5447(.a(_w_7349),.q(_w_7350));
  bfr _b_9791(.a(_w_11693),.q(_w_11694));
  or_bb g998(.a(n951_0),.b(n997_0),.q(n998));
  bfr _b_5448(.a(_w_7350),.q(_w_7351));
  bfr _b_5449(.a(_w_7351),.q(_w_7352));
  bfr _b_5451(.a(_w_7353),.q(_w_7354));
  bfr _b_9482(.a(_w_11384),.q(_w_11385));
  bfr _b_5453(.a(_w_7355),.q(_w_7356));
  bfr _b_11422(.a(_w_13324),.q(_w_13325));
  bfr _b_7127(.a(_w_9029),.q(_w_9030));
  spl2 g356_s_0(.a(n356),.q0(n356_0),.q1(n356_1));
  bfr _b_5455(.a(_w_7357),.q(_w_7358));
  spl2 g400_s_0(.a(n400),.q0(n400_0),.q1(_w_7543));
  bfr _b_7253(.a(_w_9155),.q(_w_9156));
  and_bb g1734(.a(N205_17),.b(N494_16),.q(_w_14218));
  bfr _b_5456(.a(_w_7358),.q(_w_7359));
  bfr _b_4823(.a(_w_6725),.q(_w_6726));
  and_bi g585(.a(n584_0),.b(n528_0),.q(n585));
  bfr _b_5459(.a(_w_7361),.q(_w_7362));
  bfr _b_5460(.a(_w_7362),.q(_w_7363));
  bfr _b_7522(.a(_w_9424),.q(_w_9425));
  bfr _b_5462(.a(_w_7364),.q(_w_7365));
  bfr _b_9479(.a(_w_11381),.q(_w_11382));
  bfr _b_5464(.a(_w_7366),.q(_w_7367));
  bfr _b_5465(.a(_w_7367),.q(_w_7368));
  bfr _b_10010(.a(_w_11912),.q(_w_11913));
  bfr _b_5466(.a(_w_7368),.q(_w_7369));
  bfr _b_5467(.a(_w_7369),.q(_w_7370));
  bfr _b_12633(.a(_w_14535),.q(_w_14536));
  bfr _b_3868(.a(_w_5770),.q(_w_5771));
  bfr _b_5468(.a(_w_7370),.q(_w_7371));
  bfr _b_10055(.a(_w_11957),.q(_w_11958));
  bfr _b_5472(.a(_w_7374),.q(N86_2));
  bfr _b_11232(.a(_w_13134),.q(_w_13135));
  bfr _b_3932(.a(_w_5834),.q(n974_1));
  bfr _b_5473(.a(_w_7375),.q(_w_7376));
  bfr _b_5476(.a(_w_7378),.q(_w_7379));
  bfr _b_9512(.a(_w_11414),.q(_w_11415));
  bfr _b_5953(.a(_w_7855),.q(_w_7856));
  bfr _b_5477(.a(_w_7379),.q(_w_7380));
  bfr _b_5478(.a(_w_7380),.q(_w_7381));
  bfr _b_7107(.a(_w_9009),.q(_w_9010));
  bfr _b_3732(.a(_w_5634),.q(_w_5635));
  bfr _b_3547(.a(_w_5449),.q(_w_5450));
  bfr _b_5481(.a(_w_7383),.q(_w_7384));
  spl2 g1647_s_0(.a(n1647),.q0(n1647_0),.q1(_w_10885));
  bfr _b_10240(.a(_w_12142),.q(_w_12143));
  bfr _b_5482(.a(_w_7384),.q(_w_7385));
  bfr _b_7171(.a(_w_9073),.q(_w_9074));
  bfr _b_12416(.a(_w_14318),.q(_w_14319));
  bfr _b_10102(.a(_w_12004),.q(_w_12005));
  bfr _b_13627(.a(N171),.q(_w_15529));
  bfr _b_5483(.a(_w_7385),.q(_w_7386));
  bfr _b_4023(.a(_w_5925),.q(_w_5926));
  bfr _b_5485(.a(_w_7387),.q(_w_7388));
  bfr _b_5044(.a(_w_6946),.q(_w_6947));
  bfr _b_5486(.a(_w_7388),.q(_w_7389));
  bfr _b_5487(.a(_w_7389),.q(_w_7390));
  bfr _b_7929(.a(_w_9831),.q(_w_9832));
  bfr _b_9189(.a(_w_11091),.q(_w_11092));
  bfr _b_5494(.a(_w_7396),.q(_w_7397));
  bfr _b_7938(.a(_w_9840),.q(_w_9841));
  bfr _b_8196(.a(_w_10098),.q(_w_10099));
  bfr _b_5495(.a(_w_7397),.q(_w_7398));
  bfr _b_8447(.a(_w_10349),.q(_w_10350));
  bfr _b_5496(.a(_w_7398),.q(_w_7399));
  bfr _b_5497(.a(_w_7399),.q(_w_7400));
  bfr _b_5501(.a(_w_7403),.q(_w_7404));
  bfr _b_5502(.a(_w_7404),.q(_w_7405));
  bfr _b_5504(.a(_w_7406),.q(_w_7407));
  bfr _b_6184(.a(_w_8086),.q(_w_8087));
  bfr _b_5505(.a(_w_7407),.q(_w_7408));
  bfr _b_5507(.a(_w_7409),.q(_w_7410));
  bfr _b_5508(.a(_w_7410),.q(_w_7411));
  bfr _b_11449(.a(_w_13351),.q(_w_13352));
  bfr _b_5511(.a(_w_7413),.q(_w_7414));
  spl2 g905_s_0(.a(n905),.q0(n905_0),.q1(_w_5849));
  bfr _b_6079(.a(_w_7981),.q(_w_7982));
  bfr _b_8860(.a(_w_10762),.q(_w_10763));
  bfr _b_7969(.a(_w_9871),.q(_w_9872));
  and_bi g1152(.a(n1151_0),.b(n1050_0),.q(n1152));
  bfr _b_5512(.a(_w_7414),.q(_w_7415));
  bfr _b_5513(.a(_w_7415),.q(_w_7416));
  bfr _b_7220(.a(_w_9122),.q(_w_9123));
  bfr _b_10461(.a(_w_12363),.q(n1333_1));
  bfr _b_5514(.a(_w_7416),.q(_w_7417));
  bfr _b_5939(.a(_w_7841),.q(_w_7842));
  bfr _b_8937(.a(_w_10839),.q(_w_10840));
  bfr _b_5523(.a(_w_7425),.q(_w_7426));
  bfr _b_5525(.a(_w_7427),.q(_w_7428));
  bfr _b_4329(.a(_w_6231),.q(N120_14));
  bfr _b_9913(.a(_w_11815),.q(n1483));
  and_bi g1158(.a(n1157_0),.b(n1046_1),.q(n1158));
  bfr _b_5526(.a(_w_7428),.q(_w_7429));
  bfr _b_8955(.a(_w_10857),.q(_w_10858));
  bfr _b_5528(.a(_w_7430),.q(_w_7431));
  spl2 g186_s_0(.a(n186),.q0(n186_0),.q1(n186_1));
  bfr _b_5530(.a(_w_7432),.q(_w_7433));
  bfr _b_11693(.a(_w_13595),.q(_w_13596));
  bfr _b_9452(.a(_w_11354),.q(_w_11355));
  bfr _b_12703(.a(_w_14605),.q(_w_14606));
  bfr _b_5531(.a(_w_7433),.q(_w_7434));
  and_bb g1543(.a(N188_15),.b(N460_15),.q(_w_11146));
  bfr _b_5532(.a(_w_7434),.q(_w_7435));
  bfr _b_5534(.a(_w_7436),.q(_w_7437));
  bfr _b_5536(.a(_w_7438),.q(_w_7439));
  bfr _b_5537(.a(_w_7439),.q(_w_7440));
  bfr _b_5538(.a(_w_7440),.q(_w_7441));
  bfr _b_12037(.a(_w_13939),.q(n644));
  bfr _b_5540(.a(_w_7442),.q(_w_7443));
  bfr _b_8468(.a(_w_10370),.q(_w_10371));
  bfr _b_6552(.a(_w_8454),.q(_w_8455));
  bfr _b_5541(.a(_w_7443),.q(_w_7444));
  spl2 g1367_s_0(.a(n1367),.q0(n1367_0),.q1(n1367_1));
  bfr _b_6035(.a(_w_7937),.q(_w_7938));
  bfr _b_6702(.a(_w_8604),.q(_w_8605));
  bfr _b_5543(.a(_w_7445),.q(_w_7446));
  bfr _b_5544(.a(_w_7446),.q(_w_7447));
  bfr _b_8336(.a(_w_10238),.q(_w_10239));
  bfr _b_5545(.a(_w_7447),.q(_w_7448));
  bfr _b_8670(.a(_w_10572),.q(n855));
  and_bi g487(.a(n486_0),.b(n446_0),.q(n487));
  bfr _b_5546(.a(_w_7448),.q(_w_7449));
  bfr _b_8305(.a(_w_10207),.q(_w_10208));
  bfr _b_5548(.a(_w_7450),.q(_w_7451));
  spl2 g387_s_0(.a(n387),.q0(n387_0),.q1(n387_1));
  bfr _b_5549(.a(_w_7451),.q(_w_7452));
  and_bi g1810(.a(n1779_1),.b(n1808_1),.q(_w_12079));
  bfr _b_5551(.a(_w_7453),.q(_w_7454));
  bfr _b_9358(.a(_w_11260),.q(_w_11261));
  bfr _b_5552(.a(_w_7454),.q(_w_7455));
  and_bb g1090(.a(n1071_1),.b(n1088_1),.q(_w_8201));
  or_bb g214(.a(n185_0),.b(n213_0),.q(n214));
  bfr _b_5553(.a(_w_7455),.q(_w_7456));
  bfr _b_8979(.a(_w_10881),.q(n316));
  bfr _b_12088(.a(_w_13990),.q(_w_13991));
  bfr _b_5557(.a(_w_7459),.q(_w_7460));
  bfr _b_5558(.a(_w_7460),.q(_w_7461));
  spl2 g988_s_0(.a(n988),.q0(n988_0),.q1(n988_1));
  bfr _b_7932(.a(_w_9834),.q(_w_9835));
  bfr _b_5560(.a(_w_7462),.q(N86_3));
  bfr _b_5564(.a(_w_7466),.q(n814_1));
  bfr _b_9186(.a(_w_11088),.q(_w_11089));
  bfr _b_5565(.a(_w_7467),.q(_w_7468));
  bfr _b_5566(.a(_w_7468),.q(_w_7469));
  bfr _b_10884(.a(_w_12786),.q(_w_12787));
  spl2 g769_s_0(.a(n769),.q0(n769_0),.q1(n769_1));
  bfr _b_5567(.a(_w_7469),.q(_w_7470));
  bfr _b_12727(.a(_w_14629),.q(_w_14630));
  bfr _b_5571(.a(_w_7473),.q(_w_7474));
  bfr _b_5825(.a(_w_7727),.q(_w_7728));
  bfr _b_5574(.a(_w_7476),.q(_w_7477));
  spl2 g1009_s_0(.a(n1009),.q0(n1009_0),.q1(n1009_1));
  bfr _b_5575(.a(_w_7477),.q(_w_7478));
  bfr _b_5578(.a(_w_7480),.q(_w_7481));
  and_bb g739(.a(N239_5),.b(N273_18),.q(_w_13003));
  bfr _b_5829(.a(_w_7731),.q(_w_7732));
  bfr _b_5579(.a(_w_7481),.q(_w_7482));
  bfr _b_5580(.a(_w_7482),.q(_w_7483));
  bfr _b_5582(.a(_w_7484),.q(_w_7485));
  bfr _b_5583(.a(_w_7485),.q(_w_7486));
  bfr _b_11487(.a(_w_13389),.q(_w_13390));
  bfr _b_4715(.a(_w_6617),.q(_w_6618));
  or_bb g640(.a(n542_1),.b(n639_0),.q(n640));
  bfr _b_8085(.a(_w_9987),.q(n74));
  bfr _b_9995(.a(_w_11897),.q(_w_11898));
  bfr _b_5591(.a(_w_7493),.q(_w_7494));
  bfr _b_5592(.a(_w_7494),.q(_w_7495));
  bfr _b_5394(.a(_w_7296),.q(_w_7297));
  bfr _b_5597(.a(_w_7499),.q(_w_7500));
  bfr _b_6478(.a(_w_8380),.q(n1054));
  bfr _b_5598(.a(_w_7500),.q(_w_7501));
  bfr _b_6196(.a(_w_8098),.q(_w_8099));
  bfr _b_5604(.a(_w_7506),.q(_w_7507));
  spl2 g1845_s_0(.a(n1845),.q0(n1845_0),.q1(_w_11624));
  bfr _b_5605(.a(_w_7507),.q(_w_7508));
  bfr _b_5607(.a(_w_7509),.q(_w_7510));
  bfr _b_5608(.a(_w_7510),.q(N69_15));
  bfr _b_5610(.a(_w_7512),.q(_w_7513));
  bfr _b_5611(.a(_w_7513),.q(_w_7514));
  bfr _b_7400(.a(_w_9302),.q(_w_9303));
  spl4L N103_s_1(.a(N103_0),.q0(N103_4),.q1(N103_5),.q2(_w_6882),.q3(_w_6884));
  bfr _b_5773(.a(_w_7675),.q(_w_7676));
  bfr _b_5613(.a(_w_7515),.q(_w_7516));
  bfr _b_3511(.a(_w_5413),.q(_w_5414));
  and_bi g572(.a(n570_0),.b(n571),.q(n572));
  bfr _b_5614(.a(_w_7516),.q(_w_7517));
  bfr _b_10974(.a(_w_12876),.q(_w_12877));
  bfr _b_5616(.a(_w_7518),.q(_w_7519));
  bfr _b_5617(.a(_w_7519),.q(_w_7520));
  bfr _b_5619(.a(_w_7521),.q(_w_7522));
  bfr _b_5623(.a(_w_7525),.q(_w_7526));
  bfr _b_5627(.a(_w_7529),.q(_w_7530));
  bfr _b_5524(.a(_w_7426),.q(_w_7427));
  bfr _b_5628(.a(_w_7530),.q(_w_7531));
  bfr _b_5629(.a(_w_7531),.q(_w_7532));
  bfr _b_8084(.a(_w_9986),.q(_w_9987));
  bfr _b_8505(.a(_w_10407),.q(_w_10408));
  bfr _b_5632(.a(_w_7534),.q(N69_11));
  or_bb g430(.a(n361_0),.b(n429_0),.q(n430));
  bfr _b_9434(.a(_w_11336),.q(_w_11337));
  bfr _b_5633(.a(_w_7535),.q(_w_7536));
  bfr _b_5635(.a(_w_7537),.q(_w_7538));
  bfr _b_8178(.a(_w_10080),.q(_w_10081));
  bfr _b_12048(.a(_w_13950),.q(n1586));
  spl2 g1178_s_0(.a(n1178),.q0(n1178_0),.q1(n1178_1));
  bfr _b_5638(.a(_w_7540),.q(_w_7541));
  bfr _b_3484(.a(_w_5386),.q(_w_5387));
  bfr _b_5640(.a(_w_7542),.q(n312_1));
  bfr _b_11926(.a(_w_13828),.q(_w_13829));
  bfr _b_5985(.a(_w_7887),.q(_w_7888));
  bfr _b_5641(.a(_w_7543),.q(_w_7544));
  bfr _b_12460(.a(_w_14362),.q(_w_14363));
  bfr _b_6551(.a(_w_8453),.q(_w_8454));
  bfr _b_7608(.a(_w_9510),.q(_w_9511));
  bfr _b_5643(.a(_w_7545),.q(_w_7546));
  bfr _b_10054(.a(_w_11956),.q(_w_11957));
  bfr _b_7592(.a(_w_9494),.q(_w_9495));
  bfr _b_5644(.a(_w_7546),.q(n400_1));
  bfr _b_5326(.a(_w_7228),.q(_w_7229));
  bfr _b_5646(.a(_w_7548),.q(_w_7549));
  bfr _b_13122(.a(_w_15024),.q(_w_15025));
  bfr _b_10837(.a(_w_12739),.q(_w_12740));
  bfr _b_5647(.a(_w_7549),.q(_w_7550));
  bfr _b_5736(.a(_w_7638),.q(_w_7639));
  and_bb g1084(.a(n1073_1),.b(n1082_1),.q(_w_8202));
  bfr _b_7109(.a(_w_9011),.q(_w_9012));
  bfr _b_7817(.a(_w_9719),.q(_w_9720));
  bfr _b_5648(.a(_w_7550),.q(_w_7551));
  bfr _b_5649(.a(_w_7551),.q(_w_7552));
  bfr _b_6018(.a(_w_7920),.q(_w_7921));
  bfr _b_12041(.a(_w_13943),.q(n1580));
  bfr _b_8090(.a(_w_9992),.q(n206));
  bfr _b_9830(.a(_w_11732),.q(_w_11733));
  bfr _b_11623(.a(_w_13525),.q(_w_13526));
  bfr _b_3967(.a(_w_5869),.q(_w_5870));
  bfr _b_5653(.a(_w_7555),.q(_w_7556));
  bfr _b_5654(.a(_w_7556),.q(_w_7557));
  bfr _b_5656(.a(_w_7558),.q(_w_7559));
  bfr _b_8235(.a(_w_10137),.q(_w_10138));
  bfr _b_9752(.a(_w_11654),.q(_w_11655));
  bfr _b_5658(.a(_w_7560),.q(_w_7561));
  bfr _b_4767(.a(_w_6669),.q(_w_6670));
  bfr _b_6724(.a(_w_8626),.q(_w_8627));
  bfr _b_5660(.a(_w_7562),.q(_w_7563));
  bfr _b_10675(.a(_w_12577),.q(_w_12578));
  and_bi g845(.a(n742_1),.b(n745_1),.q(n845));
  bfr _b_5662(.a(_w_7564),.q(_w_7565));
  bfr _b_12524(.a(_w_14426),.q(_w_14427));
  bfr _b_5664(.a(_w_7566),.q(_w_7567));
  bfr _b_6048(.a(_w_7950),.q(_w_7951));
  bfr _b_3688(.a(_w_5590),.q(N256_16));
  bfr _b_5665(.a(_w_7567),.q(_w_7568));
  bfr _b_8778(.a(_w_10680),.q(_w_10681));
  bfr _b_7259(.a(_w_9161),.q(n1630));
  bfr _b_5666(.a(_w_7568),.q(_w_7569));
  bfr _b_12747(.a(_w_14649),.q(_w_14650));
  bfr _b_11696(.a(_w_13598),.q(_w_13599));
  spl2 g1500_s_0(.a(n1500),.q0(n1500_0),.q1(n1500_1));
  bfr _b_7650(.a(_w_9552),.q(_w_9553));
  bfr _b_5668(.a(_w_7570),.q(N154_11));
  bfr _b_5670(.a(_w_7572),.q(_w_7573));
  bfr _b_10020(.a(_w_11922),.q(_w_11923));
  or_bb g1356(.a(n1354_0),.b(n1355),.q(n1356));
  bfr _b_5671(.a(_w_7573),.q(_w_7574));
  bfr _b_5588(.a(_w_7490),.q(_w_7491));
  bfr _b_5673(.a(_w_7575),.q(_w_7576));
  bfr _b_5674(.a(_w_7576),.q(N222_20));
  bfr _b_5675(.a(_w_7577),.q(_w_7578));
  bfr _b_7767(.a(_w_9669),.q(_w_9670));
  bfr _b_9786(.a(_w_11688),.q(_w_11689));
  bfr _b_5677(.a(_w_7579),.q(_w_7580));
  bfr _b_5678(.a(_w_7580),.q(_w_7581));
  bfr _b_10818(.a(_w_12720),.q(N86_15));
  bfr _b_5680(.a(_w_7582),.q(_w_7583));
  bfr _b_5683(.a(_w_7585),.q(_w_7586));
  bfr _b_14343(.a(_w_16245),.q(_w_16246));
  bfr _b_7178(.a(_w_9080),.q(_w_9081));
  bfr _b_5685(.a(_w_7587),.q(_w_7588));
  bfr _b_5686(.a(_w_7588),.q(_w_7589));
  bfr _b_10571(.a(_w_12473),.q(_w_12474));
  bfr _b_5345(.a(_w_7247),.q(_w_7248));
  bfr _b_8359(.a(_w_10261),.q(_w_10262));
  bfr _b_5688(.a(_w_7590),.q(_w_7591));
  bfr _b_5689(.a(_w_7591),.q(_w_7592));
  bfr _b_13286(.a(_w_15188),.q(_w_15189));
  bfr _b_5693(.a(_w_7595),.q(_w_7596));
  bfr _b_11806(.a(_w_13708),.q(_w_13709));
  bfr _b_5695(.a(_w_7597),.q(_w_7598));
  bfr _b_5697(.a(_w_7599),.q(_w_7600));
  bfr _b_5698(.a(_w_7600),.q(_w_7601));
  bfr _b_5699(.a(_w_7601),.q(N222_16));
  bfr _b_13978(.a(_w_15880),.q(_w_15881));
  bfr _b_6432(.a(_w_8334),.q(_w_8335));
  bfr _b_5701(.a(_w_7603),.q(_w_7604));
  and_bi g414(.a(n412_0),.b(n413),.q(n414));
  bfr _b_6545(.a(_w_8447),.q(_w_8448));
  and_bb g1786(.a(N256_9),.b(N460_19),.q(_w_14349));
  bfr _b_7040(.a(_w_8942),.q(n514_1));
  bfr _b_10166(.a(_w_12068),.q(_w_12069));
  bfr _b_7648(.a(_w_9550),.q(_w_9551));
  spl2 g1401_s_0(.a(n1401),.q0(n1401_0),.q1(n1401_1));
  bfr _b_5702(.a(_w_7604),.q(N222_17));
  bfr _b_5919(.a(_w_7821),.q(_w_7822));
  bfr _b_5703(.a(_w_7605),.q(_w_7606));
  bfr _b_5706(.a(_w_7608),.q(_w_7609));
  spl2 g878_s_0(.a(n878),.q0(n878_0),.q1(n878_1));
  bfr _b_5707(.a(_w_7609),.q(_w_7610));
  bfr _b_7116(.a(_w_9018),.q(_w_9019));
  bfr _b_8257(.a(_w_10159),.q(_w_10160));
  bfr _b_5151(.a(_w_7053),.q(N103_3));
  bfr _b_5710(.a(_w_7612),.q(_w_7613));
  bfr _b_11511(.a(_w_13413),.q(_w_13414));
  bfr _b_8728(.a(_w_10630),.q(_w_10631));
  bfr _b_5711(.a(_w_7613),.q(_w_7614));
  bfr _b_9393(.a(_w_11295),.q(_w_11296));
  bfr _b_5713(.a(_w_7615),.q(_w_7616));
  bfr _b_5714(.a(_w_7616),.q(_w_7617));
  bfr _b_5717(.a(_w_7619),.q(_w_7620));
  bfr _b_5718(.a(_w_7620),.q(_w_7621));
  bfr _b_5719(.a(_w_7621),.q(_w_7622));
  bfr _b_5723(.a(_w_7625),.q(_w_7626));
  bfr _b_5724(.a(_w_7626),.q(_w_7627));
  bfr _b_5727(.a(_w_7629),.q(_w_7630));
  and_bb g1807(.a(n1780_1),.b(n1805_1),.q(_w_14540));
  bfr _b_5731(.a(_w_7633),.q(_w_7634));
  bfr _b_8348(.a(_w_10250),.q(_w_10251));
  bfr _b_5733(.a(_w_7635),.q(N222_9));
  bfr _b_5737(.a(_w_7639),.q(N222_10));
  or_bb g435(.a(n433_0),.b(n434),.q(_w_10459));
  bfr _b_5742(.a(_w_7644),.q(_w_7645));
  bfr _b_8818(.a(_w_10720),.q(_w_10721));
  bfr _b_14161(.a(_w_16063),.q(_w_16064));
  bfr _b_5747(.a(_w_7649),.q(_w_7650));
  bfr _b_12010(.a(_w_13912),.q(_w_13913));
  bfr _b_5751(.a(_w_7653),.q(_w_7654));
  and_bi g409(.a(n408_0),.b(n368_0),.q(n409));
  bfr _b_5794(.a(_w_7696),.q(_w_7697));
  bfr _b_5753(.a(_w_7655),.q(_w_7656));
  bfr _b_10125(.a(_w_12027),.q(_w_12028));
  bfr _b_5754(.a(_w_7656),.q(_w_7657));
  bfr _b_8668(.a(_w_10570),.q(n1692_1));
  bfr _b_11841(.a(_w_13743),.q(_w_13744));
  bfr _b_5756(.a(_w_7658),.q(_w_7659));
  bfr _b_12761(.a(_w_14663),.q(_w_14664));
  bfr _b_5757(.a(_w_7659),.q(_w_7660));
  bfr _b_9849(.a(_w_11751),.q(_w_11752));
  bfr _b_5758(.a(_w_7660),.q(_w_7661));
  bfr _b_9767(.a(_w_11669),.q(_w_11670));
  bfr _b_9129(.a(_w_11031),.q(_w_11032));
  and_bb g938(.a(N35_18),.b(N511_6),.q(_w_8579));
  bfr _b_5761(.a(_w_7663),.q(_w_7664));
  bfr _b_11149(.a(_w_13051),.q(_w_13052));
  bfr _b_5763(.a(_w_7665),.q(_w_7666));
  bfr _b_5765(.a(_w_7667),.q(_w_7668));
  bfr _b_5766(.a(_w_7668),.q(_w_7669));
  and_bi g288(.a(n286_0),.b(n287),.q(n288));
  bfr _b_8012(.a(_w_9914),.q(_w_9915));
  bfr _b_5767(.a(_w_7669),.q(_w_7670));
  bfr _b_4944(.a(_w_6846),.q(_w_6847));
  bfr _b_6486(.a(_w_8388),.q(n1440_1));
  bfr _b_5049(.a(_w_6951),.q(_w_6952));
  spl2 g1024_s_0(.a(n1024),.q0(n1024_0),.q1(n1024_1));
  bfr _b_5768(.a(_w_7670),.q(_w_7671));
  bfr _b_10418(.a(_w_12320),.q(_w_12321));
  bfr _b_5769(.a(_w_7671),.q(_w_7672));
  bfr _b_6431(.a(_w_8333),.q(_w_8334));
  bfr _b_13710(.a(_w_15612),.q(_w_15613));
  bfr _b_5771(.a(_w_7673),.q(_w_7674));
  bfr _b_5772(.a(_w_7674),.q(_w_7675));
  and_bi g955(.a(n869_1),.b(n872_1),.q(n955));
  bfr _b_5778(.a(_w_7680),.q(_w_7681));
  bfr _b_5779(.a(_w_7681),.q(_w_7682));
  bfr _b_5780(.a(_w_7682),.q(_w_7683));
  bfr _b_6344(.a(_w_8246),.q(_w_8247));
  bfr _b_5781(.a(_w_7683),.q(_w_7684));
  and_bb g1541(.a(N171_16),.b(N477_14),.q(n1541));
  bfr _b_3721(.a(_w_5623),.q(_w_5624));
  bfr _b_5471(.a(_w_7373),.q(_w_7374));
  bfr _b_9947(.a(_w_11849),.q(_w_11850));
  bfr _b_5784(.a(_w_7686),.q(_w_7687));
  bfr _b_12862(.a(_w_14764),.q(n1747_1));
  bfr _b_5785(.a(_w_7687),.q(_w_7688));
  bfr _b_7029(.a(_w_8931),.q(_w_8932));
  spl2 g944_s_0(.a(n944),.q0(n944_0),.q1(n944_1));
  bfr _b_10114(.a(_w_12016),.q(_w_12017));
  bfr _b_5786(.a(_w_7688),.q(_w_7689));
  bfr _b_5789(.a(_w_7691),.q(_w_7692));
  bfr _b_4048(.a(_w_5950),.q(_w_5951));
  bfr _b_3949(.a(_w_5851),.q(_w_5852));
  bfr _b_6797(.a(_w_8699),.q(_w_8700));
  bfr _b_8270(.a(_w_10172),.q(_w_10173));
  bfr _b_5790(.a(_w_7692),.q(_w_7693));
  bfr _b_6774(.a(_w_8676),.q(N222_12));
  spl2 g1282_s_0(.a(n1282),.q0(n1282_0),.q1(n1282_1));
  bfr _b_5791(.a(_w_7693),.q(_w_7694));
  bfr _b_5792(.a(_w_7694),.q(_w_7695));
  bfr _b_5796(.a(_w_7698),.q(_w_7699));
  bfr _b_5973(.a(_w_7875),.q(_w_7876));
  spl3L g308_s_0(.a(n308),.q0(n308_0),.q1(_w_14302),.q2(_w_14304));
  bfr _b_5798(.a(_w_7700),.q(_w_7701));
  bfr _b_14164(.a(_w_16066),.q(_w_16067));
  bfr _b_10954(.a(_w_12856),.q(n269));
  bfr _b_5799(.a(_w_7701),.q(_w_7702));
  bfr _b_5802(.a(_w_7704),.q(_w_7705));
  bfr _b_10784(.a(_w_12686),.q(_w_12687));
  or_bb g201(.a(n199_0),.b(n200),.q(n201));
  bfr _b_9084(.a(_w_10986),.q(_w_10987));
  bfr _b_9184(.a(_w_11086),.q(_w_11087));
  bfr _b_5804(.a(_w_7706),.q(_w_7707));
  bfr _b_5807(.a(_w_7709),.q(_w_7710));
  spl2 g1839_s_0(.a(n1839),.q0(n1839_0),.q1(_w_15040));
  bfr _b_9311(.a(_w_11213),.q(_w_11214));
  bfr _b_7820(.a(_w_9722),.q(_w_9723));
  bfr _b_5810(.a(_w_7712),.q(_w_7713));
  bfr _b_5811(.a(_w_7713),.q(_w_7714));
  bfr _b_5812(.a(_w_7714),.q(_w_7715));
  bfr _b_5813(.a(_w_7715),.q(_w_7716));
  bfr _b_11594(.a(_w_13496),.q(_w_13497));
  bfr _b_5815(.a(_w_7717),.q(_w_7718));
  bfr _b_5817(.a(_w_7719),.q(N222_6));
  bfr _b_14055(.a(_w_15957),.q(_w_15958));
  bfr _b_5821(.a(_w_7723),.q(_w_7724));
  bfr _b_5058(.a(_w_6960),.q(_w_6961));
  bfr _b_5822(.a(_w_7724),.q(_w_7725));
  bfr _b_5823(.a(_w_7725),.q(_w_7726));
  bfr _b_14157(.a(_w_16059),.q(_w_16060));
  bfr _b_5824(.a(_w_7726),.q(_w_7727));
  bfr _b_9661(.a(_w_11563),.q(_w_11564));
  bfr _b_5826(.a(_w_7728),.q(_w_7729));
  bfr _b_9398(.a(_w_11300),.q(_w_11301));
  bfr _b_5827(.a(_w_7729),.q(_w_7730));
  bfr _b_5828(.a(_w_7730),.q(_w_7731));
  bfr _b_14021(.a(_w_15923),.q(_w_15924));
  bfr _b_5830(.a(_w_7732),.q(_w_7733));
  bfr _b_8184(.a(_w_10086),.q(_w_10087));
  bfr _b_5834(.a(_w_7736),.q(_w_7737));
  bfr _b_5942(.a(_w_7844),.q(_w_7845));
  bfr _b_5835(.a(_w_7737),.q(_w_7738));
  bfr _b_8278(.a(_w_10180),.q(n1729));
  bfr _b_11609(.a(_w_13511),.q(n1367));
  bfr _b_4097(.a(_w_5999),.q(_w_6000));
  bfr _b_5838(.a(_w_7740),.q(_w_7741));
  bfr _b_3860(.a(_w_5762),.q(_w_5763));
  bfr _b_5840(.a(_w_7742),.q(_w_7743));
  bfr _b_5843(.a(_w_7745),.q(_w_7746));
  bfr _b_5845(.a(_w_7747),.q(_w_7748));
  bfr _b_10911(.a(_w_12813),.q(_w_12814));
  bfr _b_5847(.a(_w_7749),.q(_w_7750));
  bfr _b_12671(.a(_w_14573),.q(_w_14574));
  bfr _b_5848(.a(_w_7750),.q(_w_7751));
  bfr _b_5850(.a(_w_7752),.q(_w_7753));
  bfr _b_5851(.a(_w_7753),.q(_w_7754));
  bfr _b_14068(.a(_w_15970),.q(_w_15971));
  bfr _b_4196(.a(_w_6098),.q(_w_6099));
  bfr _b_3767(.a(_w_5669),.q(_w_5670));
  bfr _b_5855(.a(_w_7757),.q(_w_7758));
  bfr _b_7994(.a(_w_9896),.q(_w_9897));
  bfr _b_8464(.a(_w_10366),.q(_w_10367));
  bfr _b_5857(.a(_w_7759),.q(N222_7));
  bfr _b_4711(.a(_w_6613),.q(_w_6614));
  bfr _b_9206(.a(_w_11108),.q(n565));
  bfr _b_12034(.a(_w_13936),.q(_w_13937));
  bfr _b_5859(.a(_w_7761),.q(_w_7762));
  and_bi g410(.a(n368_1),.b(n408_1),.q(_w_15109));
  bfr _b_10126(.a(_w_12028),.q(_w_12029));
  bfr _b_5861(.a(_w_7763),.q(_w_7764));
  bfr _b_5865(.a(_w_7767),.q(_w_7768));
  bfr _b_6157(.a(_w_8059),.q(_w_8060));
  bfr _b_5866(.a(_w_7768),.q(_w_7769));
  bfr _b_3573(.a(_w_5475),.q(_w_5476));
  bfr _b_5867(.a(_w_7769),.q(_w_7770));
  bfr _b_14352(.a(_w_16254),.q(_w_16255));
  bfr _b_5871(.a(_w_7773),.q(_w_7774));
  bfr _b_6011(.a(_w_7913),.q(_w_7914));
  bfr _b_14050(.a(_w_15952),.q(_w_15953));
  and_bb g912(.a(n827_1),.b(n910_1),.q(_w_8779));
  bfr _b_5876(.a(_w_7778),.q(_w_7779));
  bfr _b_7202(.a(_w_9104),.q(_w_9105));
  bfr _b_5881(.a(_w_7783),.q(_w_7784));
  bfr _b_5884(.a(_w_7786),.q(_w_7787));
  bfr _b_5886(.a(_w_7788),.q(_w_7789));
  bfr _b_9686(.a(_w_11588),.q(_w_11589));
  bfr _b_5888(.a(_w_7790),.q(_w_7791));
  bfr _b_5889(.a(_w_7791),.q(_w_7792));
  bfr _b_5890(.a(_w_7792),.q(_w_7793));
  bfr _b_5892(.a(_w_7794),.q(_w_7795));
  bfr _b_5893(.a(_w_7795),.q(_w_7796));
  bfr _b_12074(.a(_w_13976),.q(n1633));
  bfr _b_6756(.a(_w_8658),.q(_w_8659));
  or_bb g1242(.a(n1168_0),.b(n1241_0),.q(n1242));
  bfr _b_5895(.a(_w_7797),.q(_w_7798));
  bfr _b_10898(.a(_w_12800),.q(_w_12801));
  bfr _b_5896(.a(_w_7798),.q(_w_7799));
  bfr _b_6509(.a(_w_8411),.q(_w_8412));
  bfr _b_3869(.a(_w_5771),.q(_w_5772));
  bfr _b_9737(.a(_w_11639),.q(_w_11640));
  bfr _b_7729(.a(_w_9631),.q(_w_9632));
  bfr _b_6953(.a(_w_8855),.q(_w_8856));
  bfr _b_9070(.a(_w_10972),.q(_w_10973));
  bfr _b_5900(.a(_w_7802),.q(_w_7803));
  bfr _b_13015(.a(_w_14917),.q(_w_14918));
  bfr _b_5901(.a(_w_7803),.q(_w_7804));
  bfr _b_5902(.a(_w_7804),.q(_w_7805));
  bfr _b_9607(.a(_w_11509),.q(_w_11510));
  bfr _b_10789(.a(_w_12691),.q(_w_12692));
  bfr _b_9743(.a(_w_11645),.q(_w_11646));
  bfr _b_10670(.a(_w_12572),.q(_w_12573));
  and_bi g1560(.a(n1558_0),.b(n1559),.q(n1560));
  bfr _b_5903(.a(_w_7805),.q(_w_7806));
  bfr _b_5307(.a(_w_7209),.q(_w_7210));
  bfr _b_5904(.a(_w_7806),.q(_w_7807));
  bfr _b_14173(.a(_w_16075),.q(_w_16076));
  bfr _b_13338(.a(_w_15240),.q(_w_15241));
  bfr _b_9181(.a(_w_11083),.q(_w_11084));
  bfr _b_12229(.a(_w_14131),.q(_w_14132));
  bfr _b_11226(.a(_w_13128),.q(_w_13129));
  bfr _b_5905(.a(_w_7807),.q(_w_7808));
  bfr _b_5906(.a(_w_7808),.q(N222_0));
  bfr _b_5964(.a(_w_7866),.q(_w_7867));
  bfr _b_3666(.a(_w_5568),.q(n998_1));
  or_bb g1844(.a(n1842_0),.b(n1843),.q(n1844));
  spl2 g1302_s_0(.a(n1302),.q0(n1302_0),.q1(n1302_1));
  bfr _b_5907(.a(_w_7809),.q(_w_7810));
  bfr _b_5912(.a(_w_7814),.q(_w_7815));
  spl2 g673_s_0(.a(n673),.q0(n673_0),.q1(n673_1));
  bfr _b_5915(.a(_w_7817),.q(_w_7818));
  bfr _b_5916(.a(_w_7818),.q(_w_7819));
  bfr _b_5917(.a(_w_7819),.q(_w_7820));
  bfr _b_5925(.a(_w_7827),.q(_w_7828));
  or_bb g208(.a(n187_0),.b(n207_0),.q(n208));
  bfr _b_5931(.a(_w_7833),.q(_w_7834));
  bfr _b_11401(.a(_w_13303),.q(_w_13304));
  bfr _b_5936(.a(_w_7838),.q(_w_7839));
  bfr _b_7714(.a(_w_9616),.q(_w_9617));
  bfr _b_11741(.a(_w_13643),.q(_w_13644));
  bfr _b_11639(.a(_w_13541),.q(n146_1));
  bfr _b_8162(.a(_w_10064),.q(_w_10065));
  bfr _b_5937(.a(_w_7839),.q(_w_7840));
  bfr _b_12260(.a(_w_14162),.q(_w_14163));
  bfr _b_6568(.a(_w_8470),.q(N205_2));
  bfr _b_9744(.a(_w_11646),.q(_w_11647));
  bfr _b_14017(.a(_w_15919),.q(_w_15920));
  bfr _b_5940(.a(_w_7842),.q(_w_7843));
  bfr _b_5408(.a(_w_7310),.q(_w_7311));
  bfr _b_5943(.a(_w_7845),.q(_w_7846));
  bfr _b_5944(.a(_w_7846),.q(_w_7847));
  spl2 g62_s_0(.a(n62),.q0(n62_0),.q1(n62_1));
  bfr _b_8737(.a(_w_10639),.q(_w_10640));
  bfr _b_5955(.a(_w_7857),.q(_w_7858));
  bfr _b_5957(.a(_w_7859),.q(_w_7860));
  bfr _b_4989(.a(_w_6891),.q(_w_6892));
  bfr _b_5958(.a(_w_7860),.q(_w_7861));
  bfr _b_5960(.a(_w_7862),.q(_w_7863));
  bfr _b_14084(.a(_w_15986),.q(_w_15987));
  bfr _b_5961(.a(_w_7863),.q(_w_7864));
  bfr _b_5963(.a(_w_7865),.q(_w_7866));
  bfr _b_4895(.a(_w_6797),.q(_w_6798));
  and_bi g1030(.a(n1028_0),.b(n1029),.q(n1030));
  bfr _b_5965(.a(_w_7867),.q(_w_7868));
  or_bb g1811(.a(n1809_0),.b(n1810),.q(n1811));
  bfr _b_5967(.a(_w_7869),.q(_w_7870));
  bfr _b_5968(.a(_w_7870),.q(_w_7871));
  bfr _b_8597(.a(_w_10499),.q(_w_10500));
  bfr _b_11001(.a(_w_12903),.q(_w_12904));
  bfr _b_3819(.a(_w_5721),.q(_w_5722));
  bfr _b_9878(.a(_w_11780),.q(_w_11781));
  bfr _b_5969(.a(_w_7871),.q(_w_7872));
  bfr _b_9695(.a(_w_11597),.q(n638));
  bfr _b_12893(.a(_w_14795),.q(_w_14796));
  bfr _b_5970(.a(_w_7872),.q(_w_7873));
  bfr _b_8917(.a(_w_10819),.q(n812));
  spl4L N35_s_3(.a(N35_2),.q0(N35_12),.q1(_w_12446),.q2(_w_12454),.q3(_w_12466));
  bfr _b_5975(.a(_w_7877),.q(_w_7878));
  or_bb g150(.a(n108_1),.b(n149_0),.q(n150));
  bfr _b_5976(.a(_w_7878),.q(_w_7879));
  bfr _b_11643(.a(_w_13545),.q(_w_13546));
  bfr _b_9079(.a(_w_10981),.q(n873));
  bfr _b_5437(.a(_w_7339),.q(_w_7340));
  bfr _b_5977(.a(_w_7879),.q(_w_7880));
  bfr _b_5978(.a(_w_7880),.q(n1485_1));
  spl4L N290_s_4(.a(N290_3),.q0(N290_16),.q1(N290_17),.q2(N290_18),.q3(_w_7889));
  bfr _b_4760(.a(_w_6662),.q(_w_6663));
  bfr _b_5980(.a(_w_7882),.q(_w_7883));
  or_bb g477(.a(n475_0),.b(n476),.q(n477));
  bfr _b_8153(.a(_w_10055),.q(_w_10056));
  bfr _b_5982(.a(_w_7884),.q(n502_1));
  bfr _b_4532(.a(_w_6434),.q(_w_6435));
  bfr _b_9292(.a(_w_11194),.q(_w_11195));
  bfr _b_5986(.a(_w_7888),.q(n456_2));
  bfr _b_14072(.a(_w_15974),.q(_w_15975));
  spl2 g1268_s_0(.a(n1268),.q0(n1268_0),.q1(n1268_1));
  bfr _b_5987(.a(_w_7889),.q(_w_7890));
  and_bi g1495(.a(n1464_1),.b(n1493_1),.q(_w_12032));
  bfr _b_5988(.a(_w_7890),.q(_w_7891));
  bfr _b_5989(.a(_w_7891),.q(N290_19));
  bfr _b_5991(.a(_w_7893),.q(n378_1));
  bfr _b_5993(.a(_w_7895),.q(n378_2));
  bfr _b_7541(.a(_w_9443),.q(_w_9444));
  bfr _b_5994(.a(_w_7896),.q(_w_7897));
  bfr _b_13079(.a(_w_14981),.q(_w_14982));
  bfr _b_5995(.a(_w_7897),.q(_w_7898));
  bfr _b_3537(.a(_w_5439),.q(_w_5440));
  bfr _b_5996(.a(_w_7898),.q(_w_7899));
  bfr _b_7905(.a(_w_9807),.q(_w_9808));
  and_bb g1005(.a(n1003_1),.b(n949_1),.q(_w_8361));
  bfr _b_5997(.a(_w_7899),.q(_w_7900));
  spl4L N120_s_2(.a(N120_1),.q0(N120_8),.q1(N120_9),.q2(N120_10),.q3(_w_6244));
  spl2 g114_s_0(.a(n114),.q0(n114_0),.q1(n114_1));
  bfr _b_5998(.a(_w_7900),.q(_w_7901));
  bfr _b_11852(.a(_w_13754),.q(_w_13755));
  bfr _b_11099(.a(_w_13001),.q(n1201));
  bfr _b_6001(.a(_w_7903),.q(N188_13));
  bfr _b_4724(.a(_w_6626),.q(_w_6627));
  bfr _b_6002(.a(_w_7904),.q(_w_7905));
  bfr _b_7339(.a(_w_9241),.q(_w_9242));
  bfr _b_6003(.a(_w_7905),.q(_w_7906));
  bfr _b_6006(.a(_w_7908),.q(_w_7909));
  bfr _b_6532(.a(_w_8434),.q(_w_8435));
  bfr _b_6007(.a(_w_7909),.q(_w_7910));
  and_bi g1555(.a(n1554_0),.b(n1549_0),.q(n1555));
  bfr _b_6008(.a(_w_7910),.q(_w_7911));
  and_bb g325(.a(n303_1),.b(n323_1),.q(_w_11026));
  bfr _b_6009(.a(_w_7911),.q(_w_7912));
  bfr _b_12777(.a(_w_14679),.q(_w_14680));
  bfr _b_6013(.a(_w_7915),.q(N188_14));
  bfr _b_9412(.a(_w_11314),.q(_w_11315));
  bfr _b_6017(.a(_w_7919),.q(_w_7920));
  bfr _b_6020(.a(_w_7922),.q(_w_7923));
  bfr _b_8080(.a(_w_9982),.q(_w_9983));
  bfr _b_12265(.a(_w_14167),.q(_w_14168));
  bfr _b_12073(.a(_w_13975),.q(n544));
  bfr _b_6027(.a(_w_7929),.q(_w_7930));
  spl2 g1677_s_0(.a(n1677),.q0(n1677_0),.q1(n1677_1));
  bfr _b_8931(.a(_w_10833),.q(_w_10834));
  or_bb g38(.a(n36_0),.b(n37),.q(_w_10882));
  bfr _b_6030(.a(_w_7932),.q(_w_7933));
  bfr _b_12739(.a(_w_14641),.q(_w_14642));
  bfr _b_6031(.a(_w_7933),.q(_w_7934));
  bfr _b_6036(.a(_w_7938),.q(_w_7939));
  bfr _b_7532(.a(_w_9434),.q(_w_9435));
  bfr _b_6037(.a(_w_7939),.q(_w_7940));
  bfr _b_7782(.a(_w_9684),.q(n1862));
  bfr _b_6038(.a(_w_7940),.q(_w_7941));
  bfr _b_6039(.a(_w_7941),.q(_w_7942));
  bfr _b_6040(.a(_w_7942),.q(_w_7943));
  bfr _b_9018(.a(_w_10920),.q(_w_10921));
  bfr _b_6042(.a(_w_7944),.q(_w_7945));
  bfr _b_6043(.a(_w_7945),.q(_w_7946));
  and_bi g1586(.a(n1539_1),.b(n1584_1),.q(_w_13950));
  bfr _b_6044(.a(_w_7946),.q(_w_7947));
  bfr _b_6515(.a(_w_8417),.q(_w_8418));
  bfr _b_6045(.a(_w_7947),.q(_w_7948));
  and_bb g1243(.a(n1168_1),.b(n1241_1),.q(_w_8925));
  bfr _b_6703(.a(_w_8605),.q(_w_8606));
  bfr _b_13295(.a(_w_15197),.q(_w_15198));
  bfr _b_6047(.a(_w_7949),.q(_w_7950));
  bfr _b_14381(.a(_w_16283),.q(_w_16284));
  bfr _b_3774(.a(_w_5676),.q(_w_5677));
  bfr _b_6053(.a(_w_7955),.q(N188_7));
  bfr _b_6055(.a(_w_7957),.q(_w_7958));
  bfr _b_6056(.a(_w_7958),.q(_w_7959));
  bfr _b_7524(.a(_w_9426),.q(_w_9427));
  bfr _b_6058(.a(_w_7960),.q(_w_7961));
  bfr _b_6059(.a(_w_7961),.q(n246_1));
  bfr _b_6061(.a(_w_7963),.q(n246_2));
  bfr _b_8239(.a(_w_10141),.q(_w_10142));
  bfr _b_13741(.a(_w_15643),.q(_w_15644));
  spl2 g1058_s_0(.a(n1058),.q0(n1058_0),.q1(n1058_1));
  bfr _b_6064(.a(_w_7966),.q(_w_7967));
  bfr _b_6065(.a(_w_7967),.q(_w_7968));
  bfr _b_6067(.a(_w_7969),.q(_w_7970));
  bfr _b_8458(.a(_w_10360),.q(_w_10361));
  bfr _b_6069(.a(_w_7971),.q(N205_13));
  bfr _b_11412(.a(_w_13314),.q(_w_13315));
  bfr _b_6070(.a(_w_7972),.q(_w_7973));
  bfr _b_6073(.a(_w_7975),.q(_w_7976));
  bfr _b_12701(.a(_w_14603),.q(_w_14604));
  bfr _b_9747(.a(_w_11649),.q(_w_11650));
  and_bb g247(.a(N137_5),.b(N273_12),.q(n247));
  bfr _b_6074(.a(_w_7976),.q(_w_7977));
  bfr _b_6075(.a(_w_7977),.q(_w_7978));
  bfr _b_8964(.a(_w_10866),.q(_w_10867));
  bfr _b_8660(.a(_w_10562),.q(_w_10563));
  bfr _b_4484(.a(_w_6386),.q(_w_6387));
  bfr _b_6078(.a(_w_7980),.q(_w_7981));
  and_bb g40(.a(N1_6),.b(N307_4),.q(_w_13571));
  bfr _b_6080(.a(_w_7982),.q(_w_7983));
  and_bi g709(.a(n708_0),.b(n612_0),.q(n709));
  bfr _b_6081(.a(_w_7983),.q(N205_14));
  bfr _b_6082(.a(_w_7984),.q(_w_7985));
  bfr _b_6083(.a(_w_7985),.q(_w_7986));
  and_bi g237(.a(n214_1),.b(n217_1),.q(n237));
  bfr _b_6085(.a(_w_7987),.q(_w_7988));
  bfr _b_7964(.a(_w_9866),.q(_w_9867));
  bfr _b_6086(.a(_w_7988),.q(_w_7989));
  bfr _b_11360(.a(_w_13262),.q(_w_13263));
  bfr _b_6088(.a(_w_7990),.q(_w_7991));
  bfr _b_5585(.a(_w_7487),.q(_w_7488));
  bfr _b_6090(.a(_w_7992),.q(_w_7993));
  bfr _b_7811(.a(_w_9713),.q(_w_9714));
  bfr _b_13030(.a(_w_14932),.q(_w_14933));
  bfr _b_6092(.a(_w_7994),.q(_w_7995));
  bfr _b_10656(.a(_w_12558),.q(_w_12559));
  bfr _b_6093(.a(_w_7995),.q(N205_15));
  bfr _b_6097(.a(_w_7999),.q(_w_8000));
  bfr _b_6098(.a(_w_8000),.q(_w_8001));
  bfr _b_12061(.a(_w_13963),.q(_w_13964));
  spl2 g1490_s_0(.a(n1490),.q0(n1490_0),.q1(n1490_1));
  bfr _b_6100(.a(_w_8002),.q(_w_8003));
  bfr _b_7318(.a(_w_9220),.q(n692));
  bfr _b_5593(.a(_w_7495),.q(_w_7496));
  bfr _b_6101(.a(_w_8003),.q(_w_8004));
  bfr _b_6102(.a(_w_8004),.q(_w_8005));
  bfr _b_6107(.a(_w_8009),.q(_w_8010));
  bfr _b_6108(.a(_w_8010),.q(_w_8011));
  bfr _b_10810(.a(_w_12712),.q(_w_12713));
  bfr _b_7430(.a(_w_9332),.q(_w_9333));
  and_bb g491(.a(n445_1),.b(n489_1),.q(_w_12364));
  bfr _b_6110(.a(_w_8012),.q(_w_8013));
  bfr _b_6569(.a(_w_8471),.q(_w_8472));
  bfr _b_6114(.a(_w_8016),.q(_w_8017));
  bfr _b_6115(.a(_w_8017),.q(_w_8018));
  bfr _b_13449(.a(_w_15351),.q(_w_15352));
  bfr _b_6120(.a(_w_8022),.q(_w_8023));
  bfr _b_7480(.a(_w_9382),.q(_w_9383));
  bfr _b_9262(.a(_w_11164),.q(_w_11165));
  bfr _b_7058(.a(_w_8960),.q(n1117));
  bfr _b_6122(.a(_w_8024),.q(_w_8025));
  bfr _b_12459(.a(_w_14361),.q(_w_14362));
  bfr _b_7281(.a(_w_9183),.q(_w_9184));
  bfr _b_6123(.a(_w_8025),.q(_w_8026));
  bfr _b_5519(.a(_w_7421),.q(_w_7422));
  bfr _b_6124(.a(_w_8026),.q(_w_8027));
  bfr _b_8970(.a(_w_10872),.q(_w_10873));
  bfr _b_6125(.a(_w_8027),.q(n1357_1));
  bfr _b_8186(.a(_w_10088),.q(_w_10089));
  or_bb g663(.a(n661_0),.b(n662),.q(n663));
  bfr _b_7520(.a(_w_9422),.q(_w_9423));
  bfr _b_6126(.a(_w_8028),.q(_w_8029));
  bfr _b_6128(.a(_w_8030),.q(_w_8031));
  spl2 g1409_s_0(.a(n1409),.q0(n1409_0),.q1(n1409_1));
  bfr _b_5380(.a(_w_7282),.q(_w_7283));
  bfr _b_6130(.a(_w_8032),.q(_w_8033));
  bfr _b_7125(.a(_w_9027),.q(_w_9028));
  bfr _b_13115(.a(_w_15017),.q(_w_15018));
  bfr _b_9050(.a(_w_10952),.q(_w_10953));
  bfr _b_6132(.a(_w_8034),.q(_w_8035));
  bfr _b_10300(.a(_w_12202),.q(_w_12203));
  spl2 g1360_s_0(.a(n1360),.q0(n1360_0),.q1(n1360_1));
  bfr _b_6133(.a(_w_8035),.q(n196_1));
  bfr _b_7967(.a(_w_9869),.q(_w_9870));
  bfr _b_6135(.a(_w_8037),.q(_w_8038));
  bfr _b_12449(.a(_w_14351),.q(_w_14352));
  bfr _b_6137(.a(_w_8039),.q(_w_8040));
  bfr _b_6139(.a(_w_8041),.q(_w_8042));
  bfr _b_6141(.a(_w_8043),.q(_w_8044));
  bfr _b_6143(.a(_w_8045),.q(_w_8046));
  bfr _b_12523(.a(_w_14425),.q(_w_14426));
  bfr _b_4938(.a(_w_6840),.q(_w_6841));
  bfr _b_5621(.a(_w_7523),.q(_w_7524));
  bfr _b_9312(.a(_w_11214),.q(_w_11215));
  bfr _b_6144(.a(_w_8046),.q(_w_8047));
  and_bi g702(.a(n700_0),.b(n701),.q(n702));
  bfr _b_6147(.a(_w_8049),.q(_w_8050));
  bfr _b_8647(.a(_w_10549),.q(_w_10550));
  bfr _b_6148(.a(_w_8050),.q(_w_8051));
  bfr _b_7593(.a(_w_9495),.q(_w_9496));
  bfr _b_11944(.a(_w_13846),.q(_w_13847));
  bfr _b_6150(.a(_w_8052),.q(_w_8053));
  bfr _b_6151(.a(_w_8053),.q(_w_8054));
  bfr _b_6019(.a(_w_7921),.q(_w_7922));
  bfr _b_6152(.a(_w_8054),.q(_w_8055));
  bfr _b_12474(.a(_w_14376),.q(_w_14377));
  bfr _b_4733(.a(_w_6635),.q(_w_6636));
  bfr _b_8959(.a(_w_10861),.q(_w_10862));
  bfr _b_10039(.a(_w_11941),.q(_w_11942));
  bfr _b_6153(.a(_w_8055),.q(_w_8056));
  bfr _b_6158(.a(_w_8060),.q(_w_8061));
  bfr _b_6531(.a(_w_8433),.q(_w_8434));
  bfr _b_6159(.a(_w_8061),.q(_w_8062));
  bfr _b_6160(.a(_w_8062),.q(_w_8063));
  bfr _b_6161(.a(_w_8063),.q(_w_8064));
  bfr _b_6162(.a(_w_8064),.q(_w_8065));
  bfr _b_9545(.a(_w_11447),.q(_w_11448));
  or_bb g135(.a(n133_0),.b(n134),.q(_w_13206));
  bfr _b_9584(.a(_w_11486),.q(_w_11487));
  bfr _b_6163(.a(_w_8065),.q(_w_8066));
  bfr _b_6165(.a(_w_8067),.q(_w_8068));
  bfr _b_5379(.a(_w_7281),.q(_w_7282));
  bfr _b_6169(.a(_w_8071),.q(_w_8072));
  bfr _b_12153(.a(_w_14055),.q(_w_14056));
  bfr _b_6170(.a(_w_8072),.q(_w_8073));
  bfr _b_7588(.a(_w_9490),.q(_w_9491));
  bfr _b_6171(.a(_w_8073),.q(_w_8074));
  bfr _b_9263(.a(_w_11165),.q(_w_11166));
  bfr _b_6172(.a(_w_8074),.q(_w_8075));
  bfr _b_6917(.a(_w_8819),.q(_w_8820));
  bfr _b_6725(.a(_w_8627),.q(_w_8628));
  bfr _b_4954(.a(_w_6856),.q(_w_6857));
  or_bb g910(.a(n908_0),.b(n909),.q(n910));
  bfr _b_6176(.a(_w_8078),.q(_w_8079));
  bfr _b_6180(.a(_w_8082),.q(_w_8083));
  bfr _b_6182(.a(_w_8084),.q(N256_12));
  bfr _b_12958(.a(_w_14860),.q(_w_14861));
  bfr _b_6183(.a(_w_8085),.q(_w_8086));
  bfr _b_13540(.a(_w_15442),.q(_w_15443));
  bfr _b_6186(.a(_w_8088),.q(_w_8089));
  bfr _b_8421(.a(_w_10323),.q(_w_10324));
  bfr _b_9150(.a(_w_11052),.q(_w_11053));
  bfr _b_6187(.a(_w_8089),.q(_w_8090));
  bfr _b_7670(.a(_w_9572),.q(_w_9573));
  spl4L N154_s_1(.a(N154_0),.q0(N154_4),.q1(N154_5),.q2(_w_6462),.q3(_w_6464));
  and_bi g555(.a(n554_0),.b(n538_0),.q(n555));
  and_bi g550(.a(n540_1),.b(n548_1),.q(_w_12731));
  bfr _b_6189(.a(_w_8091),.q(_w_8092));
  bfr _b_13660(.a(_w_15562),.q(_w_15563));
  bfr _b_6190(.a(_w_8092),.q(_w_8093));
  bfr _b_7930(.a(_w_9832),.q(_w_9833));
  bfr _b_13143(.a(_w_15045),.q(_w_15046));
  bfr _b_8832(.a(_w_10734),.q(_w_10735));
  bfr _b_6191(.a(_w_8093),.q(_w_8094));
  bfr _b_6193(.a(_w_8095),.q(_w_8096));
  bfr _b_3892(.a(_w_5794),.q(_w_5795));
  bfr _b_9697(.a(_w_11599),.q(n148));
  bfr _b_6194(.a(_w_8096),.q(_w_8097));
  bfr _b_6197(.a(_w_8099),.q(_w_8100));
  bfr _b_6199(.a(_w_8101),.q(N256_14));
  bfr _b_10872(.a(_w_12774),.q(_w_12775));
  and_bi g708(.a(n706_0),.b(n707),.q(n708));
  and_bi g1873(.a(n1872_0),.b(n1851_0),.q(n1873));
  bfr _b_6201(.a(_w_8103),.q(_w_8104));
  spl2 g1664_s_0(.a(n1664),.q0(n1664_0),.q1(n1664_1));
  bfr _b_6202(.a(_w_8104),.q(_w_8105));
  bfr _b_9685(.a(_w_11587),.q(_w_11588));
  bfr _b_6203(.a(_w_8105),.q(_w_8106));
  bfr _b_12952(.a(_w_14854),.q(_w_14855));
  bfr _b_7152(.a(_w_9054),.q(_w_9055));
  bfr _b_11260(.a(_w_13162),.q(_w_13163));
  and_bi g661(.a(n660_0),.b(n628_0),.q(n661));
  bfr _b_6204(.a(_w_8106),.q(_w_8107));
  bfr _b_6207(.a(_w_8109),.q(_w_8110));
  bfr _b_13898(.a(_w_15800),.q(_w_15801));
  spl2 g1767_s_0(.a(n1767),.q0(n1767_0),.q1(n1767_1));
  bfr _b_9535(.a(_w_11437),.q(_w_11438));
  bfr _b_5722(.a(_w_7624),.q(_w_7625));
  spl2 g388_s_0(.a(n388),.q0(n388_0),.q1(_w_13087));
  bfr _b_6214(.a(_w_8116),.q(_w_8117));
  bfr _b_5248(.a(_w_7150),.q(_w_7151));
  bfr _b_6215(.a(_w_8117),.q(_w_8118));
  bfr _b_3833(.a(_w_5735),.q(_w_5736));
  spl2 g1263_s_0(.a(n1263),.q0(n1263_0),.q1(n1263_1));
  bfr _b_6216(.a(_w_8118),.q(N256_15));
  bfr _b_6748(.a(_w_8650),.q(_w_8651));
  bfr _b_7740(.a(_w_9642),.q(_w_9643));
  bfr _b_6219(.a(_w_8121),.q(_w_8122));
  bfr _b_6222(.a(_w_8124),.q(_w_8125));
  bfr _b_11879(.a(_w_13781),.q(_w_13782));
  bfr _b_6223(.a(_w_8125),.q(_w_8126));
  bfr _b_12075(.a(_w_13977),.q(n1642));
  and_bi g1191(.a(n1190_0),.b(n1185_0),.q(n1191));
  or_bb g973(.a(n971_0),.b(n972),.q(n973));
  bfr _b_9782(.a(_w_11684),.q(_w_11685));
  bfr _b_6224(.a(_w_8126),.q(n478_1));
  bfr _b_13713(.a(_w_15615),.q(_w_15616));
  bfr _b_4403(.a(_w_6305),.q(_w_6306));
  and_bb g245(.a(N137_4),.b(N290_12),.q(n245));
  bfr _b_6226(.a(_w_8128),.q(_w_8129));
  bfr _b_6227(.a(_w_8129),.q(_w_8130));
  bfr _b_9989(.a(_w_11891),.q(_w_11892));
  bfr _b_6228(.a(_w_8130),.q(n330_1));
  bfr _b_13154(.a(_w_15056),.q(n1428_1));
  bfr _b_6229(.a(_w_8131),.q(_w_8132));
  bfr _b_3733(.a(_w_5635),.q(_w_5636));
  bfr _b_5433(.a(_w_7335),.q(_w_7336));
  bfr _b_6230(.a(_w_8132),.q(_w_8133));
  bfr _b_6231(.a(_w_8133),.q(_w_8134));
  bfr _b_13922(.a(_w_15824),.q(_w_15825));
  bfr _b_8884(.a(_w_10786),.q(_w_10787));
  bfr _b_6232(.a(_w_8134),.q(n348_1));
  bfr _b_14223(.a(_w_16125),.q(_w_16126));
  bfr _b_6602(.a(_w_8504),.q(_w_8505));
  spl2 g184_s_0(.a(n184),.q0(n184_0),.q1(n184_1));
  and_bi g1366(.a(n1345_1),.b(n1348_1),.q(n1366));
  bfr _b_6234(.a(_w_8136),.q(_w_8137));
  bfr _b_6239(.a(_w_8141),.q(_w_8142));
  bfr _b_7483(.a(_w_9385),.q(_w_9386));
  bfr _b_6240(.a(_w_8142),.q(n986_1));
  bfr _b_7095(.a(_w_8997),.q(_w_8998));
  bfr _b_8515(.a(_w_10417),.q(_w_10418));
  and_bb g1068(.a(N188_10),.b(N375_15),.q(_w_8182));
  bfr _b_6243(.a(_w_8145),.q(_w_8146));
  bfr _b_6244(.a(_w_8146),.q(n130_1));
  bfr _b_12202(.a(_w_14104),.q(_w_14105));
  bfr _b_6248(.a(_w_8150),.q(N392_19));
  bfr _b_10932(.a(_w_12834),.q(_w_12835));
  bfr _b_6119(.a(_w_8021),.q(N205_6));
  bfr _b_6249(.a(_w_8151),.q(n248));
  bfr _b_6250(.a(_w_8152),.q(n1132));
  bfr _b_14315(.a(_w_16217),.q(_w_16218));
  and_bi g1436(.a(n1434_0),.b(n1435),.q(n1436));
  bfr _b_6252(.a(_w_8154),.q(n607));
  bfr _b_6254(.a(_w_8156),.q(_w_8157));
  bfr _b_4095(.a(_w_5997),.q(_w_5998));
  bfr _b_7836(.a(_w_9738),.q(n1531));
  bfr _b_6255(.a(_w_8157),.q(_w_8158));
  bfr _b_6257(.a(_w_8159),.q(_w_8160));
  bfr _b_6258(.a(_w_8160),.q(_w_8161));
  bfr _b_7341(.a(_w_9243),.q(n683));
  bfr _b_6261(.a(_w_8163),.q(_w_8164));
  bfr _b_6262(.a(_w_8164),.q(_w_8165));
  bfr _b_11348(.a(_w_13250),.q(_w_13251));
  bfr _b_6792(.a(_w_8694),.q(_w_8695));
  or_bb g1155(.a(n1049_0),.b(n1154_0),.q(n1155));
  bfr _b_6263(.a(_w_8165),.q(_w_8166));
  bfr _b_6265(.a(_w_8167),.q(_w_8168));
  bfr _b_8068(.a(_w_9970),.q(_w_9971));
  bfr _b_6267(.a(_w_8169),.q(_w_8170));
  bfr _b_6270(.a(_w_8172),.q(_w_8173));
  bfr _b_8181(.a(_w_10083),.q(_w_10084));
  spl2 g866_s_0(.a(n866),.q0(n866_0),.q1(n866_1));
  bfr _b_6271(.a(_w_8173),.q(_w_8174));
  bfr _b_6272(.a(_w_8174),.q(_w_8175));
  bfr _b_6273(.a(_w_8175),.q(_w_8176));
  bfr _b_6274(.a(_w_8176),.q(_w_8177));
  bfr _b_14065(.a(_w_15967),.q(_w_15968));
  bfr _b_6275(.a(_w_8177),.q(_w_8178));
  bfr _b_6277(.a(_w_8179),.q(n1114));
  spl4L N256_s_1(.a(N256_0),.q0(N256_4),.q1(_w_5591),.q2(_w_5627),.q3(_w_5663));
  bfr _b_6278(.a(_w_8180),.q(n1108));
  bfr _b_6282(.a(_w_8184),.q(_w_8185));
  bfr _b_3905(.a(_w_5807),.q(_w_5808));
  bfr _b_6283(.a(_w_8185),.q(_w_8186));
  bfr _b_10600(.a(_w_12502),.q(_w_12503));
  spl2 g887_s_0(.a(n887),.q0(n887_0),.q1(_w_11063));
  bfr _b_6284(.a(_w_8186),.q(_w_8187));
  bfr _b_6285(.a(_w_8187),.q(_w_8188));
  bfr _b_6289(.a(_w_8191),.q(_w_8192));
  bfr _b_5187(.a(_w_7089),.q(_w_7090));
  bfr _b_6290(.a(_w_8192),.q(_w_8193));
  bfr _b_6297(.a(_w_8199),.q(n1111));
  bfr _b_11036(.a(_w_12938),.q(_w_12939));
  bfr _b_6298(.a(_w_8200),.q(n1093));
  bfr _b_6299(.a(_w_8201),.q(n1090));
  bfr _b_11990(.a(_w_13892),.q(_w_13893));
  bfr _b_4439(.a(_w_6341),.q(n1113_1));
  bfr _b_7688(.a(_w_9590),.q(_w_9591));
  spl2 g892_s_0(.a(n892),.q0(n892_0),.q1(n892_1));
  bfr _b_6301(.a(_w_8203),.q(n1660));
  bfr _b_12734(.a(_w_14636),.q(_w_14637));
  bfr _b_8904(.a(_w_10806),.q(_w_10807));
  bfr _b_6303(.a(_w_8205),.q(n1081));
  bfr _b_6304(.a(_w_8206),.q(n407));
  bfr _b_9074(.a(_w_10976),.q(_w_10977));
  and_bb g1171(.a(N120_15),.b(N460_11),.q(_w_11069));
  bfr _b_6305(.a(_w_8207),.q(n1648));
  bfr _b_4113(.a(_w_6015),.q(_w_6016));
  bfr _b_7213(.a(_w_9115),.q(_w_9116));
  bfr _b_4710(.a(_w_6612),.q(_w_6613));
  and_bi g350(.a(n348_0),.b(n349),.q(n350));
  bfr _b_9276(.a(_w_11178),.q(_w_11179));
  bfr _b_13510(.a(_w_15412),.q(_w_15413));
  bfr _b_6309(.a(_w_8211),.q(_w_8212));
  bfr _b_8566(.a(_w_10468),.q(_w_10469));
  bfr _b_8102(.a(_w_10004),.q(_w_10005));
  bfr _b_12868(.a(_w_14770),.q(n1885));
  bfr _b_6311(.a(_w_8213),.q(_w_8214));
  bfr _b_6312(.a(_w_8214),.q(_w_8215));
  bfr _b_6315(.a(_w_8217),.q(_w_8218));
  bfr _b_12736(.a(_w_14638),.q(_w_14639));
  bfr _b_6317(.a(_w_8219),.q(n917_1));
  bfr _b_6943(.a(_w_8845),.q(_w_8846));
  bfr _b_5053(.a(_w_6955),.q(_w_6956));
  bfr _b_6318(.a(_w_8220),.q(_w_8221));
  bfr _b_6319(.a(_w_8221),.q(_w_8222));
  bfr _b_6322(.a(_w_8224),.q(_w_8225));
  bfr _b_8571(.a(_w_10473),.q(_w_10474));
  bfr _b_10703(.a(_w_12605),.q(_w_12606));
  bfr _b_3425(.a(_w_5327),.q(_w_5328));
  bfr _b_6324(.a(_w_8226),.q(_w_8227));
  bfr _b_12405(.a(_w_14307),.q(n1766));
  bfr _b_7146(.a(_w_9048),.q(_w_9049));
  bfr _b_6325(.a(_w_8227),.q(n1242_1));
  bfr _b_8177(.a(_w_10079),.q(_w_10080));
  bfr _b_6328(.a(_w_8230),.q(_w_8231));
  spl2 g690_s_0(.a(n690),.q0(n690_0),.q1(n690_1));
  bfr _b_6480(.a(_w_8382),.q(_w_8383));
  spl2 g213_s_0(.a(n213),.q0(n213_0),.q1(n213_1));
  bfr _b_6329(.a(_w_8231),.q(_w_8232));
  bfr _b_7197(.a(_w_9099),.q(_w_9100));
  bfr _b_6330(.a(_w_8232),.q(_w_8233));
  bfr _b_6332(.a(_w_8234),.q(_w_8235));
  bfr _b_6335(.a(_w_8237),.q(_w_8238));
  bfr _b_7662(.a(_w_9564),.q(_w_9565));
  bfr _b_6336(.a(_w_8238),.q(_w_8239));
  bfr _b_6585(.a(_w_8487),.q(_w_8488));
  bfr _b_6337(.a(_w_8239),.q(_w_8240));
  bfr _b_8666(.a(_w_10568),.q(_w_10569));
  bfr _b_10579(.a(_w_12481),.q(_w_12482));
  and_bb g565(.a(n535_1),.b(n563_1),.q(_w_11108));
  bfr _b_6338(.a(_w_8240),.q(_w_8241));
  bfr _b_6339(.a(_w_8241),.q(_w_8242));
  bfr _b_6342(.a(_w_8244),.q(_w_8245));
  bfr _b_3406(.a(_w_5308),.q(_w_5309));
  bfr _b_6345(.a(_w_8247),.q(_w_8248));
  bfr _b_14311(.a(_w_16213),.q(_w_16214));
  bfr _b_4262(.a(_w_6164),.q(n1010_1));
  bfr _b_9052(.a(_w_10954),.q(n254));
  bfr _b_6346(.a(_w_8248),.q(_w_8249));
  bfr _b_3845(.a(_w_5747),.q(_w_5748));
  bfr _b_6347(.a(_w_8249),.q(_w_8250));
  bfr _b_10085(.a(_w_11987),.q(_w_11988));
  bfr _b_4969(.a(_w_6871),.q(_w_6872));
  bfr _b_6348(.a(_w_8250),.q(_w_8251));
  bfr _b_6352(.a(_w_8254),.q(_w_8255));
  bfr _b_12028(.a(_w_13930),.q(_w_13931));
  bfr _b_10424(.a(_w_12326),.q(_w_12327));
  bfr _b_8424(.a(_w_10326),.q(_w_10327));
  bfr _b_8974(.a(_w_10876),.q(_w_10877));
  bfr _b_12169(.a(_w_14071),.q(_w_14072));
  bfr _b_6355(.a(_w_8257),.q(_w_8258));
  bfr _b_6356(.a(_w_8258),.q(_w_8259));
  spl2 g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1));
  bfr _b_6357(.a(_w_8259),.q(_w_8260));
  bfr _b_9632(.a(_w_11534),.q(_w_11535));
  bfr _b_6359(.a(_w_8261),.q(_w_8262));
  bfr _b_6744(.a(_w_8646),.q(_w_8647));
  bfr _b_6360(.a(_w_8262),.q(_w_8263));
  bfr _b_13927(.a(_w_15829),.q(_w_15830));
  bfr _b_6361(.a(_w_8263),.q(_w_8264));
  bfr _b_6366(.a(_w_8268),.q(_w_8269));
  bfr _b_7336(.a(_w_9238),.q(_w_9239));
  bfr _b_5439(.a(_w_7341),.q(_w_7342));
  bfr _b_6367(.a(_w_8269),.q(_w_8270));
  bfr _b_6370(.a(_w_8272),.q(n1869));
  bfr _b_6371(.a(_w_8273),.q(_w_8274));
  or_bb g1515(.a(n1457_0),.b(n1514_0),.q(n1515));
  bfr _b_6372(.a(_w_8274),.q(_w_8275));
  spl2 g1886_s_0(.a(n1886),.q0(n1886_0),.q1(n1886_1));
  bfr _b_6373(.a(_w_8275),.q(_w_8276));
  bfr _b_6374(.a(_w_8276),.q(_w_8277));
  bfr _b_10812(.a(_w_12714),.q(_w_12715));
  bfr _b_6377(.a(_w_8279),.q(_w_8280));
  bfr _b_9503(.a(_w_11405),.q(n509));
  bfr _b_6378(.a(_w_8280),.q(_w_8281));
  bfr _b_6380(.a(_w_8282),.q(_w_8283));
  bfr _b_6381(.a(_w_8283),.q(_w_8284));
  bfr _b_6384(.a(_w_8286),.q(_w_8287));
  bfr _b_7920(.a(_w_9822),.q(_w_9823));
  bfr _b_6385(.a(_w_8287),.q(_w_8288));
  bfr _b_6387(.a(_w_8289),.q(_w_8290));
  bfr _b_13254(.a(_w_15156),.q(_w_15157));
  bfr _b_8334(.a(_w_10236),.q(_w_10237));
  bfr _b_13774(.a(_w_15676),.q(_w_15677));
  bfr _b_6389(.a(_w_8291),.q(_w_8292));
  bfr _b_6392(.a(_w_8294),.q(_w_8295));
  bfr _b_6393(.a(_w_8295),.q(_w_8296));
  bfr _b_6396(.a(_w_8298),.q(_w_8299));
  bfr _b_6398(.a(_w_8300),.q(_w_8301));
  bfr _b_6399(.a(_w_8301),.q(_w_8302));
  bfr _b_14366(.a(_w_16268),.q(_w_16269));
  bfr _b_6969(.a(_w_8871),.q(_w_8872));
  bfr _b_6401(.a(_w_8303),.q(_w_8304));
  bfr _b_6404(.a(_w_8306),.q(_w_8307));
  bfr _b_6217(.a(_w_8119),.q(_w_8120));
  bfr _b_6410(.a(_w_8312),.q(_w_8313));
  bfr _b_12573(.a(_w_14475),.q(_w_14476));
  bfr _b_6411(.a(_w_8313),.q(_w_8314));
  bfr _b_6412(.a(_w_8314),.q(_w_8315));
  bfr _b_7502(.a(_w_9404),.q(_w_9405));
  bfr _b_6279(.a(_w_8181),.q(n260));
  bfr _b_6413(.a(_w_8315),.q(_w_8316));
  bfr _b_11762(.a(_w_13664),.q(_w_13665));
  bfr _b_6414(.a(_w_8316),.q(_w_8317));
  bfr _b_8712(.a(_w_10614),.q(_w_10615));
  spl2 g1437_s_0(.a(n1437),.q0(n1437_0),.q1(n1437_1));
  bfr _b_9897(.a(_w_11799),.q(_w_11800));
  bfr _b_6416(.a(_w_8318),.q(_w_8319));
  bfr _b_8375(.a(_w_10277),.q(_w_10278));
  bfr _b_6417(.a(_w_8319),.q(_w_8320));
  bfr _b_10762(.a(_w_12664),.q(_w_12665));
  bfr _b_7022(.a(_w_8924),.q(N5971));
  bfr _b_6418(.a(_w_8320),.q(_w_8321));
  bfr _b_7725(.a(_w_9627),.q(_w_9628));
  bfr _b_6422(.a(_w_8324),.q(_w_8325));
  bfr _b_10216(.a(_w_12118),.q(_w_12119));
  bfr _b_10090(.a(_w_11992),.q(_w_11993));
  bfr _b_5164(.a(_w_7066),.q(_w_7067));
  bfr _b_6423(.a(_w_8325),.q(_w_8326));
  bfr _b_6776(.a(_w_8678),.q(_w_8679));
  bfr _b_9036(.a(_w_10938),.q(_w_10939));
  spl2 g1514_s_0(.a(n1514),.q0(n1514_0),.q1(n1514_1));
  bfr _b_6427(.a(_w_8329),.q(_w_8330));
  bfr _b_6428(.a(_w_8330),.q(_w_8331));
  bfr _b_6434(.a(_w_8336),.q(_w_8337));
  bfr _b_11672(.a(_w_13574),.q(_w_13575));
  bfr _b_6436(.a(_w_8338),.q(_w_8339));
  bfr _b_11819(.a(_w_13721),.q(_w_13722));
  bfr _b_6887(.a(_w_8789),.q(_w_8790));
  bfr _b_9054(.a(_w_10956),.q(_w_10957));
  bfr _b_7828(.a(_w_9730),.q(_w_9731));
  bfr _b_6437(.a(_w_8339),.q(_w_8340));
  bfr _b_6440(.a(_w_8342),.q(_w_8343));
  bfr _b_6441(.a(_w_8343),.q(_w_8344));
  bfr _b_6443(.a(_w_8345),.q(_w_8346));
  bfr _b_5081(.a(_w_6983),.q(_w_6984));
  bfr _b_6444(.a(_w_8346),.q(_w_8347));
  bfr _b_6686(.a(_w_8588),.q(_w_8589));
  bfr _b_6446(.a(_w_8348),.q(_w_8349));
  bfr _b_8735(.a(_w_10637),.q(_w_10638));
  bfr _b_12276(.a(_w_14178),.q(_w_14179));
  bfr _b_6448(.a(_w_8350),.q(_w_8351));
  bfr _b_10088(.a(_w_11990),.q(_w_11991));
  bfr _b_6449(.a(_w_8351),.q(_w_8352));
  bfr _b_6450(.a(_w_8352),.q(_w_8353));
  bfr _b_3620(.a(_w_5522),.q(_w_5523));
  bfr _b_6156(.a(_w_8058),.q(_w_8059));
  bfr _b_6452(.a(_w_8354),.q(_w_8355));
  spl2 g657_s_0(.a(n657),.q0(n657_0),.q1(n657_1));
  bfr _b_8455(.a(_w_10357),.q(_w_10358));
  bfr _b_9401(.a(_w_11303),.q(_w_11304));
  bfr _b_6458(.a(_w_8360),.q(n1029));
  bfr _b_6459(.a(_w_8361),.q(n1005));
  bfr _b_7311(.a(_w_9213),.q(_w_9214));
  bfr _b_14270(.a(_w_16172),.q(_w_16173));
  and_bi g1115(.a(n1113_0),.b(n1114),.q(n1115));
  bfr _b_6460(.a(_w_8362),.q(n1002));
  or_bb g1557(.a(n1555_0),.b(n1556),.q(n1557));
  bfr _b_6461(.a(_w_8363),.q(n999));
  bfr _b_6462(.a(_w_8364),.q(_w_8365));
  bfr _b_6466(.a(_w_8368),.q(n990));
  bfr _b_5189(.a(_w_7091),.q(_w_7092));
  bfr _b_6468(.a(_w_8370),.q(_w_8371));
  bfr _b_14289(.a(_w_16191),.q(_w_16192));
  bfr _b_6469(.a(_w_8371),.q(_w_8372));
  and_bb g1618(.a(N222_10),.b(N443_17),.q(_w_13966));
  bfr _b_6470(.a(_w_8372),.q(n967));
  bfr _b_6471(.a(_w_8373),.q(_w_8374));
  bfr _b_7274(.a(_w_9176),.q(n734));
  bfr _b_10939(.a(_w_12841),.q(_w_12842));
  bfr _b_6473(.a(_w_8375),.q(_w_8376));
  bfr _b_6014(.a(_w_7916),.q(_w_7917));
  bfr _b_6477(.a(_w_8379),.q(_w_8380));
  bfr _b_6113(.a(_w_8015),.q(_w_8016));
  bfr _b_6479(.a(_w_8381),.q(_w_8382));
  bfr _b_6481(.a(_w_8383),.q(n964));
  and_bi g1135(.a(n1056_1),.b(n1133_1),.q(_w_13204));
  bfr _b_9595(.a(_w_11497),.q(_w_11498));
  and_bb g738(.a(n637_1),.b(n737_0),.q(n738));
  bfr _b_6482(.a(_w_8384),.q(n1708));
  and_bi g223(.a(n222_0),.b(n182_0),.q(n223));
  bfr _b_8933(.a(_w_10835),.q(_w_10836));
  bfr _b_6484(.a(_w_8386),.q(_w_8387));
  bfr _b_6485(.a(_w_8387),.q(_w_8388));
  bfr _b_6488(.a(_w_8390),.q(n290));
  bfr _b_6490(.a(_w_8392),.q(_w_8393));
  bfr _b_6491(.a(_w_8393),.q(_w_8394));
  spl4L N18_s_1(.a(N18_0),.q0(N18_4),.q1(N18_5),.q2(_w_15485),.q3(_w_15487));
  bfr _b_6492(.a(_w_8394),.q(_w_8395));
  bfr _b_6493(.a(_w_8395),.q(_w_8396));
  bfr _b_6494(.a(_w_8396),.q(_w_8397));
  bfr _b_6496(.a(_w_8398),.q(_w_8399));
  bfr _b_8906(.a(_w_10808),.q(_w_10809));
  bfr _b_6498(.a(_w_8400),.q(_w_8401));
  bfr _b_12511(.a(_w_14413),.q(_w_14414));
  bfr _b_6885(.a(_w_8787),.q(_w_8788));
  bfr _b_7256(.a(_w_9158),.q(_w_9159));
  bfr _b_6500(.a(_w_8402),.q(_w_8403));
  bfr _b_6501(.a(_w_8403),.q(_w_8404));
  bfr _b_8112(.a(_w_10014),.q(_w_10015));
  bfr _b_10428(.a(_w_12330),.q(_w_12331));
  bfr _b_4610(.a(_w_6512),.q(_w_6513));
  bfr _b_6503(.a(_w_8405),.q(_w_8406));
  bfr _b_6506(.a(_w_8408),.q(_w_8409));
  bfr _b_6508(.a(_w_8410),.q(_w_8411));
  bfr _b_5806(.a(_w_7708),.q(_w_7709));
  bfr _b_6510(.a(_w_8412),.q(_w_8413));
  bfr _b_9093(.a(_w_10995),.q(_w_10996));
  bfr _b_12205(.a(_w_14107),.q(n879));
  bfr _b_11470(.a(_w_13372),.q(n1325));
  bfr _b_6513(.a(_w_8415),.q(_w_8416));
  spl2 g1728_s_0(.a(n1728),.q0(n1728_0),.q1(n1728_1));
  bfr _b_6516(.a(_w_8418),.q(_w_8419));
  and_bb g832(.a(N103_13),.b(N426_10),.q(n832));
  bfr _b_5584(.a(_w_7486),.q(N69_13));
  bfr _b_6519(.a(_w_8421),.q(_w_8422));
  bfr _b_9882(.a(_w_11784),.q(_w_11785));
  bfr _b_6520(.a(_w_8422),.q(_w_8423));
  bfr _b_6521(.a(_w_8423),.q(_w_8424));
  bfr _b_6524(.a(_w_8426),.q(_w_8427));
  bfr _b_6594(.a(_w_8496),.q(_w_8497));
  bfr _b_8921(.a(_w_10823),.q(_w_10824));
  bfr _b_6526(.a(_w_8428),.q(_w_8429));
  bfr _b_6527(.a(_w_8429),.q(_w_8430));
  bfr _b_6529(.a(_w_8431),.q(_w_8432));
  bfr _b_6530(.a(_w_8432),.q(_w_8433));
  bfr _b_13923(.a(_w_15825),.q(_w_15826));
  bfr _b_6534(.a(_w_8436),.q(_w_8437));
  bfr _b_6535(.a(_w_8437),.q(_w_8438));
  bfr _b_13907(.a(_w_15809),.q(_w_15810));
  and_bi g1234(.a(n1171_1),.b(n1232_1),.q(_w_13010));
  bfr _b_6536(.a(_w_8438),.q(_w_8439));
  bfr _b_7359(.a(_w_9261),.q(n656));
  bfr _b_6537(.a(_w_8439),.q(_w_8440));
  bfr _b_6539(.a(_w_8441),.q(_w_8442));
  bfr _b_6541(.a(_w_8443),.q(_w_8444));
  bfr _b_6542(.a(_w_8444),.q(_w_8445));
  bfr _b_6547(.a(_w_8449),.q(_w_8450));
  bfr _b_7809(.a(_w_9711),.q(_w_9712));
  bfr _b_6548(.a(_w_8450),.q(_w_8451));
  bfr _b_6549(.a(_w_8451),.q(_w_8452));
  bfr _b_6553(.a(_w_8455),.q(_w_8456));
  bfr _b_6554(.a(_w_8456),.q(_w_8457));
  bfr _b_6796(.a(_w_8698),.q(_w_8699));
  bfr _b_5498(.a(_w_7400),.q(_w_7401));
  spl2 g1357_s_0(.a(n1357),.q0(n1357_0),.q1(_w_8024));
  bfr _b_6555(.a(_w_8457),.q(_w_8458));
  bfr _b_6556(.a(_w_8458),.q(_w_8459));
  bfr _b_6558(.a(_w_8460),.q(_w_8461));
  and_bi g510(.a(n508_0),.b(n509),.q(n510));
  bfr _b_6559(.a(_w_8461),.q(_w_8462));
  bfr _b_6560(.a(_w_8462),.q(_w_8463));
  bfr _b_4890(.a(_w_6792),.q(_w_6793));
  bfr _b_6561(.a(_w_8463),.q(_w_8464));
  and_bb g251(.a(n192_2),.b(n249_1),.q(_w_12490));
  bfr _b_6593(.a(_w_8495),.q(_w_8496));
  bfr _b_6562(.a(_w_8464),.q(_w_8465));
  bfr _b_12726(.a(_w_14628),.q(_w_14629));
  bfr _b_6566(.a(_w_8468),.q(_w_8469));
  bfr _b_7939(.a(_w_9841),.q(_w_9842));
  bfr _b_6571(.a(_w_8473),.q(_w_8474));
  bfr _b_6573(.a(_w_8475),.q(_w_8476));
  bfr _b_6574(.a(_w_8476),.q(_w_8477));
  bfr _b_6576(.a(_w_8478),.q(_w_8479));
  or_bb g693(.a(n691_0),.b(n692),.q(n693));
  bfr _b_6579(.a(_w_8481),.q(_w_8482));
  bfr _b_11500(.a(_w_13402),.q(_w_13403));
  bfr _b_6407(.a(_w_8309),.q(_w_8310));
  bfr _b_9896(.a(_w_11798),.q(_w_11799));
  bfr _b_4773(.a(_w_6675),.q(_w_6676));
  bfr _b_9892(.a(_w_11794),.q(_w_11795));
  bfr _b_6581(.a(_w_8483),.q(_w_8484));
  spl2 g1724_s_0(.a(n1724),.q0(n1724_0),.q1(n1724_1));
  bfr _b_6582(.a(_w_8484),.q(_w_8485));
  bfr _b_5729(.a(_w_7631),.q(N222_8));
  bfr _b_6583(.a(_w_8485),.q(_w_8486));
  bfr _b_12731(.a(_w_14633),.q(_w_14634));
  bfr _b_6588(.a(_w_8490),.q(_w_8491));
  and_bi g1718(.a(n1716_0),.b(n1717),.q(n1718));
  bfr _b_6425(.a(_w_8327),.q(_w_8328));
  bfr _b_6928(.a(_w_8830),.q(_w_8831));
  bfr _b_6589(.a(_w_8491),.q(_w_8492));
  bfr _b_6592(.a(_w_8494),.q(_w_8495));
  bfr _b_6595(.a(_w_8497),.q(_w_8498));
  bfr _b_9750(.a(_w_11652),.q(_w_11653));
  bfr _b_5492(.a(_w_7394),.q(_w_7395));
  bfr _b_6596(.a(_w_8498),.q(_w_8499));
  bfr _b_6599(.a(_w_8501),.q(_w_8502));
  bfr _b_6600(.a(_w_8502),.q(_w_8503));
  bfr _b_10591(.a(_w_12493),.q(_w_12494));
  bfr _b_6603(.a(_w_8505),.q(_w_8506));
  bfr _b_7370(.a(_w_9272),.q(_w_9273));
  bfr _b_13994(.a(_w_15896),.q(_w_15897));
  bfr _b_9589(.a(_w_11491),.q(_w_11492));
  bfr _b_6604(.a(_w_8506),.q(_w_8507));
  bfr _b_6979(.a(_w_8881),.q(_w_8882));
  bfr _b_8671(.a(_w_10573),.q(n473));
  bfr _b_6237(.a(_w_8139),.q(_w_8140));
  bfr _b_6379(.a(_w_8281),.q(_w_8282));
  bfr _b_9040(.a(_w_10942),.q(_w_10943));
  bfr _b_6606(.a(_w_8508),.q(_w_8509));
  bfr _b_7299(.a(_w_9201),.q(n712));
  bfr _b_10965(.a(_w_12867),.q(_w_12868));
  bfr _b_5297(.a(_w_7199),.q(_w_7200));
  bfr _b_6607(.a(_w_8509),.q(_w_8510));
  bfr _b_6608(.a(_w_8510),.q(_w_8511));
  bfr _b_6609(.a(_w_8511),.q(_w_8512));
  bfr _b_6610(.a(_w_8512),.q(_w_8513));
  bfr _b_8940(.a(_w_10842),.q(n1375));
  bfr _b_6611(.a(_w_8513),.q(_w_8514));
  spl2 g1659_s_0(.a(n1659),.q0(n1659_0),.q1(_w_9257));
  bfr _b_7909(.a(_w_9811),.q(_w_9812));
  bfr _b_6613(.a(_w_8515),.q(_w_8516));
  bfr _b_13836(.a(_w_15738),.q(_w_15739));
  or_bb g1248(.a(n1166_0),.b(n1247_0),.q(n1248));
  bfr _b_7305(.a(_w_9207),.q(n720));
  bfr _b_13290(.a(_w_15192),.q(_w_15193));
  bfr _b_6614(.a(_w_8516),.q(_w_8517));
  bfr _b_6616(.a(_w_8518),.q(_w_8519));
  bfr _b_6778(.a(_w_8680),.q(_w_8681));
  bfr _b_12262(.a(_w_14164),.q(_w_14165));
  bfr _b_9723(.a(_w_11625),.q(_w_11626));
  bfr _b_6618(.a(_w_8520),.q(_w_8521));
  bfr _b_13850(.a(_w_15752),.q(_w_15753));
  bfr _b_13401(.a(_w_15303),.q(n1206_1));
  bfr _b_6755(.a(_w_8657),.q(_w_8658));
  bfr _b_6619(.a(_w_8521),.q(_w_8522));
  bfr _b_13145(.a(_w_15047),.q(n1515_1));
  bfr _b_10985(.a(_w_12887),.q(n1268));
  bfr _b_6620(.a(_w_8522),.q(_w_8523));
  bfr _b_6621(.a(_w_8523),.q(_w_8524));
  bfr _b_11771(.a(_w_13673),.q(_w_13674));
  bfr _b_7966(.a(_w_9868),.q(_w_9869));
  bfr _b_12499(.a(_w_14401),.q(_w_14402));
  bfr _b_6622(.a(_w_8524),.q(_w_8525));
  and_bi g1215(.a(n1214_0),.b(n1177_0),.q(n1215));
  bfr _b_6623(.a(_w_8525),.q(_w_8526));
  bfr _b_8944(.a(_w_10846),.q(_w_10847));
  bfr _b_8056(.a(_w_9958),.q(n67));
  bfr _b_6624(.a(_w_8526),.q(_w_8527));
  bfr _b_3577(.a(_w_5479),.q(_w_5480));
  bfr _b_4877(.a(_w_6779),.q(_w_6780));
  spl2 g796_s_0(.a(n796),.q0(n796_0),.q1(_w_7058));
  or_bb g1670(.a(n1668_0),.b(n1669),.q(_w_14010));
  bfr _b_6626(.a(_w_8528),.q(_w_8529));
  bfr _b_6627(.a(_w_8529),.q(_w_8530));
  bfr _b_6628(.a(_w_8530),.q(_w_8531));
  bfr _b_6633(.a(_w_8535),.q(_w_8536));
  bfr _b_6634(.a(_w_8536),.q(_w_8537));
  bfr _b_9004(.a(_w_10906),.q(_w_10907));
  bfr _b_12049(.a(_w_13951),.q(n975));
  bfr _b_5720(.a(_w_7622),.q(_w_7623));
  bfr _b_9660(.a(_w_11562),.q(_w_11563));
  bfr _b_6636(.a(_w_8538),.q(_w_8539));
  bfr _b_6637(.a(_w_8539),.q(_w_8540));
  bfr _b_6638(.a(_w_8540),.q(_w_8541));
  bfr _b_11650(.a(_w_13552),.q(_w_13553));
  bfr _b_6888(.a(_w_8790),.q(_w_8791));
  or_bb g986(.a(n955_0),.b(n985_0),.q(n986));
  bfr _b_6639(.a(_w_8541),.q(_w_8542));
  bfr _b_10727(.a(_w_12629),.q(_w_12630));
  bfr _b_6640(.a(_w_8542),.q(_w_8543));
  spl2 g167_s_0(.a(n167),.q0(n167_0),.q1(n167_1));
  bfr _b_6641(.a(_w_8543),.q(_w_8544));
  bfr _b_6642(.a(_w_8544),.q(_w_8545));
  bfr _b_6643(.a(_w_8545),.q(_w_8546));
  bfr _b_12493(.a(_w_14395),.q(_w_14396));
  bfr _b_6645(.a(_w_8547),.q(_w_8548));
  spl2 g1236_s_0(.a(n1236),.q0(n1236_0),.q1(_w_14977));
  bfr _b_6648(.a(_w_8550),.q(_w_8551));
  bfr _b_6649(.a(_w_8551),.q(_w_8552));
  bfr _b_9879(.a(_w_11781),.q(_w_11782));
  bfr _b_6651(.a(_w_8553),.q(_w_8554));
  and_bi g1556(.a(n1549_1),.b(n1554_1),.q(_w_13932));
  bfr _b_6653(.a(_w_8555),.q(_w_8556));
  bfr _b_6656(.a(_w_8558),.q(N205_3));
  bfr _b_6658(.a(_w_8560),.q(_w_8561));
  bfr _b_6659(.a(_w_8561),.q(_w_8562));
  bfr _b_10235(.a(_w_12137),.q(_w_12138));
  bfr _b_12191(.a(_w_14093),.q(_w_14094));
  bfr _b_6661(.a(_w_8563),.q(n262_1));
  and_bi g1482(.a(n1481_0),.b(n1468_0),.q(n1482));
  bfr _b_6666(.a(_w_8568),.q(_w_8569));
  bfr _b_9032(.a(_w_10934),.q(_w_10935));
  bfr _b_7501(.a(_w_9403),.q(_w_9404));
  bfr _b_6667(.a(_w_8569),.q(_w_8570));
  bfr _b_12750(.a(_w_14652),.q(_w_14653));
  bfr _b_8027(.a(_w_9929),.q(_w_9930));
  bfr _b_6670(.a(_w_8572),.q(_w_8573));
  bfr _b_7324(.a(_w_9226),.q(n686));
  and_bi g1534(.a(n1521_1),.b(n1524_1),.q(n1534));
  bfr _b_6402(.a(_w_8304),.q(_w_8305));
  bfr _b_6671(.a(_w_8573),.q(_w_8574));
  bfr _b_6675(.a(_w_8577),.q(_w_8578));
  and_bb g1156(.a(n1049_1),.b(n1154_1),.q(_w_12863));
  bfr _b_6676(.a(_w_8578),.q(n374));
  bfr _b_12498(.a(_w_14400),.q(_w_14401));
  bfr _b_4453(.a(_w_6355),.q(_w_6356));
  bfr _b_6678(.a(_w_8580),.q(_w_8581));
  bfr _b_6680(.a(_w_8582),.q(_w_8583));
  bfr _b_9069(.a(_w_10971),.q(_w_10972));
  bfr _b_10059(.a(_w_11961),.q(_w_11962));
  bfr _b_6681(.a(_w_8583),.q(_w_8584));
  bfr _b_11809(.a(_w_13711),.q(_w_13712));
  and_bi g311(.a(n310),.b(n308_0),.q(n311));
  bfr _b_7298(.a(_w_9200),.q(_w_9201));
  bfr _b_8817(.a(_w_10719),.q(_w_10720));
  bfr _b_6683(.a(_w_8585),.q(_w_8586));
  bfr _b_8200(.a(_w_10102),.q(_w_10103));
  bfr _b_6685(.a(_w_8587),.q(_w_8588));
  bfr _b_6687(.a(_w_8589),.q(_w_8590));
  bfr _b_9961(.a(_w_11863),.q(_w_11864));
  bfr _b_6688(.a(_w_8590),.q(_w_8591));
  bfr _b_6689(.a(_w_8591),.q(_w_8592));
  bfr _b_10999(.a(_w_12901),.q(_w_12902));
  bfr _b_5313(.a(_w_7215),.q(_w_7216));
  bfr _b_6806(.a(_w_8708),.q(_w_8709));
  bfr _b_7949(.a(_w_9851),.q(_w_9852));
  bfr _b_9680(.a(_w_11582),.q(_w_11583));
  bfr _b_9594(.a(_w_11496),.q(_w_11497));
  bfr _b_6690(.a(_w_8592),.q(_w_8593));
  bfr _b_10510(.a(_w_12412),.q(_w_12413));
  bfr _b_7399(.a(_w_9301),.q(_w_9302));
  bfr _b_8057(.a(_w_9959),.q(n386));
  bfr _b_6693(.a(_w_8595),.q(_w_8596));
  bfr _b_6694(.a(_w_8596),.q(_w_8597));
  bfr _b_11740(.a(_w_13642),.q(_w_13643));
  bfr _b_6697(.a(_w_8599),.q(_w_8600));
  bfr _b_9217(.a(_w_11119),.q(_w_11120));
  bfr _b_6699(.a(_w_8601),.q(_w_8602));
  bfr _b_14361(.a(_w_16263),.q(_w_16264));
  bfr _b_6700(.a(_w_8602),.q(_w_8603));
  bfr _b_9997(.a(_w_11899),.q(_w_11900));
  bfr _b_6701(.a(_w_8603),.q(_w_8604));
  bfr _b_6705(.a(_w_8607),.q(_w_8608));
  bfr _b_12125(.a(_w_14027),.q(_w_14028));
  bfr _b_9112(.a(_w_11014),.q(n552_1));
  bfr _b_3648(.a(_w_5550),.q(n1635_1));
  bfr _b_6706(.a(_w_8608),.q(_w_8609));
  or_bb g753(.a(n751_0),.b(n752),.q(n753));
  bfr _b_6708(.a(_w_8610),.q(_w_8611));
  bfr _b_6709(.a(_w_8611),.q(_w_8612));
  bfr _b_9148(.a(_w_11050),.q(_w_11051));
  bfr _b_7464(.a(_w_9366),.q(_w_9367));
  bfr _b_6710(.a(_w_8612),.q(_w_8613));
  bfr _b_6723(.a(_w_8625),.q(_w_8626));
  bfr _b_9219(.a(_w_11121),.q(_w_11122));
  bfr _b_10505(.a(_w_12407),.q(_w_12408));
  and_bi g84(.a(n82_0),.b(n83),.q(n84));
  bfr _b_6711(.a(_w_8613),.q(_w_8614));
  bfr _b_9593(.a(_w_11495),.q(_w_11496));
  spl2 g345_s_0(.a(n345),.q0(n345_0),.q1(n345_1));
  bfr _b_6712(.a(_w_8614),.q(_w_8615));
  bfr _b_6713(.a(_w_8615),.q(_w_8616));
  bfr _b_7557(.a(_w_9459),.q(_w_9460));
  bfr _b_8773(.a(_w_10675),.q(_w_10676));
  bfr _b_6714(.a(_w_8616),.q(_w_8617));
  bfr _b_12236(.a(_w_14138),.q(_w_14139));
  bfr _b_10419(.a(_w_12321),.q(_w_12322));
  bfr _b_6715(.a(_w_8617),.q(_w_8618));
  spl2 g321_s_0(.a(n321),.q0(n321_0),.q1(n321_1));
  bfr _b_6717(.a(_w_8619),.q(_w_8620));
  bfr _b_4659(.a(_w_6561),.q(_w_6562));
  bfr _b_6106(.a(_w_8008),.q(_w_8009));
  bfr _b_9810(.a(_w_11712),.q(_w_11713));
  bfr _b_10140(.a(_w_12042),.q(_w_12043));
  bfr _b_10241(.a(_w_12143),.q(_w_12144));
  bfr _b_6719(.a(_w_8621),.q(_w_8622));
  bfr _b_11475(.a(_w_13377),.q(_w_13378));
  bfr _b_10021(.a(_w_11923),.q(_w_11924));
  bfr _b_6720(.a(_w_8622),.q(_w_8623));
  bfr _b_6721(.a(_w_8623),.q(_w_8624));
  bfr _b_9413(.a(_w_11315),.q(_w_11316));
  bfr _b_6727(.a(_w_8629),.q(_w_8630));
  bfr _b_3488(.a(_w_5390),.q(_w_5391));
  bfr _b_6429(.a(_w_8331),.q(_w_8332));
  bfr _b_6944(.a(_w_8846),.q(_w_8847));
  bfr _b_6729(.a(_w_8631),.q(_w_8632));
  bfr _b_6731(.a(_w_8633),.q(_w_8634));
  bfr _b_3527(.a(_w_5429),.q(_w_5430));
  bfr _b_6733(.a(_w_8635),.q(_w_8636));
  spl2 g232_s_0(.a(n232),.q0(n232_0),.q1(n232_1));
  bfr _b_6736(.a(_w_8638),.q(_w_8639));
  bfr _b_6737(.a(_w_8639),.q(_w_8640));
  bfr _b_6105(.a(_w_8007),.q(_w_8008));
  bfr _b_6740(.a(_w_8642),.q(_w_8643));
  bfr _b_11526(.a(_w_13428),.q(_w_13429));
  bfr _b_6741(.a(_w_8643),.q(_w_8644));
  spl2 g273_s_0(.a(n273),.q0(n273_0),.q1(n273_1));
  bfr _b_6742(.a(_w_8644),.q(_w_8645));
  bfr _b_6743(.a(_w_8645),.q(_w_8646));
  bfr _b_6745(.a(_w_8647),.q(_w_8648));
  bfr _b_11408(.a(_w_13310),.q(_w_13311));
  bfr _b_6746(.a(_w_8648),.q(_w_8649));
  bfr _b_6747(.a(_w_8649),.q(_w_8650));
  bfr _b_9339(.a(_w_11241),.q(_w_11242));
  bfr _b_11854(.a(_w_13756),.q(n1438));
  bfr _b_6750(.a(_w_8652),.q(_w_8653));
  bfr _b_6753(.a(_w_8655),.q(_w_8656));
  bfr _b_13446(.a(_w_15348),.q(_w_15349));
  bfr _b_12599(.a(_w_14501),.q(_w_14502));
  bfr _b_6759(.a(_w_8661),.q(_w_8662));
  spl2 g423_s_0(.a(n423),.q0(n423_0),.q1(n423_1));
  bfr _b_7320(.a(_w_9222),.q(_w_9223));
  bfr _b_3599(.a(_w_5501),.q(_w_5502));
  bfr _b_6760(.a(_w_8662),.q(_w_8663));
  bfr _b_3505(.a(_w_5407),.q(_w_5408));
  bfr _b_6761(.a(_w_8663),.q(_w_8664));
  bfr _b_6762(.a(_w_8664),.q(_w_8665));
  bfr _b_6764(.a(_w_8666),.q(_w_8667));
  bfr _b_6767(.a(_w_8669),.q(_w_8670));
  bfr _b_6769(.a(_w_8671),.q(_w_8672));
  bfr _b_6770(.a(_w_8672),.q(_w_8673));
  bfr _b_6771(.a(_w_8673),.q(_w_8674));
  bfr _b_4827(.a(_w_6729),.q(_w_6730));
  bfr _b_4327(.a(_w_6229),.q(_w_6230));
  bfr _b_6773(.a(_w_8675),.q(_w_8676));
  bfr _b_8760(.a(_w_10662),.q(_w_10663));
  bfr _b_13450(.a(_w_15352),.q(_w_15353));
  spl2 g348_s_0(.a(n348),.q0(n348_0),.q1(_w_8131));
  bfr _b_9551(.a(_w_11453),.q(_w_11454));
  bfr _b_5642(.a(_w_7544),.q(_w_7545));
  bfr _b_6777(.a(_w_8679),.q(_w_8680));
  bfr _b_11641(.a(_w_13543),.q(n146_2));
  bfr _b_5882(.a(_w_7784),.q(_w_7785));
  bfr _b_7103(.a(_w_9005),.q(_w_9006));
  bfr _b_6781(.a(_w_8683),.q(_w_8684));
  bfr _b_3985(.a(_w_5887),.q(_w_5888));
  bfr _b_10244(.a(_w_12146),.q(_w_12147));
  bfr _b_6782(.a(_w_8684),.q(_w_8685));
  bfr _b_6783(.a(_w_8685),.q(_w_8686));
  bfr _b_7169(.a(_w_9071),.q(_w_9072));
  bfr _b_6784(.a(_w_8686),.q(_w_8687));
  or_bb g285(.a(n283_0),.b(n284),.q(n285));
  bfr _b_6785(.a(_w_8687),.q(_w_8688));
  bfr _b_6786(.a(_w_8688),.q(_w_8689));
  bfr _b_9120(.a(_w_11022),.q(n574));
  bfr _b_6787(.a(_w_8689),.q(_w_8690));
  bfr _b_13955(.a(_w_15857),.q(_w_15858));
  spl2 g1109_s_0(.a(n1109),.q0(n1109_0),.q1(n1109_1));
  bfr _b_6793(.a(_w_8695),.q(_w_8696));
  bfr _b_11454(.a(_w_13356),.q(_w_13357));
  bfr _b_7079(.a(_w_8981),.q(_w_8982));
  bfr _b_10106(.a(_w_12008),.q(_w_12009));
  bfr _b_6798(.a(_w_8700),.q(N222_14));
  bfr _b_8089(.a(_w_9991),.q(n280_1));
  bfr _b_6799(.a(_w_8701),.q(_w_8702));
  spl2 g1442_s_0(.a(n1442),.q0(n1442_0),.q1(n1442_1));
  bfr _b_6800(.a(_w_8702),.q(_w_8703));
  bfr _b_9356(.a(_w_11258),.q(_w_11259));
  bfr _b_6803(.a(_w_8705),.q(_w_8706));
  bfr _b_11544(.a(_w_13446),.q(n1358));
  bfr _b_3959(.a(_w_5861),.q(_w_5862));
  bfr _b_5894(.a(_w_7796),.q(_w_7797));
  bfr _b_6805(.a(_w_8707),.q(_w_8708));
  bfr _b_9361(.a(_w_11263),.q(_w_11264));
  bfr _b_6807(.a(_w_8709),.q(_w_8710));
  bfr _b_9016(.a(_w_10918),.q(_w_10919));
  bfr _b_6808(.a(_w_8710),.q(_w_8711));
  bfr _b_6809(.a(_w_8711),.q(_w_8712));
  bfr _b_8722(.a(_w_10624),.q(n287));
  bfr _b_3459(.a(_w_5361),.q(_w_5362));
  bfr _b_6810(.a(_w_8712),.q(_w_8713));
  bfr _b_11573(.a(_w_13475),.q(_w_13476));
  bfr _b_7716(.a(_w_9618),.q(_w_9619));
  bfr _b_9267(.a(_w_11169),.q(_w_11170));
  bfr _b_9776(.a(_w_11678),.q(_w_11679));
  bfr _b_3568(.a(_w_5470),.q(_w_5471));
  bfr _b_6812(.a(_w_8714),.q(_w_8715));
  bfr _b_8563(.a(_w_10465),.q(_w_10466));
  bfr _b_11836(.a(_w_13738),.q(_w_13739));
  bfr _b_6814(.a(_w_8716),.q(_w_8717));
  bfr _b_13337(.a(_w_15239),.q(_w_15240));
  spl2 g973_s_0(.a(n973),.q0(n973_0),.q1(n973_1));
  bfr _b_6817(.a(_w_8719),.q(_w_8720));
  bfr _b_6819(.a(_w_8721),.q(_w_8722));
  bfr _b_11340(.a(_w_13242),.q(_w_13243));
  bfr _b_7181(.a(_w_9083),.q(_w_9084));
  bfr _b_6820(.a(_w_8722),.q(_w_8723));
  bfr _b_3609(.a(_w_5511),.q(_w_5512));
  bfr _b_6826(.a(_w_8728),.q(n1078));
  bfr _b_7829(.a(_w_9731),.q(_w_9732));
  bfr _b_6828(.a(_w_8730),.q(n665));
  bfr _b_12275(.a(_w_14177),.q(_w_14178));
  bfr _b_5663(.a(_w_7565),.q(_w_7566));
  bfr _b_6829(.a(_w_8731),.q(_w_8732));
  and_bb g736(.a(N205_6),.b(N307_16),.q(_w_14292));
  bfr _b_6831(.a(_w_8733),.q(_w_8734));
  bfr _b_9047(.a(_w_10949),.q(_w_10950));
  bfr _b_6833(.a(_w_8735),.q(_w_8736));
  bfr _b_11760(.a(_w_13662),.q(_w_13663));
  bfr _b_8946(.a(_w_10848),.q(_w_10849));
  bfr _b_12657(.a(_w_14559),.q(_w_14560));
  bfr _b_11881(.a(_w_13783),.q(_w_13784));
  bfr _b_11138(.a(_w_13040),.q(_w_13041));
  bfr _b_6834(.a(_w_8736),.q(_w_8737));
  bfr _b_6835(.a(_w_8737),.q(_w_8738));
  bfr _b_6836(.a(_w_8738),.q(n1739));
  bfr _b_7515(.a(_w_9417),.q(_w_9418));
  bfr _b_6837(.a(_w_8739),.q(n915));
  bfr _b_6839(.a(_w_8741),.q(_w_8742));
  bfr _b_10753(.a(_w_12655),.q(_w_12656));
  or_bb g94(.a(n73_0),.b(n93_0),.q(n94));
  bfr _b_8380(.a(_w_10282),.q(N5672));
  bfr _b_6840(.a(_w_8742),.q(_w_8743));
  bfr _b_11873(.a(_w_13775),.q(_w_13776));
  spl2 g1218_s_0(.a(n1218),.q0(n1218_0),.q1(_w_11593));
  bfr _b_6841(.a(_w_8743),.q(_w_8744));
  bfr _b_4761(.a(_w_6663),.q(_w_6664));
  bfr _b_6845(.a(_w_8747),.q(n100));
  bfr _b_6847(.a(_w_8749),.q(_w_8750));
  bfr _b_11272(.a(_w_13174),.q(_w_13175));
  bfr _b_10273(.a(_w_12175),.q(_w_12176));
  bfr _b_6848(.a(_w_8750),.q(_w_8751));
  bfr _b_6850(.a(_w_8752),.q(_w_8753));
  bfr _b_11082(.a(_w_12984),.q(_w_12985));
  bfr _b_6851(.a(_w_8753),.q(_w_8754));
  bfr _b_8325(.a(_w_10227),.q(_w_10228));
  bfr _b_6852(.a(_w_8754),.q(_w_8755));
  bfr _b_10997(.a(_w_12899),.q(_w_12900));
  and_bb g1177(.a(N171_12),.b(N409_14),.q(n1177));
  bfr _b_9965(.a(_w_11867),.q(_w_11868));
  bfr _b_6853(.a(_w_8755),.q(_w_8756));
  bfr _b_6854(.a(_w_8756),.q(_w_8757));
  bfr _b_8058(.a(_w_9960),.q(n586));
  bfr _b_8096(.a(_w_9998),.q(_w_9999));
  bfr _b_6857(.a(_w_8759),.q(_w_8760));
  bfr _b_6858(.a(_w_8760),.q(_w_8761));
  bfr _b_9051(.a(_w_10953),.q(N6190));
  bfr _b_6860(.a(_w_8762),.q(_w_8763));
  bfr _b_6861(.a(_w_8763),.q(_w_8764));
  or_bb g904(.a(n902_0),.b(n903),.q(n904));
  bfr _b_6862(.a(_w_8764),.q(n838));
  bfr _b_6864(.a(_w_8766),.q(_w_8767));
  bfr _b_6866(.a(_w_8768),.q(_w_8769));
  bfr _b_6867(.a(_w_8769),.q(_w_8770));
  bfr _b_6868(.a(_w_8770),.q(n846));
  bfr _b_10342(.a(_w_12244),.q(_w_12245));
  bfr _b_6869(.a(_w_8771),.q(n897));
  bfr _b_5241(.a(_w_7143),.q(_w_7144));
  bfr _b_6870(.a(_w_8772),.q(n885));
  bfr _b_6872(.a(_w_8774),.q(n671));
  bfr _b_6873(.a(_w_8775),.q(n1240));
  bfr _b_6876(.a(_w_8778),.q(n864));
  bfr _b_12946(.a(_w_14848),.q(_w_14849));
  bfr _b_6879(.a(_w_8781),.q(_w_8782));
  bfr _b_6881(.a(_w_8783),.q(_w_8784));
  spl2 g1043_s_0(.a(n1043),.q0(n1043_0),.q1(n1043_1));
  bfr _b_6882(.a(_w_8784),.q(n1870_1));
  bfr _b_12047(.a(_w_13949),.q(n1583));
  bfr _b_8341(.a(_w_10243),.q(_w_10244));
  bfr _b_6884(.a(_w_8786),.q(_w_8787));
  bfr _b_6893(.a(_w_8795),.q(_w_8796));
  bfr _b_6889(.a(_w_8791),.q(_w_8792));
  bfr _b_11652(.a(_w_13554),.q(_w_13555));
  bfr _b_7594(.a(_w_9496),.q(_w_9497));
  bfr _b_6891(.a(_w_8793),.q(_w_8794));
  bfr _b_6892(.a(_w_8794),.q(_w_8795));
  or_bb g1839(.a(n1821_0),.b(n1838_0),.q(n1839));
  bfr _b_6895(.a(_w_8797),.q(_w_8798));
  bfr _b_10181(.a(_w_12083),.q(n1173));
  bfr _b_6897(.a(_w_8799),.q(_w_8800));
  and_bb g197(.a(n146_2),.b(n195_1),.q(_w_10627));
  bfr _b_10046(.a(_w_11948),.q(_w_11949));
  bfr _b_13174(.a(_w_15076),.q(_w_15077));
  spl2 g1095_s_0(.a(n1095),.q0(n1095_0),.q1(_w_13864));
  bfr _b_6902(.a(_w_8804),.q(_w_8805));
  bfr _b_6908(.a(_w_8810),.q(_w_8811));
  bfr _b_6910(.a(_w_8812),.q(_w_8813));
  bfr _b_6911(.a(_w_8813),.q(_w_8814));
  bfr _b_6913(.a(_w_8815),.q(_w_8816));
  bfr _b_7123(.a(_w_9025),.q(_w_9026));
  bfr _b_6918(.a(_w_8820),.q(_w_8821));
  bfr _b_8757(.a(_w_10659),.q(_w_10660));
  bfr _b_6922(.a(_w_8824),.q(_w_8825));
  bfr _b_10257(.a(_w_12159),.q(_w_12160));
  bfr _b_11558(.a(_w_13460),.q(_w_13461));
  bfr _b_6925(.a(_w_8827),.q(_w_8828));
  bfr _b_4842(.a(_w_6744),.q(_w_6745));
  bfr _b_6926(.a(_w_8828),.q(_w_8829));
  bfr _b_6927(.a(_w_8829),.q(_w_8830));
  bfr _b_6932(.a(_w_8834),.q(_w_8835));
  bfr _b_6933(.a(_w_8835),.q(_w_8836));
  bfr _b_10664(.a(_w_12566),.q(_w_12567));
  bfr _b_6936(.a(_w_8838),.q(_w_8839));
  bfr _b_7606(.a(_w_9508),.q(_w_9509));
  bfr _b_9519(.a(_w_11421),.q(_w_11422));
  bfr _b_6937(.a(_w_8839),.q(_w_8840));
  bfr _b_12195(.a(_w_14097),.q(_w_14098));
  bfr _b_6938(.a(_w_8840),.q(_w_8841));
  bfr _b_7471(.a(_w_9373),.q(_w_9374));
  bfr _b_6941(.a(_w_8843),.q(_w_8844));
  bfr _b_6942(.a(_w_8844),.q(_w_8845));
  bfr _b_13452(.a(_w_15354),.q(_w_15355));
  bfr _b_6946(.a(_w_8848),.q(_w_8849));
  bfr _b_6947(.a(_w_8849),.q(_w_8850));
  bfr _b_8121(.a(_w_10023),.q(_w_10024));
  bfr _b_11607(.a(_w_13509),.q(_w_13510));
  bfr _b_8845(.a(_w_10747),.q(_w_10748));
  bfr _b_6948(.a(_w_8850),.q(_w_8851));
  bfr _b_6949(.a(_w_8851),.q(_w_8852));
  bfr _b_7371(.a(_w_9273),.q(n1616));
  spl2 g1552_s_0(.a(n1552),.q0(n1552_0),.q1(_w_8364));
  bfr _b_6951(.a(_w_8853),.q(_w_8854));
  bfr _b_6954(.a(_w_8856),.q(N137_11));
  and_bb g1882(.a(n1879_1),.b(n1880_1),.q(_w_14769));
  bfr _b_6955(.a(_w_8857),.q(_w_8858));
  bfr _b_6959(.a(_w_8861),.q(_w_8862));
  bfr _b_9290(.a(_w_11192),.q(_w_11193));
  bfr _b_6960(.a(_w_8862),.q(_w_8863));
  bfr _b_6961(.a(_w_8863),.q(_w_8864));
  bfr _b_9516(.a(_w_11418),.q(_w_11419));
  bfr _b_7703(.a(_w_9605),.q(_w_9606));
  bfr _b_6962(.a(_w_8864),.q(_w_8865));
  bfr _b_13845(.a(_w_15747),.q(_w_15748));
  bfr _b_6967(.a(_w_8869),.q(_w_8870));
  bfr _b_6974(.a(_w_8876),.q(_w_8877));
  bfr _b_6975(.a(_w_8877),.q(_w_8878));
  bfr _b_6977(.a(_w_8879),.q(_w_8880));
  bfr _b_4518(.a(_w_6420),.q(_w_6421));
  bfr _b_6981(.a(_w_8883),.q(_w_8884));
  bfr _b_4519(.a(_w_6421),.q(_w_6422));
  bfr _b_8932(.a(_w_10834),.q(_w_10835));
  bfr _b_6983(.a(_w_8885),.q(_w_8886));
  bfr _b_6985(.a(_w_8887),.q(_w_8888));
  bfr _b_9542(.a(_w_11444),.q(_w_11445));
  bfr _b_6986(.a(_w_8888),.q(_w_8889));
  bfr _b_6987(.a(_w_8889),.q(_w_8890));
  bfr _b_6988(.a(_w_8890),.q(_w_8891));
  or_bb g1520(.a(n1518_0),.b(n1519),.q(n1520));
  bfr _b_4068(.a(_w_5970),.q(_w_5971));
  bfr _b_6989(.a(_w_8891),.q(_w_8892));
  bfr _b_5083(.a(_w_6985),.q(_w_6986));
  bfr _b_6993(.a(_w_8895),.q(_w_8896));
  bfr _b_6994(.a(_w_8896),.q(_w_8897));
  bfr _b_8630(.a(_w_10532),.q(_w_10533));
  bfr _b_11874(.a(_w_13776),.q(_w_13777));
  bfr _b_6997(.a(_w_8899),.q(_w_8900));
  bfr _b_12580(.a(_w_14482),.q(_w_14483));
  bfr _b_6998(.a(_w_8900),.q(_w_8901));
  bfr _b_5461(.a(_w_7363),.q(_w_7364));
  bfr _b_6999(.a(_w_8901),.q(_w_8902));
  bfr _b_12131(.a(_w_14033),.q(_w_14034));
  bfr _b_5458(.a(_w_7360),.q(_w_7361));
  bfr _b_7962(.a(_w_9864),.q(_w_9865));
  bfr _b_11583(.a(_w_13485),.q(_w_13486));
  bfr _b_9147(.a(_w_11049),.q(_w_11050));
  bfr _b_7000(.a(_w_8902),.q(_w_8903));
  bfr _b_4213(.a(_w_6115),.q(_w_6116));
  bfr _b_9384(.a(_w_11286),.q(_w_11287));
  bfr _b_7001(.a(_w_8903),.q(_w_8904));
  bfr _b_7002(.a(_w_8904),.q(_w_8905));
  bfr _b_7024(.a(_w_8926),.q(n803));
  bfr _b_3963(.a(_w_5865),.q(_w_5866));
  bfr _b_10027(.a(_w_11929),.q(_w_11930));
  bfr _b_9409(.a(_w_11311),.q(_w_11312));
  bfr _b_14058(.a(_w_15960),.q(_w_15961));
  bfr _b_9683(.a(_w_11585),.q(_w_11586));
  bfr _b_13078(.a(_w_14980),.q(n1236_1));
  bfr _b_7003(.a(_w_8905),.q(_w_8906));
  bfr _b_13505(.a(_w_15407),.q(_w_15408));
  bfr _b_7004(.a(_w_8906),.q(_w_8907));
  spl2 g787_s_0(.a(n787),.q0(n787_0),.q1(n787_1));
  bfr _b_8715(.a(_w_10617),.q(_w_10618));
  bfr _b_11937(.a(_w_13839),.q(_w_13840));
  bfr _b_9644(.a(_w_11546),.q(_w_11547));
  bfr _b_7005(.a(_w_8907),.q(_w_8908));
  bfr _b_8026(.a(_w_9928),.q(_w_9929));
  bfr _b_7009(.a(_w_8911),.q(_w_8912));
  bfr _b_8755(.a(_w_10657),.q(_w_10658));
  bfr _b_7013(.a(_w_8915),.q(_w_8916));
  bfr _b_7217(.a(_w_9119),.q(_w_9120));
  bfr _b_7015(.a(_w_8917),.q(_w_8918));
  or_bb g1722(.a(n1672_0),.b(n1721_0),.q(n1722));
  and_bi g1162(.a(n1149_1),.b(n1152_1),.q(n1162));
  bfr _b_7016(.a(_w_8918),.q(_w_8919));
  bfr _b_7945(.a(_w_9847),.q(_w_9848));
  and_bb g532(.a(N103_10),.b(N375_10),.q(_w_14524));
  bfr _b_7017(.a(_w_8919),.q(_w_8920));
  bfr _b_7019(.a(_w_8921),.q(_w_8922));
  bfr _b_11379(.a(_w_13281),.q(_w_13282));
  and_bb g1207(.a(n1180_1),.b(n1205_1),.q(_w_8369));
  bfr _b_7020(.a(_w_8922),.q(_w_8923));
  bfr _b_8583(.a(_w_10485),.q(_w_10486));
  bfr _b_7025(.a(_w_8927),.q(_w_8928));
  bfr _b_7028(.a(_w_8930),.q(_w_8931));
  bfr _b_7031(.a(_w_8933),.q(_w_8934));
  bfr _b_4605(.a(_w_6507),.q(_w_6508));
  bfr _b_7032(.a(_w_8934),.q(_w_8935));
  bfr _b_7033(.a(_w_8935),.q(_w_8936));
  bfr _b_8849(.a(_w_10751),.q(_w_10752));
  bfr _b_7034(.a(_w_8936),.q(_w_8937));
  bfr _b_7035(.a(_w_8937),.q(_w_8938));
  bfr _b_7036(.a(_w_8938),.q(n828));
  spl2 g1269_s_0(.a(n1269),.q0(n1269_0),.q1(n1269_1));
  bfr _b_7037(.a(_w_8939),.q(_w_8940));
  bfr _b_7038(.a(_w_8940),.q(_w_8941));
  bfr _b_12512(.a(_w_14414),.q(_w_14415));
  bfr _b_7039(.a(_w_8941),.q(_w_8942));
  or_bb g1130(.a(n1128_0),.b(n1129),.q(n1130));
  bfr _b_8499(.a(_w_10401),.q(_w_10402));
  bfr _b_9324(.a(_w_11226),.q(n151));
  bfr _b_7041(.a(_w_8943),.q(n797));
  bfr _b_4369(.a(_w_6271),.q(N120_7));
  bfr _b_7043(.a(_w_8945),.q(_w_8946));
  bfr _b_7045(.a(_w_8947),.q(n274_1));
  bfr _b_8137(.a(_w_10039),.q(_w_10040));
  bfr _b_7046(.a(_w_8948),.q(n794));
  bfr _b_7047(.a(_w_8949),.q(n470));
  bfr _b_12199(.a(_w_14101),.q(_w_14102));
  bfr _b_9378(.a(_w_11280),.q(_w_11281));
  bfr _b_7049(.a(_w_8951),.q(_w_8952));
  bfr _b_7050(.a(_w_8952),.q(_w_8953));
  spl2 g297_s_0(.a(n297),.q0(n297_0),.q1(n297_1));
  bfr _b_9618(.a(_w_11520),.q(_w_11521));
  bfr _b_7055(.a(_w_8957),.q(_w_8958));
  bfr _b_11198(.a(_w_13100),.q(n1812_1));
  bfr _b_7465(.a(_w_9367),.q(n1564_1));
  bfr _b_11644(.a(_w_13546),.q(_w_13547));
  bfr _b_8331(.a(_w_10233),.q(_w_10234));
  bfr _b_7056(.a(_w_8958),.q(_w_8959));
  bfr _b_7061(.a(_w_8963),.q(_w_8964));
  bfr _b_4916(.a(_w_6818),.q(_w_6819));
  and_bb g950(.a(N137_12),.b(N409_12),.q(n950));
  bfr _b_7062(.a(_w_8964),.q(_w_8965));
  bfr _b_13636(.a(N290),.q(_w_15538));
  bfr _b_7064(.a(_w_8966),.q(_w_8967));
  bfr _b_7066(.a(_w_8968),.q(_w_8969));
  bfr _b_7067(.a(_w_8969),.q(_w_8970));
  bfr _b_4616(.a(_w_6518),.q(_w_6519));
  bfr _b_7068(.a(_w_8970),.q(_w_8971));
  bfr _b_7072(.a(_w_8974),.q(_w_8975));
  bfr _b_7073(.a(_w_8975),.q(_w_8976));
  bfr _b_12413(.a(_w_14315),.q(_w_14316));
  bfr _b_9835(.a(_w_11737),.q(_w_11738));
  bfr _b_7075(.a(_w_8977),.q(_w_8978));
  bfr _b_7076(.a(_w_8978),.q(_w_8979));
  bfr _b_7078(.a(_w_8980),.q(_w_8981));
  bfr _b_7080(.a(_w_8982),.q(_w_8983));
  bfr _b_11312(.a(_w_13214),.q(_w_13215));
  bfr _b_4889(.a(_w_6791),.q(_w_6792));
  bfr _b_9754(.a(_w_11656),.q(_w_11657));
  bfr _b_8574(.a(_w_10476),.q(_w_10477));
  bfr _b_7085(.a(_w_8987),.q(_w_8988));
  bfr _b_8395(.a(_w_10297),.q(n188));
  bfr _b_7086(.a(_w_8988),.q(_w_8989));
  bfr _b_7087(.a(_w_8989),.q(_w_8990));
  bfr _b_7089(.a(_w_8991),.q(_w_8992));
  and_bi g1749(.a(n1747_0),.b(n1748),.q(n1749));
  bfr _b_7090(.a(_w_8992),.q(_w_8993));
  bfr _b_10442(.a(_w_12344),.q(_w_12345));
  bfr _b_7092(.a(_w_8994),.q(_w_8995));
  bfr _b_14348(.a(_w_16250),.q(_w_16251));
  bfr _b_14249(.a(_w_16151),.q(_w_16152));
  bfr _b_9540(.a(_w_11442),.q(_w_11443));
  or_bb g669(.a(n667_0),.b(n668),.q(n669));
  bfr _b_7093(.a(_w_8995),.q(_w_8996));
  bfr _b_12023(.a(_w_13925),.q(_w_13926));
  bfr _b_9268(.a(_w_11170),.q(_w_11171));
  bfr _b_12527(.a(_w_14429),.q(_w_14430));
  bfr _b_6704(.a(_w_8606),.q(_w_8607));
  bfr _b_7094(.a(_w_8996),.q(_w_8997));
  bfr _b_7096(.a(_w_8998),.q(_w_8999));
  bfr _b_5782(.a(_w_7684),.q(_w_7685));
  bfr _b_7098(.a(_w_9000),.q(_w_9001));
  bfr _b_13839(.a(_w_15741),.q(_w_15742));
  bfr _b_7104(.a(_w_9006),.q(_w_9007));
  and_bi g1425(.a(n1424_0),.b(n1371_0),.q(n1425));
  bfr _b_7105(.a(_w_9007),.q(_w_9008));
  spl2 g1139_s_0(.a(n1139),.q0(n1139_0),.q1(n1139_1));
  bfr _b_7108(.a(_w_9010),.q(_w_9011));
  bfr _b_7113(.a(_w_9015),.q(_w_9016));
  bfr _b_7114(.a(_w_9016),.q(_w_9017));
  bfr _b_7552(.a(_w_9454),.q(_w_9455));
  bfr _b_7118(.a(_w_9020),.q(_w_9021));
  bfr _b_7119(.a(_w_9021),.q(_w_9022));
  bfr _b_7121(.a(_w_9023),.q(_w_9024));
  bfr _b_7122(.a(_w_9024),.q(_w_9025));
  bfr _b_7124(.a(_w_9026),.q(_w_9027));
  bfr _b_7129(.a(_w_9031),.q(_w_9032));
  bfr _b_7130(.a(_w_9032),.q(_w_9033));
  bfr _b_7131(.a(_w_9033),.q(_w_9034));
  bfr _b_8233(.a(_w_10135),.q(_w_10136));
  bfr _b_11316(.a(_w_13218),.q(_w_13219));
  bfr _b_7132(.a(_w_9034),.q(_w_9035));
  spl4L N188_s_1(.a(N188_0),.q0(N188_4),.q1(N188_5),.q2(_w_7952),.q3(_w_7954));
  bfr _b_4252(.a(_w_6154),.q(_w_6155));
  bfr _b_7133(.a(_w_9035),.q(_w_9036));
  bfr _b_11416(.a(_w_13318),.q(_w_13319));
  bfr _b_9813(.a(_w_11715),.q(_w_11716));
  bfr _b_6677(.a(_w_8579),.q(_w_8580));
  bfr _b_7297(.a(_w_9199),.q(_w_9200));
  bfr _b_7135(.a(_w_9037),.q(_w_9038));
  bfr _b_11012(.a(_w_12914),.q(_w_12915));
  bfr _b_7142(.a(_w_9044),.q(_w_9045));
  bfr _b_7147(.a(_w_9049),.q(_w_9050));
  bfr _b_12124(.a(_w_14026),.q(_w_14027));
  bfr _b_7148(.a(_w_9050),.q(_w_9051));
  bfr _b_12690(.a(_w_14592),.q(_w_14593));
  bfr _b_7149(.a(_w_9051),.q(_w_9052));
  bfr _b_7151(.a(_w_9053),.q(_w_9054));
  and_bb g822(.a(N18_18),.b(N511_5),.q(_w_11158));
  bfr _b_7153(.a(_w_9055),.q(_w_9056));
  bfr _b_7154(.a(_w_9056),.q(_w_9057));
  bfr _b_7155(.a(_w_9057),.q(_w_9058));
  bfr _b_9240(.a(_w_11142),.q(_w_11143));
  bfr _b_7157(.a(_w_9059),.q(_w_9060));
  bfr _b_6859(.a(_w_8761),.q(_w_8762));
  bfr _b_8223(.a(_w_10125),.q(_w_10126));
  and_bb g1072(.a(N222_16),.b(N341_17),.q(n1072));
  bfr _b_7161(.a(_w_9063),.q(_w_9064));
  bfr _b_7756(.a(_w_9658),.q(n1600_1));
  bfr _b_7162(.a(_w_9064),.q(_w_9065));
  bfr _b_7165(.a(_w_9067),.q(_w_9068));
  bfr _b_9210(.a(_w_11112),.q(_w_11113));
  bfr _b_7166(.a(_w_9068),.q(_w_9069));
  bfr _b_7173(.a(_w_9075),.q(_w_9076));
  bfr _b_12716(.a(_w_14618),.q(_w_14619));
  bfr _b_7175(.a(_w_9077),.q(_w_9078));
  bfr _b_5097(.a(_w_6999),.q(_w_7000));
  bfr _b_7176(.a(_w_9078),.q(_w_9079));
  bfr _b_7183(.a(_w_9085),.q(_w_9086));
  bfr _b_5793(.a(_w_7695),.q(_w_7696));
  bfr _b_9019(.a(_w_10921),.q(_w_10922));
  and_bb g1054(.a(N494_8),.b(N69_17),.q(_w_8373));
  bfr _b_10203(.a(_w_12105),.q(_w_12106));
  bfr _b_9445(.a(_w_11347),.q(_w_11348));
  bfr _b_7187(.a(_w_9089),.q(_w_9090));
  bfr _b_7188(.a(_w_9090),.q(_w_9091));
  bfr _b_7190(.a(_w_9092),.q(_w_9093));
  bfr _b_12910(.a(_w_14812),.q(_w_14813));
  bfr _b_5350(.a(_w_7252),.q(_w_7253));
  bfr _b_8150(.a(_w_10052),.q(_w_10053));
  bfr _b_7191(.a(_w_9093),.q(_w_9094));
  bfr _b_7192(.a(_w_9094),.q(_w_9095));
  bfr _b_7194(.a(_w_9096),.q(_w_9097));
  bfr _b_7195(.a(_w_9097),.q(_w_9098));
  bfr _b_7196(.a(_w_9098),.q(_w_9099));
  and_bb g203(.a(n189_1),.b(n201_1),.q(_w_11629));
  bfr _b_7198(.a(_w_9100),.q(_w_9101));
  bfr _b_7200(.a(_w_9102),.q(_w_9103));
  bfr _b_7201(.a(_w_9103),.q(_w_9104));
  bfr _b_7210(.a(_w_9112),.q(_w_9113));
  bfr _b_7211(.a(_w_9113),.q(_w_9114));
  bfr _b_7212(.a(_w_9114),.q(_w_9115));
  bfr _b_8997(.a(_w_10899),.q(_w_10900));
  bfr _b_7215(.a(_w_9117),.q(_w_9118));
  bfr _b_12667(.a(_w_14569),.q(n467));
  bfr _b_7216(.a(_w_9118),.q(_w_9119));
  spl2 g1257_s_0(.a(n1257),.q0(n1257_0),.q1(n1257_1));
  bfr _b_6909(.a(_w_8811),.q(_w_8812));
  bfr _b_9608(.a(_w_11510),.q(_w_11511));
  bfr _b_7222(.a(_w_9124),.q(_w_9125));
  bfr _b_7474(.a(_w_9376),.q(_w_9377));
  bfr _b_7223(.a(_w_9125),.q(_w_9126));
  bfr _b_7224(.a(_w_9126),.q(_w_9127));
  bfr _b_13735(.a(_w_15637),.q(_w_15638));
  bfr _b_7225(.a(_w_9127),.q(_w_9128));
  and_bi g1452(.a(n1446_1),.b(n1449_1),.q(n1452));
  bfr _b_9090(.a(_w_10992),.q(_w_10993));
  bfr _b_7226(.a(_w_9128),.q(N188_3));
  bfr _b_7229(.a(_w_9131),.q(n770));
  bfr _b_7230(.a(_w_9132),.q(n1023));
  spl2 g1067_s_0(.a(n1067),.q0(n1067_0),.q1(n1067_1));
  bfr _b_7231(.a(_w_9133),.q(n1258));
  spl2 g408_s_0(.a(n408),.q0(n408_0),.q1(n408_1));
  bfr _b_7233(.a(_w_9135),.q(n764));
  bfr _b_13152(.a(_w_15054),.q(_w_15055));
  spl2 g1793_s_0(.a(n1793),.q0(n1793_0),.q1(n1793_1));
  bfr _b_7234(.a(_w_9136),.q(n758));
  bfr _b_7235(.a(_w_9137),.q(n755));
  bfr _b_7236(.a(_w_9138),.q(n752));
  bfr _b_7238(.a(_w_9140),.q(n743));
  bfr _b_8957(.a(_w_10859),.q(n1020));
  bfr _b_7239(.a(_w_9141),.q(_w_9142));
  bfr _b_7240(.a(_w_9142),.q(_w_9143));
  bfr _b_13481(.a(_w_15383),.q(_w_15384));
  bfr _b_3433(.a(_w_5335),.q(_w_5336));
  bfr _b_7241(.a(_w_9143),.q(_w_9144));
  spl2 g1086_s_0(.a(n1086),.q0(n1086_0),.q1(n1086_1));
  bfr _b_9157(.a(_w_11059),.q(n612));
  spl4L N460_s_2(.a(N460_1),.q0(N460_8),.q1(N460_9),.q2(N460_10),.q3(N460_11));
  bfr _b_7242(.a(_w_9144),.q(_w_9145));
  bfr _b_13826(.a(_w_15728),.q(_w_15729));
  bfr _b_10301(.a(_w_12203),.q(_w_12204));
  bfr _b_7243(.a(_w_9145),.q(_w_9146));
  bfr _b_9161(.a(_w_11063),.q(_w_11064));
  bfr _b_7244(.a(_w_9146),.q(_w_9147));
  bfr _b_7251(.a(_w_9153),.q(_w_9154));
  bfr _b_14118(.a(_w_16020),.q(_w_16021));
  bfr _b_13066(.a(_w_14968),.q(n1568));
  bfr _b_12026(.a(_w_13928),.q(_w_13929));
  bfr _b_7254(.a(_w_9156),.q(_w_9157));
  spl2 g863_s_0(.a(n863),.q0(n863_0),.q1(_w_6276));
  bfr _b_3580(.a(_w_5482),.q(_w_5483));
  bfr _b_8126(.a(_w_10028),.q(_w_10029));
  bfr _b_7260(.a(_w_9162),.q(n1032));
  bfr _b_7262(.a(_w_9164),.q(_w_9165));
  and_bb g142(.a(N324_7),.b(N52_7),.q(_w_9687));
  spl2 g994_s_0(.a(n994),.q0(n994_0),.q1(n994_1));
  bfr _b_7263(.a(_w_9165),.q(_w_9166));
  bfr _b_12838(.a(_w_14740),.q(_w_14741));
  bfr _b_9565(.a(_w_11467),.q(_w_11468));
  spl2 g1161_s_0(.a(n1161),.q0(n1161_0),.q1(n1161_1));
  bfr _b_7264(.a(_w_9166),.q(_w_9167));
  bfr _b_12448(.a(_w_14350),.q(_w_14351));
  bfr _b_7266(.a(_w_9168),.q(_w_9169));
  bfr _b_13352(.a(_w_15254),.q(_w_15255));
  bfr _b_7267(.a(_w_9169),.q(_w_9170));
  bfr _b_7940(.a(_w_9842),.q(_w_9843));
  bfr _b_7273(.a(_w_9175),.q(_w_9176));
  bfr _b_6996(.a(_w_8898),.q(_w_8899));
  bfr _b_7276(.a(_w_9178),.q(_w_9179));
  bfr _b_7755(.a(_w_9657),.q(_w_9658));
  bfr _b_4932(.a(_w_6834),.q(_w_6835));
  bfr _b_7278(.a(_w_9180),.q(_w_9181));
  bfr _b_10752(.a(_w_12654),.q(_w_12655));
  bfr _b_8740(.a(_w_10642),.q(_w_10643));
  bfr _b_9165(.a(_w_11067),.q(n1751));
  bfr _b_7279(.a(_w_9181),.q(_w_9182));
  bfr _b_10001(.a(_w_11903),.q(_w_11904));
  bfr _b_11413(.a(_w_13315),.q(_w_13316));
  bfr _b_7280(.a(_w_9182),.q(_w_9183));
  bfr _b_7649(.a(_w_9551),.q(_w_9552));
  bfr _b_7286(.a(_w_9188),.q(_w_9189));
  bfr _b_13272(.a(_w_15174),.q(_w_15175));
  bfr _b_6242(.a(_w_8144),.q(_w_8145));
  bfr _b_7288(.a(_w_9190),.q(_w_9191));
  bfr _b_7289(.a(_w_9191),.q(_w_9192));
  bfr _b_12375(.a(_w_14277),.q(_w_14278));
  bfr _b_10742(.a(_w_12644),.q(_w_12645));
  bfr _b_7291(.a(_w_9193),.q(_w_9194));
  bfr _b_14339(.a(_w_16241),.q(_w_16242));
  bfr _b_7293(.a(_w_9195),.q(_w_9196));
  bfr _b_9359(.a(_w_11261),.q(_w_11262));
  bfr _b_7102(.a(_w_9004),.q(_w_9005));
  bfr _b_7295(.a(_w_9197),.q(_w_9198));
  bfr _b_13080(.a(_w_14982),.q(_w_14983));
  bfr _b_7300(.a(_w_9202),.q(n641));
  bfr _b_12127(.a(_w_14029),.q(_w_14030));
  bfr _b_7301(.a(_w_9203),.q(n1129));
  bfr _b_7721(.a(_w_9623),.q(_w_9624));
  spl2 g1465_s_0(.a(n1465),.q0(n1465_0),.q1(n1465_1));
  bfr _b_6474(.a(_w_8376),.q(_w_8377));
  bfr _b_7302(.a(_w_9204),.q(_w_9205));
  bfr _b_12126(.a(_w_14028),.q(_w_14029));
  bfr _b_9520(.a(_w_11422),.q(_w_11423));
  bfr _b_12612(.a(_w_14514),.q(_w_14515));
  bfr _b_7303(.a(_w_9205),.q(_w_9206));
  bfr _b_12325(.a(_w_14227),.q(_w_14228));
  bfr _b_8922(.a(_w_10824),.q(_w_10825));
  bfr _b_7306(.a(_w_9208),.q(n969));
  bfr _b_9985(.a(_w_11887),.q(_w_11888));
  bfr _b_7307(.a(_w_9209),.q(n1804));
  bfr _b_8008(.a(_w_9910),.q(_w_9911));
  bfr _b_7312(.a(_w_9214),.q(_w_9215));
  bfr _b_7313(.a(_w_9215),.q(_w_9216));
  bfr _b_7134(.a(_w_9036),.q(_w_9037));
  bfr _b_9860(.a(_w_11762),.q(_w_11763));
  bfr _b_4669(.a(_w_6571),.q(_w_6572));
  bfr _b_7322(.a(_w_9224),.q(_w_9225));
  bfr _b_6791(.a(_w_8693),.q(_w_8694));
  bfr _b_7923(.a(_w_9825),.q(_w_9826));
  bfr _b_7327(.a(_w_9229),.q(_w_9230));
  bfr _b_7328(.a(_w_9230),.q(_w_9231));
  or_bb g174(.a(n137_0),.b(n173_0),.q(n174));
  bfr _b_7329(.a(_w_9231),.q(_w_9232));
  bfr _b_7331(.a(_w_9233),.q(_w_9234));
  bfr _b_7332(.a(_w_9234),.q(_w_9235));
  bfr _b_7333(.a(_w_9235),.q(_w_9236));
  bfr _b_7334(.a(_w_9236),.q(_w_9237));
  bfr _b_10206(.a(_w_12108),.q(_w_12109));
  bfr _b_7338(.a(_w_9240),.q(_w_9241));
  bfr _b_9464(.a(_w_11366),.q(_w_11367));
  bfr _b_7343(.a(_w_9245),.q(n773));
  and_bi g1761(.a(n1759_0),.b(n1760),.q(n1761));
  bfr _b_7345(.a(_w_9247),.q(n662));
  bfr _b_7347(.a(_w_9249),.q(n1138));
  bfr _b_5625(.a(_w_7527),.q(_w_7528));
  bfr _b_9757(.a(_w_11659),.q(_w_11660));
  bfr _b_7350(.a(_w_9252),.q(n1328));
  bfr _b_6476(.a(_w_8378),.q(_w_8379));
  spl2 g848_s_0(.a(n848),.q0(n848_0),.q1(n848_1));
  bfr _b_8847(.a(_w_10749),.q(_w_10750));
  bfr _b_12815(.a(_w_14717),.q(_w_14718));
  bfr _b_7357(.a(_w_9259),.q(_w_9260));
  bfr _b_9928(.a(_w_11830),.q(_w_11831));
  bfr _b_4995(.a(_w_6897),.q(_w_6898));
  bfr _b_7361(.a(_w_9263),.q(_w_9264));
  bfr _b_7365(.a(_w_9267),.q(_w_9268));
  bfr _b_4140(.a(_w_6042),.q(_w_6043));
  bfr _b_7367(.a(_w_9269),.q(_w_9270));
  bfr _b_7368(.a(_w_9270),.q(_w_9271));
  bfr _b_7372(.a(_w_9274),.q(_w_9275));
  bfr _b_11552(.a(_w_13454),.q(_w_13455));
  bfr _b_7373(.a(_w_9275),.q(_w_9276));
  or_bb g681(.a(n679_0),.b(n680),.q(n681));
  bfr _b_7376(.a(_w_9278),.q(_w_9279));
  bfr _b_7379(.a(_w_9281),.q(_w_9282));
  spl2 g46_s_0(.a(n46),.q0(n46_0),.q1(_w_13850));
  bfr _b_7381(.a(_w_9283),.q(_w_9284));
  bfr _b_7382(.a(_w_9284),.q(_w_9285));
  bfr _b_7386(.a(_w_9288),.q(_w_9289));
  bfr _b_7388(.a(_w_9290),.q(n650));
  bfr _b_7591(.a(_w_9493),.q(_w_9494));
  spl2 g696_s_0(.a(n696),.q0(n696_0),.q1(n696_1));
  bfr _b_7389(.a(_w_9291),.q(n701));
  bfr _b_13651(.a(_w_15553),.q(_w_15554));
  bfr _b_7392(.a(_w_9294),.q(_w_9295));
  bfr _b_7393(.a(_w_9295),.q(_w_9296));
  bfr _b_8648(.a(_w_10550),.q(_w_10551));
  and_bi g1707(.a(n1706_0),.b(n1677_0),.q(n1707));
  bfr _b_7395(.a(_w_9297),.q(_w_9298));
  bfr _b_6766(.a(_w_8668),.q(_w_8669));
  bfr _b_7396(.a(_w_9298),.q(_w_9299));
  bfr _b_7397(.a(_w_9299),.q(_w_9300));
  bfr _b_7401(.a(_w_9303),.q(_w_9304));
  spl4L N511_s_1(.a(N511_0),.q0(N511_4),.q1(N511_5),.q2(N511_6),.q3(N511_7));
  spl2 g1890_s_0(.a(n1890),.q0(n1890_0),.q1(n1890_1));
  bfr _b_7402(.a(_w_9304),.q(_w_9305));
  spl2 g840_s_0(.a(n840),.q0(n840_0),.q1(n840_1));
  bfr _b_5469(.a(_w_7371),.q(_w_7372));
  bfr _b_7404(.a(_w_9306),.q(_w_9307));
  bfr _b_14100(.a(_w_16002),.q(_w_16003));
  bfr _b_12328(.a(_w_14230),.q(_w_14231));
  bfr _b_9121(.a(_w_11023),.q(n1017));
  bfr _b_7408(.a(_w_9310),.q(_w_9311));
  bfr _b_7409(.a(_w_9311),.q(_w_9312));
  bfr _b_7411(.a(_w_9313),.q(n1601));
  bfr _b_11815(.a(_w_13717),.q(_w_13718));
  bfr _b_7414(.a(_w_9316),.q(_w_9317));
  bfr _b_7415(.a(_w_9317),.q(_w_9318));
  bfr _b_10262(.a(_w_12164),.q(_w_12165));
  bfr _b_7417(.a(_w_9319),.q(_w_9320));
  bfr _b_7420(.a(_w_9322),.q(_w_9323));
  bfr _b_7526(.a(_w_9428),.q(_w_9429));
  bfr _b_7575(.a(_w_9477),.q(_w_9478));
  bfr _b_9877(.a(_w_11779),.q(_w_11780));
  bfr _b_7421(.a(_w_9323),.q(_w_9324));
  bfr _b_8696(.a(_w_10598),.q(_w_10599));
  bfr _b_7425(.a(_w_9327),.q(_w_9328));
  bfr _b_14032(.a(_w_15934),.q(_w_15935));
  bfr _b_13384(.a(_w_15286),.q(_w_15287));
  bfr _b_7426(.a(_w_9328),.q(_w_9329));
  bfr _b_7893(.a(_w_9795),.q(_w_9796));
  bfr _b_8238(.a(_w_10140),.q(_w_10141));
  bfr _b_6164(.a(_w_8066),.q(_w_8067));
  bfr _b_7432(.a(_w_9334),.q(_w_9335));
  bfr _b_10823(.a(_w_12725),.q(_w_12726));
  bfr _b_7433(.a(_w_9335),.q(_w_9336));
  bfr _b_8195(.a(_w_10097),.q(_w_10098));
  bfr _b_13515(.a(_w_15417),.q(_w_15418));
  bfr _b_13237(.a(_w_15139),.q(_w_15140));
  or_bb g1629(.a(n1619_0),.b(n1628_0),.q(n1629));
  bfr _b_7980(.a(_w_9882),.q(N3552));
  bfr _b_7434(.a(_w_9336),.q(_w_9337));
  bfr _b_7436(.a(_w_9338),.q(n1447));
  and_bi g216(.a(n214_0),.b(n215),.q(n216));
  bfr _b_7437(.a(_w_9339),.q(_w_9340));
  bfr _b_9020(.a(_w_10922),.q(_w_10923));
  bfr _b_7441(.a(_w_9343),.q(_w_9344));
  bfr _b_7443(.a(_w_9345),.q(_w_9346));
  bfr _b_7446(.a(_w_9348),.q(_w_9349));
  bfr _b_10078(.a(_w_11980),.q(_w_11981));
  bfr _b_7450(.a(_w_9352),.q(_w_9353));
  bfr _b_7451(.a(_w_9353),.q(_w_9354));
  bfr _b_9433(.a(_w_11335),.q(_w_11336));
  or_bb g1446(.a(n1364_0),.b(n1445_0),.q(n1446));
  spl4L N341_s_3(.a(N341_2),.q0(N341_12),.q1(N341_13),.q2(N341_14),.q3(N341_15));
  and_bi g1295(.a(n1288_1),.b(n1293_1),.q(_w_13430));
  bfr _b_7453(.a(_w_9355),.q(_w_9356));
  bfr _b_7454(.a(_w_9356),.q(_w_9357));
  bfr _b_7457(.a(_w_9359),.q(_w_9360));
  bfr _b_7459(.a(_w_9361),.q(_w_9362));
  bfr _b_7460(.a(_w_9362),.q(n626));
  and_bb g870(.a(n841_1),.b(n868_1),.q(_w_11606));
  bfr _b_10100(.a(_w_12002),.q(_w_12003));
  or_bb g1521(.a(n1455_0),.b(n1520_0),.q(n1521));
  bfr _b_7461(.a(_w_9363),.q(n858));
  bfr _b_7463(.a(_w_9365),.q(_w_9366));
  bfr _b_13690(.a(_w_15592),.q(_w_15593));
  bfr _b_8203(.a(_w_10105),.q(_w_10106));
  bfr _b_6505(.a(_w_8407),.q(_w_8408));
  bfr _b_9316(.a(_w_11218),.q(_w_11219));
  bfr _b_13749(.a(_w_15651),.q(_w_15652));
  bfr _b_3984(.a(_w_5886),.q(_w_5887));
  spl2 g374_s_0(.a(n374),.q0(n374_0),.q1(n374_1));
  bfr _b_7469(.a(_w_9371),.q(n1060));
  bfr _b_12280(.a(_w_14182),.q(_w_14183));
  and_bi g1364(.a(n1351_1),.b(n1354_1),.q(n1364));
  bfr _b_7696(.a(_w_9598),.q(_w_9599));
  or_bb g380(.a(n307_1),.b(n379_0),.q(_w_12026));
  bfr _b_7470(.a(_w_9372),.q(n746));
  bfr _b_11532(.a(_w_13434),.q(n1352));
  bfr _b_7473(.a(_w_9375),.q(_w_9376));
  spl2 g774_s_0(.a(n774),.q0(n774_0),.q1(n774_1));
  bfr _b_7475(.a(_w_9377),.q(_w_9378));
  bfr _b_7476(.a(_w_9378),.q(_w_9379));
  bfr _b_11714(.a(_w_13616),.q(_w_13617));
  bfr _b_7484(.a(_w_9386),.q(_w_9387));
  bfr _b_5025(.a(_w_6927),.q(_w_6928));
  bfr _b_8146(.a(_w_10048),.q(_w_10049));
  bfr _b_7487(.a(_w_9389),.q(_w_9390));
  bfr _b_7490(.a(_w_9392),.q(_w_9393));
  bfr _b_10463(.a(_w_12365),.q(_w_12366));
  bfr _b_7491(.a(_w_9393),.q(_w_9394));
  spl2 g1597_s_0(.a(n1597),.q0(n1597_0),.q1(n1597_1));
  bfr _b_7492(.a(_w_9394),.q(_w_9395));
  bfr _b_11747(.a(_w_13649),.q(_w_13650));
  bfr _b_8250(.a(_w_10152),.q(_w_10153));
  bfr _b_7493(.a(_w_9395),.q(_w_9396));
  bfr _b_7494(.a(_w_9396),.q(N120_1));
  bfr _b_12116(.a(_w_14018),.q(_w_14019));
  and_bi g1585(.a(n1584_0),.b(n1539_0),.q(n1585));
  bfr _b_7495(.a(_w_9397),.q(_w_9398));
  bfr _b_12359(.a(_w_14261),.q(_w_14262));
  bfr _b_7496(.a(_w_9398),.q(_w_9399));
  bfr _b_7497(.a(_w_9399),.q(_w_9400));
  bfr _b_7499(.a(_w_9401),.q(_w_9402));
  bfr _b_7504(.a(_w_9406),.q(_w_9407));
  bfr _b_7507(.a(_w_9409),.q(_w_9410));
  and_bi g1708(.a(n1677_1),.b(n1706_1),.q(_w_8384));
  bfr _b_7512(.a(_w_9414),.q(_w_9415));
  bfr _b_7517(.a(_w_9419),.q(_w_9420));
  bfr _b_3824(.a(_w_5726),.q(_w_5727));
  bfr _b_7881(.a(_w_9783),.q(_w_9784));
  bfr _b_7518(.a(_w_9420),.q(_w_9421));
  bfr _b_11158(.a(_w_13060),.q(_w_13061));
  spl2 g161_s_0(.a(n161),.q0(n161_0),.q1(n161_1));
  bfr _b_7519(.a(_w_9421),.q(_w_9422));
  bfr _b_7523(.a(_w_9425),.q(_w_9426));
  bfr _b_7527(.a(_w_9429),.q(_w_9430));
  bfr _b_7529(.a(_w_9431),.q(_w_9432));
  bfr _b_9967(.a(_w_11869),.q(_w_11870));
  bfr _b_9462(.a(_w_11364),.q(_w_11365));
  bfr _b_7530(.a(_w_9432),.q(_w_9433));
  bfr _b_11325(.a(_w_13227),.q(_w_13228));
  spl2 g1494_s_0(.a(n1494),.q0(n1494_0),.q1(n1494_1));
  bfr _b_7531(.a(_w_9433),.q(_w_9434));
  bfr _b_7538(.a(_w_9440),.q(_w_9441));
  bfr _b_4878(.a(_w_6780),.q(_w_6781));
  bfr _b_6672(.a(_w_8574),.q(_w_8575));
  bfr _b_9881(.a(_w_11783),.q(_w_11784));
  bfr _b_10260(.a(_w_12162),.q(_w_12163));
  or_bb g1771(.a(n1729_0),.b(n1770_0),.q(n1771));
  bfr _b_7539(.a(_w_9441),.q(_w_9442));
  bfr _b_8808(.a(_w_10710),.q(_w_10711));
  bfr _b_7910(.a(_w_9812),.q(_w_9813));
  bfr _b_8627(.a(_w_10529),.q(_w_10530));
  bfr _b_7542(.a(_w_9444),.q(_w_9445));
  bfr _b_12059(.a(_w_13961),.q(_w_13962));
  bfr _b_7543(.a(_w_9445),.q(_w_9446));
  bfr _b_13578(.a(_w_15480),.q(_w_15481));
  bfr _b_7544(.a(_w_9446),.q(_w_9447));
  bfr _b_14224(.a(_w_16126),.q(_w_16127));
  bfr _b_7545(.a(_w_9447),.q(_w_9448));
  bfr _b_7546(.a(_w_9448),.q(_w_9449));
  bfr _b_7548(.a(_w_9450),.q(_w_9451));
  bfr _b_7549(.a(_w_9451),.q(_w_9452));
  bfr _b_9229(.a(_w_11131),.q(_w_11132));
  bfr _b_8786(.a(_w_10688),.q(_w_10689));
  bfr _b_7550(.a(_w_9452),.q(N120_2));
  bfr _b_12765(.a(_w_14667),.q(_w_14668));
  spl4L N154_s_3(.a(N154_2),.q0(N154_12),.q1(_w_6430),.q2(_w_6438),.q3(_w_6450));
  bfr _b_7554(.a(_w_9456),.q(_w_9457));
  bfr _b_7555(.a(_w_9457),.q(_w_9458));
  bfr _b_7559(.a(_w_9461),.q(_w_9462));
  bfr _b_8804(.a(_w_10706),.q(_w_10707));
  bfr _b_7561(.a(_w_9463),.q(_w_9464));
  bfr _b_7563(.a(_w_9465),.q(_w_9466));
  bfr _b_7565(.a(_w_9467),.q(_w_9468));
  bfr _b_14074(.a(_w_15976),.q(_w_15977));
  bfr _b_12414(.a(_w_14316),.q(_w_14317));
  bfr _b_7296(.a(_w_9198),.q(_w_9199));
  bfr _b_7567(.a(_w_9469),.q(_w_9470));
  bfr _b_8158(.a(_w_10060),.q(_w_10061));
  bfr _b_11350(.a(_w_13252),.q(_w_13253));
  bfr _b_7569(.a(_w_9471),.q(_w_9472));
  bfr _b_7572(.a(_w_9474),.q(_w_9475));
  bfr _b_7574(.a(_w_9476),.q(_w_9477));
  bfr _b_7576(.a(_w_9478),.q(_w_9479));
  bfr _b_3814(.a(_w_5716),.q(_w_5717));
  bfr _b_7577(.a(_w_9479),.q(_w_9480));
  bfr _b_7878(.a(_w_9780),.q(_w_9781));
  bfr _b_6543(.a(_w_8445),.q(_w_8446));
  bfr _b_7580(.a(_w_9482),.q(_w_9483));
  bfr _b_7581(.a(_w_9483),.q(_w_9484));
  bfr _b_7584(.a(_w_9486),.q(_w_9487));
  bfr _b_7585(.a(_w_9487),.q(_w_9488));
  bfr _b_7586(.a(_w_9488),.q(_w_9489));
  bfr _b_7587(.a(_w_9489),.q(_w_9490));
  bfr _b_9797(.a(_w_11699),.q(_w_11700));
  bfr _b_12330(.a(_w_14232),.q(_w_14233));
  bfr _b_6934(.a(_w_8836),.q(_w_8837));
  bfr _b_7595(.a(_w_9497),.q(_w_9498));
  bfr _b_9454(.a(_w_11356),.q(_w_11357));
  bfr _b_7599(.a(_w_9501),.q(_w_9502));
  spl2 g1829_s_0(.a(n1829),.q0(n1829_0),.q1(n1829_1));
  bfr _b_7600(.a(_w_9502),.q(_w_9503));
  bfr _b_11002(.a(_w_12904),.q(_w_12905));
  bfr _b_7607(.a(_w_9509),.q(_w_9510));
  bfr _b_4106(.a(_w_6008),.q(_w_6009));
  bfr _b_7609(.a(_w_9511),.q(_w_9512));
  bfr _b_7625(.a(_w_9527),.q(_w_9528));
  spl2 g1620_s_0(.a(n1620),.q0(n1620_0),.q1(n1620_1));
  bfr _b_7611(.a(_w_9513),.q(_w_9514));
  spl2 g1695_s_0(.a(n1695),.q0(n1695_0),.q1(n1695_1));
  bfr _b_7613(.a(_w_9515),.q(_w_9516));
  bfr _b_7614(.a(_w_9516),.q(_w_9517));
  bfr _b_7615(.a(_w_9517),.q(_w_9518));
  bfr _b_8077(.a(_w_9979),.q(_w_9980));
  bfr _b_7616(.a(_w_9518),.q(_w_9519));
  bfr _b_11929(.a(_w_13831),.q(_w_13832));
  bfr _b_9475(.a(_w_11377),.q(_w_11378));
  bfr _b_7618(.a(_w_9520),.q(_w_9521));
  bfr _b_7619(.a(_w_9521),.q(_w_9522));
  bfr _b_9973(.a(_w_11875),.q(_w_11876));
  bfr _b_7621(.a(_w_9523),.q(_w_9524));
  bfr _b_6788(.a(_w_8690),.q(_w_8691));
  bfr _b_7622(.a(_w_9524),.q(_w_9525));
  bfr _b_7624(.a(_w_9526),.q(_w_9527));
  bfr _b_8182(.a(_w_10084),.q(_w_10085));
  spl2 g591_s_0(.a(n591),.q0(n591_0),.q1(n591_1));
  bfr _b_7629(.a(_w_9531),.q(_w_9532));
  and_bi g852(.a(n849),.b(n851),.q(n852));
  bfr _b_9233(.a(_w_11135),.q(_w_11136));
  bfr _b_7630(.a(_w_9532),.q(_w_9533));
  bfr _b_7633(.a(_w_9535),.q(_w_9536));
  bfr _b_13499(.a(_w_15401),.q(_w_15402));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(n235_1));
  bfr _b_7634(.a(_w_9536),.q(_w_9537));
  and_bi g271(.a(n270_0),.b(n238_0),.q(n271));
  bfr _b_8885(.a(_w_10787),.q(_w_10788));
  bfr _b_10644(.a(_w_12546),.q(_w_12547));
  bfr _b_7636(.a(_w_9538),.q(_w_9539));
  bfr _b_7637(.a(_w_9539),.q(_w_9540));
  bfr _b_7639(.a(_w_9541),.q(_w_9542));
  bfr _b_14376(.a(_w_16278),.q(_w_16279));
  bfr _b_7640(.a(_w_9542),.q(_w_9543));
  bfr _b_7643(.a(_w_9545),.q(_w_9546));
  bfr _b_7644(.a(_w_9546),.q(_w_9547));
  bfr _b_11524(.a(_w_13426),.q(_w_13427));
  bfr _b_8419(.a(_w_10321),.q(_w_10322));
  bfr _b_7645(.a(_w_9547),.q(n1075));
  bfr _b_7646(.a(_w_9548),.q(n767));
  bfr _b_9155(.a(_w_11057),.q(_w_11058));
  bfr _b_7647(.a(_w_9549),.q(_w_9550));
  bfr _b_7653(.a(_w_9555),.q(_w_9556));
  bfr _b_7654(.a(_w_9556),.q(_w_9557));
  bfr _b_12062(.a(_w_13964),.q(_w_13965));
  bfr _b_7656(.a(_w_9558),.q(_w_9559));
  bfr _b_8672(.a(_w_10574),.q(_w_10575));
  bfr _b_7658(.a(_w_9560),.q(n616));
  bfr _b_10086(.a(_w_11988),.q(_w_11989));
  bfr _b_7660(.a(_w_9562),.q(_w_9563));
  bfr _b_7775(.a(_w_9677),.q(_w_9678));
  bfr _b_4671(.a(_w_6573),.q(_w_6574));
  bfr _b_8332(.a(_w_10234),.q(_w_10235));
  bfr _b_8470(.a(_w_10372),.q(_w_10373));
  bfr _b_7919(.a(_w_9821),.q(_w_9822));
  bfr _b_7663(.a(_w_9565),.q(n1291_1));
  bfr _b_10364(.a(_w_12266),.q(_w_12267));
  bfr _b_5587(.a(_w_7489),.q(_w_7490));
  bfr _b_7668(.a(_w_9570),.q(_w_9571));
  bfr _b_10547(.a(_w_12449),.q(_w_12450));
  or_bb g225(.a(n223_0),.b(n224),.q(n225));
  bfr _b_7669(.a(_w_9571),.q(_w_9572));
  bfr _b_9842(.a(_w_11744),.q(_w_11745));
  bfr _b_12514(.a(_w_14416),.q(_w_14417));
  bfr _b_7671(.a(_w_9573),.q(n376));
  bfr _b_7674(.a(_w_9576),.q(_w_9577));
  bfr _b_11258(.a(_w_13160),.q(_w_13161));
  bfr _b_7676(.a(_w_9578),.q(_w_9579));
  bfr _b_4195(.a(_w_6097),.q(_w_6098));
  bfr _b_5831(.a(_w_7733),.q(_w_7734));
  bfr _b_9386(.a(_w_11288),.q(_w_11289));
  bfr _b_7246(.a(_w_9148),.q(_w_9149));
  bfr _b_8231(.a(_w_10133),.q(_w_10134));
  bfr _b_7677(.a(_w_9579),.q(_w_9580));
  bfr _b_7678(.a(_w_9580),.q(_w_9581));
  bfr _b_7689(.a(_w_9591),.q(_w_9592));
  bfr _b_5432(.a(_w_7334),.q(_w_7335));
  bfr _b_7691(.a(_w_9593),.q(_w_9594));
  bfr _b_12876(.a(_w_14778),.q(_w_14779));
  bfr _b_7692(.a(_w_9594),.q(_w_9595));
  bfr _b_7812(.a(_w_9714),.q(_w_9715));
  bfr _b_7693(.a(_w_9595),.q(_w_9596));
  bfr _b_7697(.a(_w_9599),.q(_w_9600));
  bfr _b_7698(.a(_w_9600),.q(_w_9601));
  bfr _b_7701(.a(_w_9603),.q(_w_9604));
  bfr _b_7704(.a(_w_9606),.q(_w_9607));
  bfr _b_7705(.a(_w_9607),.q(_w_9608));
  bfr _b_13766(.a(_w_15668),.q(_w_15669));
  bfr _b_10469(.a(_w_12371),.q(_w_12372));
  bfr _b_7706(.a(_w_9608),.q(_w_9609));
  bfr _b_10369(.a(_w_12271),.q(_w_12272));
  bfr _b_7707(.a(_w_9609),.q(_w_9610));
  bfr _b_10732(.a(_w_12634),.q(_w_12635));
  spl2 g1169_s_0(.a(n1169),.q0(n1169_0),.q1(n1169_1));
  bfr _b_8840(.a(_w_10742),.q(_w_10743));
  bfr _b_8614(.a(_w_10516),.q(_w_10517));
  bfr _b_7708(.a(_w_9610),.q(_w_9611));
  bfr _b_7709(.a(_w_9611),.q(_w_9612));
  bfr _b_5990(.a(_w_7892),.q(_w_7893));
  bfr _b_7710(.a(_w_9612),.q(_w_9613));
  bfr _b_7712(.a(_w_9614),.q(_w_9615));
  bfr _b_6523(.a(_w_8425),.q(_w_8426));
  bfr _b_7713(.a(_w_9615),.q(_w_9616));
  bfr _b_8374(.a(_w_10276),.q(_w_10277));
  bfr _b_8994(.a(_w_10896),.q(_w_10897));
  bfr _b_7715(.a(_w_9617),.q(_w_9618));
  bfr _b_7718(.a(_w_9620),.q(N6210));
  and_bi g1896(.a(n1887_1),.b(n1890_1),.q(n1896));
  bfr _b_7722(.a(_w_9624),.q(_w_9625));
  bfr _b_6597(.a(_w_8499),.q(_w_8500));
  bfr _b_7723(.a(_w_9625),.q(_w_9626));
  bfr _b_9492(.a(_w_11394),.q(_w_11395));
  bfr _b_7724(.a(_w_9626),.q(_w_9627));
  bfr _b_7726(.a(_w_9628),.q(n144));
  bfr _b_7728(.a(_w_9630),.q(_w_9631));
  bfr _b_4982(.a(_w_6884),.q(_w_6885));
  bfr _b_7827(.a(_w_9729),.q(_w_9730));
  bfr _b_7730(.a(_w_9632),.q(_w_9633));
  bfr _b_8841(.a(_w_10743),.q(_w_10744));
  bfr _b_7731(.a(_w_9633),.q(_w_9634));
  bfr _b_7732(.a(_w_9634),.q(_w_9635));
  bfr _b_12424(.a(_w_14326),.q(_w_14327));
  bfr _b_7733(.a(_w_9635),.q(_w_9636));
  bfr _b_7734(.a(_w_9636),.q(n300));
  bfr _b_11719(.a(_w_13621),.q(_w_13622));
  bfr _b_7739(.a(_w_9641),.q(_w_9642));
  bfr _b_10435(.a(_w_12337),.q(_w_12338));
  or_bb g347(.a(n345_0),.b(n346),.q(n347));
  bfr _b_7742(.a(_w_9644),.q(_w_9645));
  bfr _b_8047(.a(_w_9949),.q(n1102));
  bfr _b_7745(.a(_w_9647),.q(_w_9648));
  bfr _b_7748(.a(_w_9650),.q(_w_9651));
  bfr _b_7749(.a(_w_9651),.q(_w_9652));
  bfr _b_7813(.a(_w_9715),.q(_w_9716));
  bfr _b_11056(.a(_w_12958),.q(_w_12959));
  bfr _b_4997(.a(_w_6899),.q(_w_6900));
  bfr _b_3579(.a(_w_5481),.q(_w_5482));
  bfr _b_7750(.a(_w_9652),.q(_w_9653));
  bfr _b_10485(.a(_w_12387),.q(_w_12388));
  bfr _b_9507(.a(_w_11409),.q(_w_11410));
  bfr _b_7757(.a(_w_9659),.q(n275));
  bfr _b_5929(.a(_w_7831),.q(_w_7832));
  bfr _b_9581(.a(_w_11483),.q(_w_11484));
  bfr _b_13472(.a(_w_15374),.q(_w_15375));
  bfr _b_9956(.a(_w_11858),.q(_w_11859));
  bfr _b_7764(.a(_w_9666),.q(_w_9667));
  bfr _b_5657(.a(_w_7559),.q(_w_7560));
  bfr _b_8011(.a(_w_9913),.q(_w_9914));
  bfr _b_13241(.a(_w_15143),.q(_w_15144));
  bfr _b_7769(.a(_w_9671),.q(_w_9672));
  bfr _b_7770(.a(_w_9672),.q(_w_9673));
  bfr _b_7771(.a(_w_9673),.q(_w_9674));
  bfr _b_6952(.a(_w_8854),.q(_w_8855));
  bfr _b_7772(.a(_w_9674),.q(_w_9675));
  spl2 g1533_s_0(.a(n1533),.q0(n1533_0),.q1(n1533_1));
  bfr _b_7774(.a(_w_9676),.q(_w_9677));
  and_bi g1098(.a(n1097_0),.b(n1068_0),.q(n1098));
  bfr _b_10079(.a(_w_11981),.q(_w_11982));
  bfr _b_10229(.a(_w_12131),.q(_w_12132));
  bfr _b_7776(.a(_w_9678),.q(_w_9679));
  bfr _b_8053(.a(_w_9955),.q(n1119_1));
  bfr _b_7779(.a(_w_9681),.q(_w_9682));
  bfr _b_7781(.a(_w_9683),.q(n1673));
  bfr _b_8179(.a(_w_10081),.q(_w_10082));
  bfr _b_8386(.a(_w_10288),.q(_w_10289));
  bfr _b_7783(.a(_w_9685),.q(n419));
  bfr _b_8319(.a(_w_10221),.q(_w_10222));
  bfr _b_7785(.a(_w_9687),.q(_w_9688));
  bfr _b_7741(.a(_w_9643),.q(_w_9644));
  bfr _b_7786(.a(_w_9688),.q(_w_9689));
  bfr _b_6978(.a(_w_8880),.q(_w_8881));
  spl4L N18_s_3(.a(N18_2),.q0(N18_12),.q1(_w_15489),.q2(_w_15497),.q3(_w_15509));
  bfr _b_7789(.a(_w_9691),.q(_w_9692));
  bfr _b_10834(.a(_w_12736),.q(_w_12737));
  bfr _b_7790(.a(_w_9692),.q(_w_9693));
  bfr _b_7791(.a(_w_9693),.q(_w_9694));
  bfr _b_7792(.a(_w_9694),.q(_w_9695));
  bfr _b_7795(.a(_w_9697),.q(_w_9698));
  bfr _b_7797(.a(_w_9699),.q(_w_9700));
  bfr _b_7798(.a(_w_9700),.q(n142));
  bfr _b_7325(.a(_w_9227),.q(_w_9228));
  bfr _b_8501(.a(_w_10403),.q(_w_10404));
  bfr _b_6286(.a(_w_8188),.q(_w_8189));
  bfr _b_9771(.a(_w_11673),.q(_w_11674));
  bfr _b_7807(.a(_w_9709),.q(_w_9710));
  bfr _b_7808(.a(_w_9710),.q(_w_9711));
  bfr _b_7810(.a(_w_9712),.q(_w_9713));
  bfr _b_7818(.a(_w_9720),.q(_w_9721));
  bfr _b_7326(.a(_w_9228),.q(_w_9229));
  bfr _b_7822(.a(_w_9724),.q(_w_9725));
  bfr _b_11699(.a(_w_13601),.q(_w_13602));
  bfr _b_9975(.a(_w_11877),.q(_w_11878));
  bfr _b_7824(.a(_w_9726),.q(_w_9727));
  and_bi g1161(.a(n1155_1),.b(n1158_1),.q(n1161));
  bfr _b_7826(.a(_w_9728),.q(_w_9729));
  bfr _b_7830(.a(_w_9732),.q(_w_9733));
  and_bi g1696(.a(n1681_1),.b(n1694_1),.q(_w_14115));
  bfr _b_7832(.a(_w_9734),.q(_w_9735));
  bfr _b_11319(.a(_w_13221),.q(_w_13222));
  bfr _b_7833(.a(_w_9735),.q(_w_9736));
  bfr _b_4295(.a(_w_6197),.q(_w_6198));
  bfr _b_8823(.a(_w_10725),.q(_w_10726));
  bfr _b_7672(.a(_w_9574),.q(_w_9575));
  bfr _b_3918(.a(_w_5820),.q(_w_5821));
  bfr _b_7834(.a(_w_9736),.q(_w_9737));
  bfr _b_7837(.a(_w_9739),.q(_w_9740));
  bfr _b_6225(.a(_w_8127),.q(_w_8128));
  bfr _b_7838(.a(_w_9740),.q(_w_9741));
  and_bi g1122(.a(n1121_0),.b(n1060_0),.q(n1122));
  bfr _b_7839(.a(_w_9741),.q(_w_9742));
  bfr _b_7840(.a(_w_9742),.q(_w_9743));
  bfr _b_7841(.a(_w_9743),.q(_w_9744));
  bfr _b_10587(.a(_w_12489),.q(n1120));
  bfr _b_9172(.a(_w_11074),.q(_w_11075));
  bfr _b_7842(.a(_w_9744),.q(_w_9745));
  bfr _b_7844(.a(_w_9746),.q(_w_9747));
  bfr _b_11851(.a(_w_13753),.q(_w_13754));
  and_bi g143(.a(n112_1),.b(n115_1),.q(n143));
  bfr _b_4049(.a(_w_5951),.q(_w_5952));
  bfr _b_7849(.a(_w_9751),.q(_w_9752));
  bfr _b_7850(.a(_w_9752),.q(n960));
  bfr _b_8212(.a(_w_10114),.q(_w_10115));
  bfr _b_10890(.a(_w_12792),.q(_w_12793));
  bfr _b_4617(.a(_w_6519),.q(_w_6520));
  bfr _b_7851(.a(_w_9753),.q(_w_9754));
  bfr _b_12875(.a(_w_14777),.q(_w_14778));
  bfr _b_7856(.a(_w_9758),.q(n454));
  and_bi g1192(.a(n1185_1),.b(n1190_1),.q(_w_12355));
  bfr _b_8418(.a(_w_10320),.q(_w_10321));
  bfr _b_4215(.a(_w_6117),.q(_w_6118));
  bfr _b_7857(.a(_w_9759),.q(_w_9760));
  bfr _b_7859(.a(_w_9761),.q(_w_9762));
  bfr _b_9576(.a(_w_11478),.q(_w_11479));
  bfr _b_7860(.a(_w_9762),.q(_w_9763));
  spl2 g329_s_0(.a(n329),.q0(n329_0),.q1(n329_1));
  bfr _b_7862(.a(_w_9764),.q(_w_9765));
  bfr _b_7864(.a(_w_9766),.q(_w_9767));
  and_bi g915(.a(n826_1),.b(n913_1),.q(_w_8739));
  bfr _b_9929(.a(_w_11831),.q(n298));
  bfr _b_7866(.a(_w_9768),.q(_w_9769));
  bfr _b_11582(.a(_w_13484),.q(_w_13485));
  spl2 g816_s_0(.a(n816),.q0(n816_0),.q1(n816_1));
  bfr _b_4756(.a(_w_6658),.q(_w_6659));
  bfr _b_6957(.a(_w_8859),.q(_w_8860));
  bfr _b_8809(.a(_w_10711),.q(_w_10712));
  bfr _b_9537(.a(_w_11439),.q(_w_11440));
  bfr _b_13123(.a(_w_15025),.q(_w_15026));
  bfr _b_7867(.a(_w_9769),.q(_w_9770));
  bfr _b_7871(.a(_w_9773),.q(_w_9774));
  bfr _b_7872(.a(_w_9774),.q(_w_9775));
  bfr _b_7874(.a(_w_9776),.q(_w_9777));
  bfr _b_4825(.a(_w_6727),.q(_w_6728));
  bfr _b_7875(.a(_w_9777),.q(_w_9778));
  bfr _b_7876(.a(_w_9778),.q(_w_9779));
  bfr _b_7882(.a(_w_9784),.q(_w_9785));
  bfr _b_7883(.a(_w_9785),.q(_w_9786));
  bfr _b_3866(.a(_w_5768),.q(_w_5769));
  bfr _b_7884(.a(_w_9786),.q(_w_9787));
  bfr _b_7885(.a(_w_9787),.q(_w_9788));
  bfr _b_7887(.a(_w_9789),.q(_w_9790));
  bfr _b_6900(.a(_w_8802),.q(_w_8803));
  bfr _b_8796(.a(_w_10698),.q(_w_10699));
  bfr _b_7888(.a(_w_9790),.q(_w_9791));
  bfr _b_6188(.a(_w_8090),.q(_w_8091));
  bfr _b_9254(.a(_w_11156),.q(_w_11157));
  bfr _b_13409(.a(_w_15311),.q(n556));
  bfr _b_7891(.a(_w_9793),.q(_w_9794));
  bfr _b_7892(.a(_w_9794),.q(_w_9795));
  bfr _b_7895(.a(_w_9797),.q(_w_9798));
  bfr _b_7896(.a(_w_9798),.q(_w_9799));
  bfr _b_7110(.a(_w_9012),.q(_w_9013));
  bfr _b_7170(.a(_w_9072),.q(_w_9073));
  bfr _b_7897(.a(_w_9799),.q(_w_9800));
  bfr _b_9596(.a(_w_11498),.q(_w_11499));
  bfr _b_7901(.a(_w_9803),.q(_w_9804));
  bfr _b_7902(.a(_w_9804),.q(_w_9805));
  bfr _b_4074(.a(_w_5976),.q(_w_5977));
  bfr _b_7904(.a(_w_9806),.q(_w_9807));
  bfr _b_7907(.a(_w_9809),.q(_w_9810));
  spl2 g1456_s_0(.a(n1456),.q0(n1456_0),.q1(n1456_1));
  bfr _b_7908(.a(_w_9810),.q(_w_9811));
  spl2 g229_s_0(.a(n229),.q0(n229_0),.q1(n229_1));
  bfr _b_8676(.a(_w_10578),.q(_w_10579));
  bfr _b_13069(.a(_w_14971),.q(_w_14972));
  spl2 g255_s_0(.a(n255),.q0(n255_0),.q1(n255_1));
  bfr _b_5344(.a(_w_7246),.q(_w_7247));
  bfr _b_7914(.a(_w_9816),.q(_w_9817));
  bfr _b_10334(.a(_w_12236),.q(_w_12237));
  bfr _b_4855(.a(_w_6757),.q(_w_6758));
  bfr _b_7915(.a(_w_9817),.q(_w_9818));
  bfr _b_10912(.a(_w_12814),.q(_w_12815));
  bfr _b_7917(.a(_w_9819),.q(_w_9820));
  bfr _b_7918(.a(_w_9820),.q(_w_9821));
  bfr _b_7921(.a(_w_9823),.q(_w_9824));
  bfr _b_7925(.a(_w_9827),.q(_w_9828));
  bfr _b_7926(.a(_w_9828),.q(_w_9829));
  bfr _b_7927(.a(_w_9829),.q(_w_9830));
  bfr _b_7933(.a(_w_9835),.q(_w_9836));
  bfr _b_8794(.a(_w_10696),.q(_w_10697));
  bfr _b_7936(.a(_w_9838),.q(_w_9839));
  bfr _b_7944(.a(_w_9846),.q(_w_9847));
  bfr _b_4544(.a(_w_6446),.q(_w_6447));
  bfr _b_7947(.a(_w_9849),.q(_w_9850));
  bfr _b_7948(.a(_w_9850),.q(_w_9851));
  spl2 g1758_s_0(.a(n1758),.q0(n1758_0),.q1(n1758_1));
  bfr _b_7954(.a(_w_9856),.q(_w_9857));
  bfr _b_7955(.a(_w_9857),.q(_w_9858));
  bfr _b_7957(.a(_w_9859),.q(_w_9860));
  bfr _b_4337(.a(_w_6239),.q(_w_6240));
  bfr _b_7959(.a(_w_9861),.q(_w_9862));
  bfr _b_3795(.a(_w_5697),.q(_w_5698));
  bfr _b_7960(.a(_w_9862),.q(_w_9863));
  spl2 g286_s_0(.a(n286),.q0(n286_0),.q1(_w_6280));
  bfr _b_7963(.a(_w_9865),.q(_w_9866));
  bfr _b_7968(.a(_w_9870),.q(_w_9871));
  bfr _b_7971(.a(_w_9873),.q(_w_9874));
  bfr _b_7974(.a(_w_9876),.q(_w_9877));
  bfr _b_9569(.a(_w_11471),.q(_w_11472));
  bfr _b_6235(.a(_w_8137),.q(_w_8138));
  bfr _b_7975(.a(_w_9877),.q(_w_9878));
  and_bi g211(.a(n210_0),.b(n186_0),.q(n211));
  bfr _b_7976(.a(_w_9878),.q(_w_9879));
  bfr _b_3914(.a(_w_5816),.q(_w_5817));
  bfr _b_7977(.a(_w_9879),.q(_w_9880));
  bfr _b_7981(.a(_w_9883),.q(n815));
  bfr _b_7982(.a(_w_9884),.q(_w_9885));
  bfr _b_13506(.a(_w_15408),.q(_w_15409));
  or_bb g576(.a(n531_0),.b(n575_0),.q(n576));
  bfr _b_10113(.a(_w_12015),.q(_w_12016));
  bfr _b_7988(.a(_w_9890),.q(_w_9891));
  bfr _b_8065(.a(_w_9967),.q(_w_9968));
  bfr _b_3572(.a(_w_5474),.q(_w_5475));
  spl2 g1294_s_0(.a(n1294),.q0(n1294_0),.q1(n1294_1));
  bfr _b_4017(.a(_w_5919),.q(_w_5920));
  bfr _b_9999(.a(_w_11901),.q(_w_11902));
  bfr _b_9105(.a(_w_11007),.q(_w_11008));
  bfr _b_7989(.a(_w_9891),.q(n238));
  bfr _b_5981(.a(_w_7883),.q(_w_7884));
  bfr _b_8802(.a(_w_10704),.q(_w_10705));
  bfr _b_7990(.a(_w_9892),.q(_w_9893));
  bfr _b_7533(.a(_w_9435),.q(_w_9436));
  bfr _b_7991(.a(_w_9893),.q(_w_9894));
  bfr _b_7993(.a(_w_9895),.q(_w_9896));
  bfr _b_7999(.a(_w_9901),.q(_w_9902));
  bfr _b_14204(.a(_w_16106),.q(_w_16107));
  bfr _b_8625(.a(_w_10527),.q(_w_10528));
  bfr _b_8002(.a(_w_9904),.q(_w_9905));
  bfr _b_4922(.a(_w_6824),.q(_w_6825));
  bfr _b_8004(.a(_w_9906),.q(_w_9907));
  bfr _b_8006(.a(_w_9908),.q(_w_9909));
  bfr _b_8007(.a(_w_9909),.q(_w_9910));
  bfr _b_11022(.a(_w_12924),.q(_w_12925));
  spl2 g744_s_0(.a(n744),.q0(n744_0),.q1(n744_1));
  bfr _b_8009(.a(_w_9911),.q(_w_9912));
  bfr _b_3452(.a(_w_5354),.q(_w_5355));
  bfr _b_8010(.a(_w_9912),.q(_w_9913));
  bfr _b_11802(.a(_w_13704),.q(_w_13705));
  spl2 g575_s_0(.a(n575),.q0(n575_0),.q1(n575_1));
  bfr _b_8013(.a(_w_9915),.q(n1365));
  bfr _b_11561(.a(_w_13463),.q(_w_13464));
  bfr _b_8014(.a(_w_9916),.q(_w_9917));
  bfr _b_8018(.a(_w_9920),.q(_w_9921));
  bfr _b_8019(.a(_w_9921),.q(_w_9922));
  spl2 g678_s_0(.a(n678),.q0(n678_0),.q1(n678_1));
  bfr _b_8021(.a(_w_9923),.q(_w_9924));
  bfr _b_8022(.a(_w_9924),.q(_w_9925));
  spl2 g1300_s_0(.a(n1300),.q0(n1300_0),.q1(n1300_1));
  bfr _b_8023(.a(_w_9925),.q(_w_9926));
  bfr _b_8024(.a(_w_9926),.q(_w_9927));
  bfr _b_8028(.a(_w_9930),.q(_w_9931));
  bfr _b_8029(.a(_w_9931),.q(_w_9932));
  bfr _b_8030(.a(_w_9932),.q(_w_9933));
  bfr _b_12379(.a(_w_14281),.q(_w_14282));
  bfr _b_8032(.a(_w_9934),.q(_w_9935));
  bfr _b_7562(.a(_w_9464),.q(_w_9465));
  bfr _b_8034(.a(_w_9936),.q(_w_9937));
  bfr _b_8038(.a(_w_9940),.q(n1666));
  and_bb g238(.a(N358_7),.b(N52_9),.q(_w_9884));
  bfr _b_8040(.a(_w_9942),.q(N290_5));
  bfr _b_10535(.a(_w_12437),.q(_w_12438));
  bfr _b_8043(.a(_w_9945),.q(_w_9946));
  and_bb g1621(.a(N256_12),.b(N409_19),.q(_w_9943));
  bfr _b_8046(.a(_w_9948),.q(n221));
  bfr _b_8048(.a(_w_9950),.q(n116));
  bfr _b_8049(.a(_w_9951),.q(n1474));
  spl2 g45_s_0(.a(n45),.q0(n45_0),.q1(n45_1));
  bfr _b_8051(.a(_w_9953),.q(_w_9954));
  bfr _b_14132(.a(_w_16034),.q(_w_16035));
  bfr _b_11542(.a(_w_13444),.q(_w_13445));
  bfr _b_8052(.a(_w_9954),.q(_w_9955));
  spl2 g469_s_0(.a(n469),.q0(n469_0),.q1(n469_1));
  bfr _b_6518(.a(_w_8420),.q(_w_8421));
  bfr _b_8059(.a(_w_9961),.q(_w_9962));
  bfr _b_13986(.a(_w_15888),.q(_w_15889));
  bfr _b_8060(.a(_w_9962),.q(_w_9963));
  bfr _b_9868(.a(_w_11770),.q(_w_11771));
  bfr _b_8061(.a(_w_9963),.q(_w_9964));
  or_bb g1391(.a(n1389_0),.b(n1390),.q(n1391));
  bfr _b_8064(.a(_w_9966),.q(_w_9967));
  bfr _b_8426(.a(_w_10328),.q(_w_10329));
  bfr _b_8066(.a(_w_9968),.q(_w_9969));
  bfr _b_8067(.a(_w_9969),.q(_w_9970));
  spl2 g1716_s_0(.a(n1716),.q0(n1716_0),.q1(_w_6346));
  and_bb g677(.a(n623_1),.b(n675_1),.q(_w_9248));
  bfr _b_10162(.a(_w_12064),.q(n360));
  bfr _b_6112(.a(_w_8014),.q(_w_8015));
  bfr _b_8072(.a(_w_9974),.q(_w_9975));
  bfr _b_8074(.a(_w_9976),.q(_w_9977));
  bfr _b_7027(.a(_w_8929),.q(_w_8930));
  bfr _b_8076(.a(_w_9978),.q(_w_9979));
  bfr _b_11038(.a(_w_12940),.q(_w_12941));
  bfr _b_8082(.a(_w_9984),.q(_w_9985));
  bfr _b_8083(.a(_w_9985),.q(_w_9986));
  bfr _b_8093(.a(_w_9995),.q(_w_9996));
  bfr _b_8095(.a(_w_9997),.q(_w_9998));
  bfr _b_8098(.a(_w_10000),.q(_w_10001));
  bfr _b_8099(.a(_w_10001),.q(_w_10002));
  bfr _b_8639(.a(_w_10541),.q(_w_10542));
  bfr _b_4490(.a(_w_6392),.q(_w_6393));
  bfr _b_8100(.a(_w_10002),.q(_w_10003));
  bfr _b_8104(.a(_w_10006),.q(_w_10007));
  bfr _b_12106(.a(_w_14008),.q(_w_14009));
  bfr _b_8105(.a(_w_10007),.q(_w_10008));
  bfr _b_8772(.a(_w_10674),.q(_w_10675));
  bfr _b_3587(.a(_w_5489),.q(_w_5490));
  and_bb g376(.a(N137_6),.b(N307_12),.q(_w_9568));
  bfr _b_8106(.a(_w_10008),.q(_w_10009));
  bfr _b_8107(.a(_w_10009),.q(_w_10010));
  bfr _b_8108(.a(_w_10010),.q(_w_10011));
  bfr _b_8110(.a(_w_10012),.q(_w_10013));
  bfr _b_8114(.a(_w_10016),.q(_w_10017));
  bfr _b_4264(.a(_w_6166),.q(_w_6167));
  or_bb g274(.a(n237_0),.b(n273_0),.q(n274));
  bfr _b_5137(.a(_w_7039),.q(_w_7040));
  bfr _b_9910(.a(_w_11812),.q(n540));
  spl2 g926_s_0(.a(n926),.q0(n926_0),.q1(n926_1));
  bfr _b_8115(.a(_w_10017),.q(_w_10018));
  bfr _b_8117(.a(_w_10019),.q(_w_10020));
  spl2 g1380_s_0(.a(n1380),.q0(n1380_0),.q1(n1380_1));
  bfr _b_9043(.a(_w_10945),.q(_w_10946));
  bfr _b_10398(.a(_w_12300),.q(n1131_1));
  bfr _b_8118(.a(_w_10020),.q(_w_10021));
  bfr _b_8120(.a(_w_10022),.q(_w_10023));
  bfr _b_8369(.a(_w_10271),.q(_w_10272));
  bfr _b_12971(.a(_w_14873),.q(_w_14874));
  bfr _b_5402(.a(_w_7304),.q(_w_7305));
  bfr _b_7682(.a(_w_9584),.q(_w_9585));
  bfr _b_8122(.a(_w_10024),.q(_w_10025));
  spl2 g1609_s_0(.a(n1609),.q0(n1609_0),.q1(n1609_1));
  bfr _b_8124(.a(_w_10026),.q(_w_10027));
  bfr _b_8127(.a(_w_10029),.q(_w_10030));
  bfr _b_4374(.a(_w_6276),.q(_w_6277));
  bfr _b_8128(.a(_w_10030),.q(_w_10031));
  bfr _b_8131(.a(_w_10033),.q(_w_10034));
  bfr _b_5527(.a(_w_7429),.q(_w_7430));
  bfr _b_8132(.a(_w_10034),.q(_w_10035));
  bfr _b_8133(.a(_w_10035),.q(_w_10036));
  bfr _b_8139(.a(_w_10041),.q(_w_10042));
  bfr _b_8415(.a(_w_10317),.q(_w_10318));
  bfr _b_8140(.a(_w_10042),.q(_w_10043));
  bfr _b_8141(.a(_w_10043),.q(_w_10044));
  bfr _b_5728(.a(_w_7630),.q(_w_7631));
  bfr _b_8144(.a(_w_10046),.q(_w_10047));
  bfr _b_9455(.a(_w_11357),.q(_w_11358));
  bfr _b_8145(.a(_w_10047),.q(_w_10048));
  bfr _b_13462(.a(_w_15364),.q(_w_15365));
  bfr _b_6718(.a(_w_8620),.q(n935));
  bfr _b_8148(.a(_w_10050),.q(_w_10051));
  bfr _b_8149(.a(_w_10051),.q(_w_10052));
  bfr _b_8154(.a(_w_10056),.q(_w_10057));
  bfr _b_8151(.a(_w_10053),.q(_w_10054));
  bfr _b_8155(.a(_w_10057),.q(_w_10058));
  spl2 g1628_s_0(.a(n1628),.q0(n1628_0),.q1(n1628_1));
  bfr _b_8156(.a(_w_10058),.q(_w_10059));
  bfr _b_8159(.a(_w_10061),.q(_w_10062));
  bfr _b_8160(.a(_w_10062),.q(_w_10063));
  bfr _b_8161(.a(_w_10063),.q(_w_10064));
  bfr _b_8164(.a(_w_10066),.q(_w_10067));
  and_bi g1731(.a(n1710_1),.b(n1713_1),.q(n1731));
  bfr _b_8167(.a(_w_10069),.q(_w_10070));
  bfr _b_9792(.a(_w_11694),.q(_w_11695));
  bfr _b_4957(.a(_w_6859),.q(_w_6860));
  bfr _b_8168(.a(_w_10070),.q(_w_10071));
  spl2 g1738_s_0(.a(n1738),.q0(n1738_0),.q1(n1738_1));
  bfr _b_6295(.a(_w_8197),.q(n1068));
  bfr _b_8169(.a(_w_10071),.q(_w_10072));
  bfr _b_13431(.a(_w_15333),.q(_w_15334));
  bfr _b_9561(.a(_w_11463),.q(_w_11464));
  bfr _b_8173(.a(_w_10075),.q(_w_10076));
  bfr _b_5832(.a(_w_7734),.q(_w_7735));
  bfr _b_8174(.a(_w_10076),.q(_w_10077));
  and_bb g1612(.a(N171_17),.b(N494_14),.q(_w_13958));
  bfr _b_8180(.a(_w_10082),.q(_w_10083));
  bfr _b_9899(.a(_w_11801),.q(_w_11802));
  bfr _b_8187(.a(_w_10089),.q(_w_10090));
  bfr _b_8189(.a(_w_10091),.q(_w_10092));
  bfr _b_8190(.a(_w_10092),.q(_w_10093));
  bfr _b_8191(.a(_w_10093),.q(_w_10094));
  bfr _b_8192(.a(_w_10094),.q(_w_10095));
  bfr _b_8337(.a(_w_10239),.q(_w_10240));
  bfr _b_8193(.a(_w_10095),.q(_w_10096));
  bfr _b_9693(.a(_w_11595),.q(_w_11596));
  bfr _b_8197(.a(_w_10099),.q(_w_10100));
  bfr _b_8198(.a(_w_10100),.q(_w_10101));
  bfr _b_8292(.a(_w_10194),.q(_w_10195));
  bfr _b_10431(.a(_w_12333),.q(n61));
  bfr _b_8201(.a(_w_10103),.q(_w_10104));
  bfr _b_8202(.a(_w_10104),.q(_w_10105));
  bfr _b_13249(.a(_w_15151),.q(_w_15152));
  bfr _b_8207(.a(_w_10109),.q(_w_10110));
  bfr _b_9391(.a(_w_11293),.q(_w_11294));
  bfr _b_8766(.a(_w_10668),.q(_w_10669));
  bfr _b_8208(.a(_w_10110),.q(_w_10111));
  bfr _b_8210(.a(_w_10112),.q(_w_10113));
  bfr _b_8214(.a(_w_10116),.q(_w_10117));
  bfr _b_8215(.a(_w_10117),.q(_w_10118));
  bfr _b_7159(.a(_w_9061),.q(_w_9062));
  bfr _b_10242(.a(_w_12144),.q(_w_12145));
  bfr _b_8216(.a(_w_10118),.q(_w_10119));
  and_bi g768(.a(n766_0),.b(n767),.q(n768));
  bfr _b_8217(.a(_w_10119),.q(_w_10120));
  bfr _b_6000(.a(_w_7902),.q(_w_7903));
  bfr _b_6314(.a(_w_8216),.q(_w_8217));
  bfr _b_8218(.a(_w_10120),.q(_w_10121));
  bfr _b_4551(.a(_w_6453),.q(_w_6454));
  and_bb g109(.a(N273_9),.b(N86_5),.q(n109));
  bfr _b_7065(.a(_w_8967),.q(_w_8968));
  bfr _b_8219(.a(_w_10121),.q(_w_10122));
  bfr _b_9436(.a(_w_11338),.q(_w_11339));
  bfr _b_8220(.a(_w_10122),.q(_w_10123));
  bfr _b_10231(.a(_w_12133),.q(_w_12134));
  bfr _b_8222(.a(_w_10124),.q(_w_10125));
  bfr _b_8224(.a(_w_10126),.q(_w_10127));
  bfr _b_8226(.a(_w_10128),.q(_w_10129));
  bfr _b_8227(.a(_w_10129),.q(_w_10130));
  bfr _b_9730(.a(_w_11632),.q(_w_11633));
  bfr _b_13791(.a(_w_15693),.q(_w_15694));
  bfr _b_11835(.a(_w_13737),.q(_w_13738));
  bfr _b_5040(.a(_w_6942),.q(_w_6943));
  bfr _b_8228(.a(_w_10130),.q(_w_10131));
  bfr _b_5144(.a(_w_7046),.q(_w_7047));
  bfr _b_8229(.a(_w_10131),.q(_w_10132));
  bfr _b_8230(.a(_w_10132),.q(_w_10133));
  bfr _b_5659(.a(_w_7561),.q(_w_7562));
  bfr _b_8232(.a(_w_10134),.q(_w_10135));
  bfr _b_8234(.a(_w_10136),.q(_w_10137));
  bfr _b_12991(.a(_w_14893),.q(_w_14894));
  bfr _b_8236(.a(_w_10138),.q(_w_10139));
  spl2 g382_s_0(.a(n382),.q0(n382_0),.q1(_w_7467));
  bfr _b_4378(.a(_w_6280),.q(_w_6281));
  bfr _b_8237(.a(_w_10139),.q(_w_10140));
  bfr _b_10194(.a(_w_12096),.q(n653));
  bfr _b_8241(.a(_w_10143),.q(_w_10144));
  and_bi g333(.a(n332_0),.b(n300_0),.q(n333));
  or_bb g256(.a(n243_0),.b(n255_0),.q(n256));
  bfr _b_8245(.a(_w_10147),.q(_w_10148));
  bfr _b_8246(.a(_w_10148),.q(N2223));
  and_bb g918(.a(n825_1),.b(n916_1),.q(_w_10441));
  bfr _b_8247(.a(_w_10149),.q(_w_10150));
  bfr _b_9506(.a(_w_11408),.q(_w_11409));
  bfr _b_8249(.a(_w_10151),.q(_w_10152));
  bfr _b_8251(.a(_w_10153),.q(_w_10154));
  bfr _b_8253(.a(_w_10155),.q(_w_10156));
  bfr _b_10248(.a(_w_12150),.q(_w_12151));
  bfr _b_3848(.a(_w_5750),.q(_w_5751));
  bfr _b_4608(.a(_w_6510),.q(_w_6511));
  bfr _b_8259(.a(_w_10161),.q(_w_10162));
  bfr _b_8260(.a(_w_10162),.q(_w_10163));
  bfr _b_5328(.a(_w_7230),.q(_w_7231));
  bfr _b_5325(.a(_w_7227),.q(_w_7228));
  bfr _b_7766(.a(_w_9668),.q(_w_9669));
  bfr _b_8266(.a(_w_10168),.q(_w_10169));
  bfr _b_14225(.a(_w_16127),.q(_w_16128));
  bfr _b_12032(.a(_w_13934),.q(_w_13935));
  bfr _b_8268(.a(_w_10170),.q(_w_10171));
  bfr _b_8271(.a(_w_10173),.q(_w_10174));
  bfr _b_8273(.a(_w_10175),.q(_w_10176));
  bfr _b_8276(.a(_w_10178),.q(_w_10179));
  bfr _b_12019(.a(_w_13921),.q(_w_13922));
  bfr _b_3473(.a(_w_5375),.q(_w_5376));
  bfr _b_8730(.a(_w_10632),.q(_w_10633));
  bfr _b_3922(.a(_w_5824),.q(_w_5825));
  bfr _b_8279(.a(_w_10181),.q(n987));
  bfr _b_8281(.a(_w_10183),.q(n1041));
  bfr _b_13375(.a(_w_15277),.q(_w_15278));
  bfr _b_8282(.a(_w_10184),.q(_w_10185));
  bfr _b_13243(.a(_w_15145),.q(_w_15146));
  bfr _b_3944(.a(_w_5846),.q(_w_5847));
  bfr _b_8284(.a(_w_10186),.q(_w_10187));
  and_bi g345(.a(n344_0),.b(n296_0),.q(n345));
  bfr _b_5899(.a(_w_7801),.q(_w_7802));
  bfr _b_8285(.a(_w_10187),.q(n1404_1));
  bfr _b_8286(.a(_w_10188),.q(_w_10189));
  bfr _b_8287(.a(_w_10189),.q(_w_10190));
  bfr _b_10207(.a(_w_12109),.q(_w_12110));
  bfr _b_8299(.a(_w_10201),.q(n401));
  bfr _b_8302(.a(_w_10204),.q(_w_10205));
  bfr _b_8309(.a(_w_10211),.q(_w_10212));
  bfr _b_9966(.a(_w_11868),.q(_w_11869));
  bfr _b_10986(.a(_w_12888),.q(n1159));
  bfr _b_8310(.a(_w_10212),.q(_w_10213));
  bfr _b_9729(.a(_w_11631),.q(_w_11632));
  bfr _b_8311(.a(_w_10213),.q(_w_10214));
  bfr _b_8617(.a(_w_10519),.q(_w_10520));
  bfr _b_8312(.a(_w_10214),.q(_w_10215));
  bfr _b_11906(.a(_w_13808),.q(_w_13809));
  bfr _b_5263(.a(_w_7165),.q(_w_7166));
  bfr _b_8314(.a(_w_10216),.q(_w_10217));
  bfr _b_12230(.a(_w_14132),.q(_w_14133));
  bfr _b_12072(.a(_w_13974),.q(n766_1));
  bfr _b_7344(.a(_w_9246),.q(n680));
  bfr _b_8315(.a(_w_10217),.q(_w_10218));
  bfr _b_8316(.a(_w_10218),.q(_w_10219));
  bfr _b_8317(.a(_w_10219),.q(_w_10220));
  bfr _b_10096(.a(_w_11998),.q(_w_11999));
  bfr _b_9468(.a(_w_11370),.q(_w_11371));
  bfr _b_8318(.a(_w_10220),.q(_w_10221));
  bfr _b_8320(.a(_w_10222),.q(_w_10223));
  bfr _b_14271(.a(_w_16173),.q(_w_16174));
  bfr _b_12764(.a(_w_14666),.q(_w_14667));
  bfr _b_8324(.a(_w_10226),.q(_w_10227));
  bfr _b_12475(.a(_w_14377),.q(_w_14378));
  bfr _b_8328(.a(_w_10230),.q(_w_10231));
  bfr _b_8329(.a(_w_10231),.q(_w_10232));
  bfr _b_7349(.a(_w_9251),.q(n1654));
  bfr _b_8330(.a(_w_10232),.q(_w_10233));
  and_bb g61(.a(n42_2),.b(n59_1),.q(_w_12333));
  bfr _b_8333(.a(_w_10235),.q(_w_10236));
  bfr _b_13012(.a(_w_14914),.q(_w_14915));
  bfr _b_4555(.a(_w_6457),.q(_w_6458));
  bfr _b_4269(.a(_w_6171),.q(_w_6172));
  bfr _b_8335(.a(_w_10237),.q(_w_10238));
  and_bi g1389(.a(n1388_0),.b(n1383_0),.q(n1389));
  bfr _b_8338(.a(_w_10240),.q(_w_10241));
  bfr _b_11967(.a(_w_13869),.q(_w_13870));
  and_bi g719(.a(n688_1),.b(n691_1),.q(n719));
  bfr _b_8339(.a(_w_10241),.q(_w_10242));
  bfr _b_7330(.a(_w_9232),.q(_w_9233));
  bfr _b_8343(.a(_w_10245),.q(_w_10246));
  bfr _b_11814(.a(_w_13716),.q(_w_13717));
  bfr _b_8345(.a(_w_10247),.q(_w_10248));
  bfr _b_8347(.a(_w_10249),.q(_w_10250));
  bfr _b_8349(.a(_w_10251),.q(_w_10252));
  bfr _b_10968(.a(_w_12870),.q(_w_12871));
  bfr _b_6350(.a(_w_8252),.q(_w_8253));
  bfr _b_8352(.a(_w_10254),.q(_w_10255));
  bfr _b_13589(.a(_w_15491),.q(_w_15492));
  bfr _b_8353(.a(_w_10255),.q(_w_10256));
  bfr _b_8354(.a(_w_10256),.q(_w_10257));
  bfr _b_8355(.a(_w_10257),.q(_w_10258));
  bfr _b_13041(.a(_w_14943),.q(_w_14944));
  bfr _b_8357(.a(_w_10259),.q(_w_10260));
  or_bb g1241(.a(n1239_0),.b(n1240),.q(n1241));
  and_bi g1591(.a(n1590_0),.b(n1537_0),.q(n1591));
  bfr _b_8358(.a(_w_10260),.q(_w_10261));
  bfr _b_8360(.a(_w_10262),.q(_w_10263));
  bfr _b_8361(.a(_w_10263),.q(_w_10264));
  bfr _b_6447(.a(_w_8349),.q(_w_8350));
  bfr _b_8362(.a(_w_10264),.q(_w_10265));
  bfr _b_8363(.a(_w_10265),.q(_w_10266));
  bfr _b_12639(.a(_w_14541),.q(_w_14542));
  bfr _b_8365(.a(_w_10267),.q(_w_10268));
  bfr _b_8366(.a(_w_10268),.q(_w_10269));
  bfr _b_4366(.a(_w_6268),.q(_w_6269));
  bfr _b_8367(.a(_w_10269),.q(_w_10270));
  bfr _b_10546(.a(_w_12448),.q(_w_12449));
  bfr _b_8371(.a(_w_10273),.q(_w_10274));
  bfr _b_8373(.a(_w_10275),.q(_w_10276));
  bfr _b_8376(.a(_w_10278),.q(_w_10279));
  bfr _b_6587(.a(_w_8489),.q(_w_8490));
  bfr _b_8377(.a(_w_10279),.q(_w_10280));
  spl2 g955_s_0(.a(n955),.q0(n955_0),.q1(n955_1));
  bfr _b_8378(.a(_w_10280),.q(_w_10281));
  bfr _b_5603(.a(_w_7505),.q(_w_7506));
  bfr _b_6827(.a(_w_8729),.q(n921));
  bfr _b_8379(.a(_w_10281),.q(_w_10282));
  bfr _b_9759(.a(_w_11661),.q(_w_11662));
  bfr _b_8381(.a(_w_10283),.q(n1231));
  bfr _b_8479(.a(_w_10381),.q(_w_10382));
  bfr _b_4620(.a(_w_6522),.q(_w_6523));
  bfr _b_8762(.a(_w_10664),.q(_w_10665));
  bfr _b_3591(.a(_w_5493),.q(_w_5494));
  bfr _b_10116(.a(_w_12018),.q(_w_12019));
  bfr _b_8382(.a(_w_10284),.q(_w_10285));
  bfr _b_12256(.a(_w_14158),.q(_w_14159));
  bfr _b_8383(.a(_w_10285),.q(_w_10286));
  and_bi g951(.a(n881_1),.b(n884_1),.q(n951));
  bfr _b_4179(.a(_w_6081),.q(_w_6082));
  bfr _b_8384(.a(_w_10286),.q(_w_10287));
  bfr _b_12833(.a(_w_14735),.q(_w_14736));
  bfr _b_9615(.a(_w_11517),.q(_w_11518));
  bfr _b_11687(.a(_w_13589),.q(_w_13590));
  bfr _b_8387(.a(_w_10289),.q(_w_10290));
  bfr _b_8388(.a(_w_10290),.q(_w_10291));
  bfr _b_8392(.a(_w_10294),.q(_w_10295));
  bfr _b_4438(.a(_w_6340),.q(_w_6341));
  bfr _b_8396(.a(_w_10298),.q(n668));
  bfr _b_11550(.a(_w_13452),.q(_w_13453));
  bfr _b_8397(.a(_w_10299),.q(_w_10300));
  bfr _b_8403(.a(_w_10305),.q(n346));
  bfr _b_10146(.a(_w_12048),.q(_w_12049));
  bfr _b_8404(.a(_w_10306),.q(n257));
  bfr _b_8405(.a(_w_10307),.q(_w_10308));
  bfr _b_8406(.a(_w_10308),.q(_w_10309));
  bfr _b_8407(.a(_w_10309),.q(_w_10310));
  bfr _b_3468(.a(_w_5370),.q(N52_11));
  bfr _b_8408(.a(_w_10310),.q(_w_10311));
  bfr _b_6288(.a(_w_8190),.q(_w_8191));
  bfr _b_8410(.a(_w_10312),.q(_w_10313));
  bfr _b_9382(.a(_w_11284),.q(_w_11285));
  bfr _b_8411(.a(_w_10313),.q(_w_10314));
  bfr _b_8412(.a(_w_10314),.q(_w_10315));
  bfr _b_13831(.a(_w_15733),.q(_w_15734));
  bfr _b_12650(.a(_w_14552),.q(_w_14553));
  spl2 g360_s_0(.a(n360),.q0(n360_0),.q1(n360_1));
  bfr _b_8413(.a(_w_10315),.q(_w_10316));
  bfr _b_9923(.a(_w_11825),.q(_w_11826));
  bfr _b_10132(.a(_w_12034),.q(n512));
  bfr _b_8414(.a(_w_10316),.q(_w_10317));
  and_bi g1080(.a(n1079_0),.b(n1074_0),.q(n1080));
  bfr _b_9582(.a(_w_11484),.q(_w_11485));
  bfr _b_8417(.a(_w_10319),.q(_w_10320));
  spl2 g1170_s_0(.a(n1170),.q0(n1170_0),.q1(n1170_1));
  bfr _b_8422(.a(_w_10324),.q(_w_10325));
  bfr _b_5074(.a(_w_6976),.q(_w_6977));
  bfr _b_9701(.a(_w_11603),.q(_w_11604));
  bfr _b_8428(.a(_w_10330),.q(_w_10331));
  bfr _b_8430(.a(_w_10332),.q(_w_10333));
  bfr _b_8433(.a(_w_10335),.q(_w_10336));
  bfr _b_13017(.a(_w_14919),.q(_w_14920));
  bfr _b_8435(.a(_w_10337),.q(_w_10338));
  bfr _b_8437(.a(_w_10339),.q(_w_10340));
  bfr _b_11060(.a(_w_12962),.q(_w_12963));
  bfr _b_8440(.a(_w_10342),.q(_w_10343));
  bfr _b_10467(.a(_w_12369),.q(_w_12370));
  bfr _b_9583(.a(_w_11485),.q(_w_11486));
  bfr _b_14369(.a(_w_16271),.q(_w_16272));
  and_bb g190(.a(N307_9),.b(N86_6),.q(_w_11631));
  bfr _b_8442(.a(_w_10344),.q(_w_10345));
  and_bb g954(.a(N171_10),.b(N375_14),.q(_w_10864));
  bfr _b_4557(.a(_w_6459),.q(_w_6460));
  bfr _b_9166(.a(_w_11068),.q(n924));
  bfr _b_8448(.a(_w_10350),.q(_w_10351));
  bfr _b_13531(.a(_w_15433),.q(_w_15434));
  bfr _b_8452(.a(_w_10354),.q(_w_10355));
  bfr _b_8453(.a(_w_10355),.q(_w_10356));
  bfr _b_8717(.a(_w_10619),.q(n52));
  bfr _b_8454(.a(_w_10356),.q(_w_10357));
  bfr _b_8460(.a(_w_10362),.q(_w_10363));
  spl2 g1121_s_0(.a(n1121),.q0(n1121_0),.q1(n1121_1));
  bfr _b_8461(.a(_w_10363),.q(_w_10364));
  bfr _b_8462(.a(_w_10364),.q(_w_10365));
  bfr _b_8463(.a(_w_10365),.q(_w_10366));
  bfr _b_12349(.a(_w_14251),.q(_w_14252));
  bfr _b_8469(.a(_w_10371),.q(_w_10372));
  bfr _b_8471(.a(_w_10373),.q(_w_10374));
  bfr _b_8472(.a(_w_10374),.q(_w_10375));
  bfr _b_8475(.a(_w_10377),.q(_w_10378));
  bfr _b_10227(.a(_w_12129),.q(_w_12130));
  bfr _b_10549(.a(_w_12451),.q(_w_12452));
  bfr _b_6726(.a(_w_8628),.q(_w_8629));
  bfr _b_8478(.a(_w_10380),.q(_w_10381));
  bfr _b_3737(.a(_w_5639),.q(_w_5640));
  bfr _b_8480(.a(_w_10382),.q(_w_10383));
  bfr _b_8481(.a(_w_10383),.q(_w_10384));
  bfr _b_3411(.a(_w_5313),.q(_w_5314));
  spl2 g1101_s_0(.a(n1101),.q0(n1101_0),.q1(_w_14298));
  bfr _b_8482(.a(_w_10384),.q(_w_10385));
  bfr _b_11890(.a(_w_13792),.q(_w_13793));
  bfr _b_8483(.a(_w_10385),.q(_w_10386));
  or_bb g1581(.a(n1579_0),.b(n1580),.q(n1581));
  bfr _b_8489(.a(_w_10391),.q(_w_10392));
  bfr _b_10221(.a(_w_12123),.q(_w_12124));
  bfr _b_8484(.a(_w_10386),.q(_w_10387));
  bfr _b_11630(.a(_w_13532),.q(_w_13533));
  bfr _b_8486(.a(_w_10388),.q(_w_10389));
  bfr _b_8565(.a(_w_10467),.q(_w_10468));
  bfr _b_8843(.a(_w_10745),.q(_w_10746));
  bfr _b_8487(.a(_w_10389),.q(_w_10390));
  bfr _b_8492(.a(_w_10394),.q(_w_10395));
  bfr _b_8496(.a(_w_10398),.q(_w_10399));
  bfr _b_8497(.a(_w_10399),.q(_w_10400));
  bfr _b_3498(.a(_w_5400),.q(_w_5401));
  bfr _b_6646(.a(_w_8548),.q(_w_8549));
  bfr _b_5839(.a(_w_7741),.q(_w_7742));
  bfr _b_8498(.a(_w_10400),.q(_w_10401));
  bfr _b_13675(.a(_w_15577),.q(_w_15578));
  and_bi g1860(.a(n1858_0),.b(n1859),.q(n1860));
  bfr _b_8600(.a(_w_10502),.q(_w_10503));
  bfr _b_8500(.a(_w_10402),.q(_w_10403));
  bfr _b_8504(.a(_w_10406),.q(_w_10407));
  or_bb g657(.a(n655_0),.b(n656),.q(n657));
  bfr _b_8507(.a(_w_10409),.q(_w_10410));
  bfr _b_8510(.a(_w_10412),.q(_w_10413));
  bfr _b_9855(.a(_w_11757),.q(_w_11758));
  bfr _b_6068(.a(_w_7970),.q(_w_7971));
  bfr _b_8511(.a(_w_10413),.q(_w_10414));
  bfr _b_4359(.a(_w_6261),.q(_w_6262));
  bfr _b_8512(.a(_w_10414),.q(_w_10415));
  bfr _b_12980(.a(_w_14882),.q(_w_14883));
  bfr _b_8513(.a(_w_10415),.q(_w_10416));
  bfr _b_8514(.a(_w_10416),.q(_w_10417));
  bfr _b_8518(.a(_w_10420),.q(_w_10421));
  bfr _b_8519(.a(_w_10421),.q(_w_10422));
  spl4L N392_s_3(.a(N392_2),.q0(N392_12),.q1(N392_13),.q2(N392_14),.q3(N392_15));
  bfr _b_8522(.a(_w_10424),.q(_w_10425));
  bfr _b_10489(.a(_w_12391),.q(_w_12392));
  bfr _b_8523(.a(_w_10425),.q(_w_10426));
  and_bi g891(.a(n834_1),.b(n889_1),.q(_w_10628));
  bfr _b_8526(.a(_w_10428),.q(_w_10429));
  spl4L N324_s_0(.a(_w_15542),.q0(N324_0),.q1(N324_1),.q2(N324_2),.q3(N324_3));
  bfr _b_5777(.a(_w_7679),.q(N222_5));
  bfr _b_8528(.a(_w_10430),.q(_w_10431));
  bfr _b_12431(.a(_w_14333),.q(_w_14334));
  bfr _b_8531(.a(_w_10433),.q(_w_10434));
  bfr _b_8952(.a(_w_10854),.q(_w_10855));
  bfr _b_8536(.a(_w_10438),.q(N3211));
  bfr _b_13381(.a(_w_15283),.q(_w_15284));
  bfr _b_8537(.a(_w_10439),.q(n479));
  spl2 g1527_s_0(.a(n1527),.q0(n1527_0),.q1(_w_10574));
  bfr _b_6775(.a(_w_8677),.q(_w_8678));
  bfr _b_8540(.a(_w_10442),.q(n562));
  bfr _b_8541(.a(_w_10443),.q(_w_10444));
  bfr _b_8544(.a(_w_10446),.q(_w_10447));
  bfr _b_8892(.a(_w_10794),.q(_w_10795));
  bfr _b_8546(.a(_w_10448),.q(_w_10449));
  bfr _b_8547(.a(_w_10449),.q(_w_10450));
  spl2 g100_s_0(.a(n100),.q0(n100_0),.q1(n100_1));
  bfr _b_8548(.a(_w_10450),.q(n1070));
  bfr _b_10294(.a(_w_12196),.q(_w_12197));
  bfr _b_8553(.a(_w_10455),.q(_w_10456));
  bfr _b_13569(.a(_w_15471),.q(_w_15472));
  bfr _b_10616(.a(_w_12518),.q(n515));
  bfr _b_8561(.a(_w_10463),.q(_w_10464));
  bfr _b_8562(.a(_w_10464),.q(_w_10465));
  bfr _b_8568(.a(_w_10470),.q(_w_10471));
  bfr _b_8569(.a(_w_10471),.q(_w_10472));
  bfr _b_8570(.a(_w_10472),.q(_w_10473));
  bfr _b_11826(.a(_w_13728),.q(_w_13729));
  and_bi g1851(.a(n1845_1),.b(n1848_1),.q(n1851));
  bfr _b_9248(.a(_w_11150),.q(_w_11151));
  bfr _b_8572(.a(_w_10474),.q(_w_10475));
  bfr _b_8573(.a(_w_10475),.q(_w_10476));
  bfr _b_8443(.a(_w_10345),.q(_w_10346));
  bfr _b_8575(.a(_w_10477),.q(_w_10478));
  bfr _b_10252(.a(_w_12154),.q(_w_12155));
  bfr _b_8576(.a(_w_10478),.q(_w_10479));
  and_bi g185(.a(n162_1),.b(n165_1),.q(n185));
  bfr _b_8581(.a(_w_10483),.q(_w_10484));
  bfr _b_8582(.a(_w_10484),.q(_w_10485));
  or_bb g1047(.a(n1045_1),.b(n935_1),.q(_w_8748));
  bfr _b_8587(.a(_w_10489),.q(_w_10490));
  and_bi g758(.a(n732_1),.b(n756_1),.q(_w_9136));
  bfr _b_8588(.a(_w_10490),.q(_w_10491));
  bfr _b_12620(.a(_w_14522),.q(n1795));
  bfr _b_8589(.a(_w_10491),.q(_w_10492));
  bfr _b_12071(.a(_w_13973),.q(_w_13974));
  spl2 g523_s_0(.a(n523),.q0(n523_0),.q1(n523_1));
  bfr _b_8590(.a(_w_10492),.q(_w_10493));
  spl4L N409_s_2(.a(N409_1),.q0(N409_8),.q1(N409_9),.q2(N409_10),.q3(N409_11));
  bfr _b_7853(.a(_w_9755),.q(_w_9756));
  bfr _b_8591(.a(_w_10493),.q(_w_10494));
  bfr _b_8601(.a(_w_10503),.q(_w_10504));
  bfr _b_13309(.a(_w_15211),.q(_w_15212));
  bfr _b_8602(.a(_w_10504),.q(_w_10505));
  bfr _b_9926(.a(_w_11828),.q(_w_11829));
  bfr _b_8646(.a(_w_10548),.q(_w_10549));
  bfr _b_8608(.a(_w_10510),.q(_w_10511));
  bfr _b_11983(.a(_w_13885),.q(n1525));
  bfr _b_11586(.a(_w_13488),.q(_w_13489));
  bfr _b_11027(.a(_w_12929),.q(n1165));
  bfr _b_8610(.a(_w_10512),.q(_w_10513));
  bfr _b_9911(.a(_w_11813),.q(n1769));
  bfr _b_7514(.a(_w_9416),.q(_w_9417));
  bfr _b_8611(.a(_w_10513),.q(_w_10514));
  bfr _b_13931(.a(_w_15833),.q(_w_15834));
  bfr _b_8613(.a(_w_10515),.q(_w_10516));
  bfr _b_13643(.a(N341),.q(_w_15546));
  bfr _b_11069(.a(_w_12971),.q(_w_12972));
  bfr _b_8714(.a(_w_10616),.q(_w_10617));
  bfr _b_8615(.a(_w_10517),.q(_w_10518));
  bfr _b_12794(.a(_w_14696),.q(_w_14697));
  bfr _b_8618(.a(_w_10520),.q(_w_10521));
  bfr _b_4794(.a(_w_6696),.q(_w_6697));
  bfr _b_5837(.a(_w_7739),.q(_w_7740));
  bfr _b_8620(.a(_w_10522),.q(_w_10523));
  bfr _b_5880(.a(_w_7782),.q(_w_7783));
  bfr _b_8621(.a(_w_10523),.q(_w_10524));
  bfr _b_8626(.a(_w_10528),.q(_w_10529));
  bfr _b_14045(.a(_w_15947),.q(_w_15948));
  bfr _b_10465(.a(_w_12367),.q(n1519));
  bfr _b_8967(.a(_w_10869),.q(_w_10870));
  bfr _b_9347(.a(_w_11249),.q(_w_11250));
  bfr _b_8633(.a(_w_10535),.q(_w_10536));
  bfr _b_11572(.a(_w_13474),.q(_w_13475));
  bfr _b_8634(.a(_w_10536),.q(_w_10537));
  or_bb g575(.a(n573_0),.b(n574),.q(n575));
  bfr _b_7738(.a(_w_9640),.q(n1298));
  bfr _b_8635(.a(_w_10537),.q(_w_10538));
  bfr _b_8636(.a(_w_10538),.q(_w_10539));
  bfr _b_6118(.a(_w_8020),.q(_w_8021));
  bfr _b_8640(.a(_w_10542),.q(_w_10543));
  bfr _b_8641(.a(_w_10543),.q(_w_10544));
  bfr _b_8642(.a(_w_10544),.q(_w_10545));
  bfr _b_4850(.a(_w_6752),.q(_w_6753));
  bfr _b_6421(.a(_w_8323),.q(_w_8324));
  bfr _b_9769(.a(_w_11671),.q(_w_11672));
  bfr _b_8644(.a(_w_10546),.q(_w_10547));
  bfr _b_8649(.a(_w_10551),.q(_w_10552));
  bfr _b_8650(.a(_w_10552),.q(_w_10553));
  bfr _b_3672(.a(_w_5574),.q(_w_5575));
  bfr _b_8654(.a(_w_10556),.q(_w_10557));
  bfr _b_8661(.a(_w_10563),.q(_w_10564));
  bfr _b_8655(.a(_w_10557),.q(_w_10558));
  bfr _b_8659(.a(_w_10561),.q(_w_10562));
  bfr _b_8663(.a(_w_10565),.q(n89));
  bfr _b_9096(.a(_w_10998),.q(_w_10999));
  bfr _b_8665(.a(_w_10567),.q(_w_10568));
  bfr _b_8669(.a(_w_10571),.q(n416));
  bfr _b_8675(.a(_w_10577),.q(_w_10578));
  bfr _b_8680(.a(_w_10582),.q(_w_10583));
  or_bb g1302(.a(n1300_0),.b(n1301),.q(n1302));
  bfr _b_8683(.a(_w_10585),.q(_w_10586));
  bfr _b_8684(.a(_w_10586),.q(_w_10587));
  bfr _b_11167(.a(_w_13069),.q(_w_13070));
  bfr _b_8686(.a(_w_10588),.q(_w_10589));
  bfr _b_8690(.a(_w_10592),.q(_w_10593));
  bfr _b_8871(.a(_w_10773),.q(_w_10774));
  bfr _b_8691(.a(_w_10593),.q(n1527_1));
  and_bi g1233(.a(n1232_0),.b(n1171_0),.q(n1233));
  bfr _b_8693(.a(_w_10595),.q(n806));
  bfr _b_5308(.a(_w_7210),.q(_w_7211));
  bfr _b_8694(.a(_w_10596),.q(_w_10597));
  bfr _b_8695(.a(_w_10597),.q(_w_10598));
  bfr _b_10820(.a(_w_12722),.q(_w_12723));
  spl2 g597_s_0(.a(n597),.q0(n597_0),.q1(n597_1));
  and_bi g829(.a(n790_1),.b(n793_1),.q(n829));
  spl2 g1271_s_0(.a(n1271),.q0(n1271_0),.q1(n1271_1));
  bfr _b_9427(.a(_w_11329),.q(_w_11330));
  bfr _b_12290(.a(_w_14192),.q(_w_14193));
  bfr _b_8698(.a(_w_10600),.q(_w_10601));
  bfr _b_8699(.a(_w_10601),.q(_w_10602));
  bfr _b_8700(.a(_w_10602),.q(_w_10603));
  bfr _b_9317(.a(_w_11219),.q(_w_11220));
  and_bi g1678(.a(n1641_1),.b(n1644_1),.q(n1678));
  spl2 g1293_s_0(.a(n1293),.q0(n1293_0),.q1(n1293_1));
  and_bb g440(.a(N35_13),.b(N426_6),.q(n440));
  bfr _b_8702(.a(_w_10604),.q(_w_10605));
  bfr _b_8703(.a(_w_10605),.q(n76));
  spl2 g1175_s_0(.a(n1175),.q0(n1175_0),.q1(n1175_1));
  bfr _b_8705(.a(_w_10607),.q(_w_10608));
  bfr _b_4427(.a(_w_6329),.q(n36_0));
  bfr _b_8708(.a(_w_10610),.q(_w_10611));
  bfr _b_5518(.a(_w_7420),.q(_w_7421));
  bfr _b_8709(.a(_w_10611),.q(_w_10612));
  bfr _b_8716(.a(_w_10618),.q(_w_10619));
  bfr _b_8718(.a(_w_10620),.q(n659));
  bfr _b_9443(.a(_w_11345),.q(_w_11346));
  bfr _b_11642(.a(_w_13544),.q(_w_13545));
  bfr _b_8720(.a(_w_10622),.q(n44));
  bfr _b_10573(.a(_w_12475),.q(_w_12476));
  bfr _b_8723(.a(_w_10625),.q(n972));
  bfr _b_8725(.a(_w_10627),.q(n197));
  bfr _b_8727(.a(_w_10629),.q(_w_10630));
  and_bi g217(.a(n216_0),.b(n184_0),.q(n217));
  bfr _b_8495(.a(_w_10397),.q(_w_10398));
  bfr _b_8729(.a(_w_10631),.q(_w_10632));
  bfr _b_8731(.a(_w_10633),.q(_w_10634));
  bfr _b_12896(.a(_w_14798),.q(_w_14799));
  bfr _b_9068(.a(_w_10970),.q(_w_10971));
  bfr _b_8734(.a(_w_10636),.q(_w_10637));
  spl4L N443_s_4(.a(N443_3),.q0(N443_16),.q1(N443_17),.q2(N443_18),.q3(N443_19));
  bfr _b_5946(.a(_w_7848),.q(_w_7849));
  bfr _b_8738(.a(_w_10640),.q(_w_10641));
  bfr _b_4493(.a(_w_6395),.q(_w_6396));
  spl2 g97_s_0(.a(n97),.q0(n97_0),.q1(n97_1));
  bfr _b_7516(.a(_w_9418),.q(_w_9419));
  bfr _b_8739(.a(_w_10641),.q(_w_10642));
  bfr _b_13763(.a(_w_15665),.q(_w_15666));
  bfr _b_8741(.a(_w_10643),.q(_w_10644));
  bfr _b_5914(.a(_w_7816),.q(_w_7817));
  bfr _b_8742(.a(_w_10644),.q(n136));
  bfr _b_8743(.a(_w_10645),.q(_w_10646));
  bfr _b_8744(.a(_w_10646),.q(_w_10647));
  bfr _b_8746(.a(_w_10648),.q(_w_10649));
  or_bb g985(.a(n983_0),.b(n984),.q(n985));
  bfr _b_10159(.a(_w_12061),.q(_w_12062));
  bfr _b_8747(.a(_w_10649),.q(_w_10650));
  bfr _b_14351(.a(_w_16253),.q(_w_16254));
  bfr _b_5045(.a(_w_6947),.q(_w_6948));
  bfr _b_8750(.a(_w_10652),.q(_w_10653));
  bfr _b_8390(.a(_w_10292),.q(_w_10293));
  bfr _b_8754(.a(_w_10656),.q(_w_10657));
  bfr _b_5800(.a(_w_7702),.q(_w_7703));
  bfr _b_8758(.a(_w_10660),.q(n182));
  bfr _b_5347(.a(_w_7249),.q(_w_7250));
  bfr _b_9380(.a(_w_11282),.q(_w_11283));
  bfr _b_8761(.a(_w_10663),.q(_w_10664));
  bfr _b_8764(.a(_w_10666),.q(_w_10667));
  bfr _b_8767(.a(_w_10669),.q(_w_10670));
  bfr _b_8768(.a(_w_10670),.q(_w_10671));
  bfr _b_5312(.a(_w_7214),.q(_w_7215));
  bfr _b_8771(.a(_w_10673),.q(_w_10674));
  bfr _b_5102(.a(_w_7004),.q(_w_7005));
  bfr _b_8775(.a(_w_10677),.q(_w_10678));
  and_bi g1121(.a(n1119_0),.b(n1120),.q(n1121));
  bfr _b_8779(.a(_w_10681),.q(_w_10682));
  and_bb g35(.a(N545_1),.b(n33_0),.q(n35));
  bfr _b_8781(.a(_w_10683),.q(_w_10684));
  bfr _b_11098(.a(_w_13000),.q(n1204));
  bfr _b_6220(.a(_w_8122),.q(n594_1));
  bfr _b_8782(.a(_w_10684),.q(_w_10685));
  spl2 g699_s_0(.a(n699),.q0(n699_0),.q1(n699_1));
  bfr _b_5212(.a(_w_7114),.q(_w_7115));
  bfr _b_8783(.a(_w_10685),.q(_w_10686));
  spl2 g872_s_0(.a(n872),.q0(n872_0),.q1(n872_1));
  bfr _b_8819(.a(_w_10721),.q(_w_10722));
  bfr _b_8785(.a(_w_10687),.q(_w_10688));
  bfr _b_7900(.a(_w_9802),.q(_w_9803));
  bfr _b_8790(.a(_w_10692),.q(_w_10693));
  bfr _b_8791(.a(_w_10693),.q(_w_10694));
  bfr _b_8185(.a(_w_10087),.q(_w_10088));
  bfr _b_8798(.a(_w_10700),.q(_w_10701));
  bfr _b_8801(.a(_w_10703),.q(_w_10704));
  bfr _b_13417(.a(_w_15319),.q(_w_15320));
  bfr _b_8803(.a(_w_10705),.q(_w_10706));
  bfr _b_13139(.a(_w_15041),.q(_w_15042));
  bfr _b_8810(.a(_w_10712),.q(_w_10713));
  bfr _b_12244(.a(_w_14146),.q(_w_14147));
  bfr _b_9098(.a(_w_11000),.q(_w_11001));
  bfr _b_7768(.a(_w_9670),.q(_w_9671));
  bfr _b_8811(.a(_w_10713),.q(_w_10714));
  bfr _b_7568(.a(_w_9470),.q(_w_9471));
  bfr _b_8812(.a(_w_10714),.q(_w_10715));
  bfr _b_11661(.a(_w_13563),.q(_w_13564));
  bfr _b_4512(.a(_w_6414),.q(_w_6415));
  bfr _b_9216(.a(_w_11118),.q(_w_11119));
  bfr _b_8813(.a(_w_10715),.q(_w_10716));
  bfr _b_8821(.a(_w_10723),.q(_w_10724));
  bfr _b_9666(.a(_w_11568),.q(_w_11569));
  bfr _b_8751(.a(_w_10653),.q(_w_10654));
  bfr _b_8822(.a(_w_10724),.q(_w_10725));
  bfr _b_12307(.a(_w_14209),.q(_w_14210));
  bfr _b_9728(.a(_w_11630),.q(n1141));
  bfr _b_8824(.a(_w_10726),.q(_w_10727));
  bfr _b_7638(.a(_w_9540),.q(N120_3));
  bfr _b_8826(.a(_w_10728),.q(_w_10729));
  bfr _b_8827(.a(_w_10729),.q(_w_10730));
  spl2 g443_s_0(.a(n443),.q0(n443_0),.q1(n443_1));
  bfr _b_6211(.a(_w_8113),.q(_w_8114));
  bfr _b_8829(.a(_w_10731),.q(_w_10732));
  and_bb g473(.a(n451_1),.b(n471_1),.q(_w_10573));
  bfr _b_9417(.a(_w_11319),.q(_w_11320));
  bfr _b_11742(.a(_w_13644),.q(_w_13645));
  bfr _b_5107(.a(_w_7009),.q(_w_7010));
  bfr _b_8830(.a(_w_10732),.q(_w_10733));
  bfr _b_8839(.a(_w_10741),.q(_w_10742));
  bfr _b_8842(.a(_w_10744),.q(_w_10745));
  bfr _b_5715(.a(_w_7617),.q(_w_7618));
  bfr _b_8846(.a(_w_10748),.q(_w_10749));
  and_bb g1102(.a(n1067_1),.b(n1100_1),.q(_w_9949));
  bfr _b_8848(.a(_w_10750),.q(_w_10751));
  or_bb g1806(.a(n1780_0),.b(n1805_0),.q(n1806));
  bfr _b_8850(.a(_w_10752),.q(_w_10753));
  bfr _b_12452(.a(_w_14354),.q(_w_14355));
  bfr _b_12277(.a(_w_14179),.q(_w_14180));
  bfr _b_8851(.a(_w_10753),.q(_w_10754));
  bfr _b_8852(.a(_w_10754),.q(_w_10755));
  bfr _b_13436(.a(_w_15338),.q(_w_15339));
  bfr _b_8854(.a(_w_10756),.q(_w_10757));
  bfr _b_8855(.a(_w_10757),.q(_w_10758));
  bfr _b_8856(.a(_w_10758),.q(_w_10759));
  bfr _b_3576(.a(_w_5478),.q(_w_5479));
  bfr _b_5030(.a(_w_6932),.q(_w_6933));
  bfr _b_8857(.a(_w_10759),.q(_w_10760));
  bfr _b_8862(.a(_w_10764),.q(_w_10765));
  bfr _b_8863(.a(_w_10765),.q(_w_10766));
  bfr _b_8864(.a(_w_10766),.q(_w_10767));
  bfr _b_12828(.a(_w_14730),.q(_w_14731));
  bfr _b_6363(.a(_w_8265),.q(_w_8266));
  bfr _b_9906(.a(_w_11808),.q(_w_11809));
  bfr _b_8865(.a(_w_10767),.q(_w_10768));
  bfr _b_4174(.a(_w_6076),.q(_w_6077));
  bfr _b_8866(.a(_w_10768),.q(_w_10769));
  bfr _b_8867(.a(_w_10769),.q(_w_10770));
  or_bb g807(.a(n805_0),.b(n806),.q(n807));
  bfr _b_8868(.a(_w_10770),.q(_w_10771));
  bfr _b_13910(.a(_w_15812),.q(_w_15813));
  bfr _b_8872(.a(_w_10774),.q(_w_10775));
  bfr _b_10101(.a(_w_12003),.q(_w_12004));
  bfr _b_8873(.a(_w_10775),.q(_w_10776));
  bfr _b_8874(.a(_w_10776),.q(_w_10777));
  bfr _b_8878(.a(_w_10780),.q(n1334));
  bfr _b_10855(.a(_w_12757),.q(_w_12758));
  bfr _b_8879(.a(_w_10781),.q(_w_10782));
  bfr _b_9486(.a(_w_11388),.q(_w_11389));
  bfr _b_4177(.a(_w_6079),.q(_w_6080));
  bfr _b_8881(.a(_w_10783),.q(_w_10784));
  bfr _b_11709(.a(_w_13611),.q(_w_13612));
  bfr _b_3641(.a(_w_5543),.q(_w_5544));
  bfr _b_8883(.a(_w_10785),.q(_w_10786));
  bfr _b_8886(.a(_w_10788),.q(_w_10789));
  bfr _b_9853(.a(_w_11755),.q(_w_11756));
  spl2 g1491_s_0(.a(n1491),.q0(n1491_0),.q1(_w_15048));
  bfr _b_8887(.a(_w_10789),.q(_w_10790));
  bfr _b_8888(.a(_w_10790),.q(_w_10791));
  bfr _b_8889(.a(_w_10791),.q(_w_10792));
  bfr _b_14005(.a(_w_15907),.q(_w_15908));
  bfr _b_8890(.a(_w_10792),.q(_w_10793));
  bfr _b_9397(.a(_w_11299),.q(_w_11300));
  bfr _b_8891(.a(_w_10793),.q(_w_10794));
  bfr _b_8893(.a(_w_10795),.q(_w_10796));
  bfr _b_8977(.a(_w_10879),.q(n954));
  bfr _b_11323(.a(_w_13225),.q(_w_13226));
  bfr _b_8894(.a(_w_10796),.q(_w_10797));
  bfr _b_9912(.a(_w_11814),.q(n506));
  bfr _b_8897(.a(_w_10799),.q(_w_10800));
  bfr _b_8898(.a(_w_10800),.q(n1052));
  bfr _b_8900(.a(_w_10802),.q(_w_10803));
  bfr _b_11569(.a(_w_13471),.q(_w_13472));
  bfr _b_8905(.a(_w_10807),.q(_w_10808));
  bfr _b_8907(.a(_w_10809),.q(_w_10810));
  bfr _b_3475(.a(_w_5377),.q(_w_5378));
  bfr _b_8909(.a(_w_10811),.q(_w_10812));
  bfr _b_14281(.a(_w_16183),.q(_w_16184));
  bfr _b_8910(.a(_w_10812),.q(_w_10813));
  bfr _b_8911(.a(_w_10813),.q(_w_10814));
  bfr _b_13552(.a(_w_15454),.q(_w_15455));
  bfr _b_8912(.a(_w_10814),.q(_w_10815));
  bfr _b_8914(.a(_w_10816),.q(_w_10817));
  bfr _b_8915(.a(_w_10817),.q(n1822));
  spl2 g94_s_0(.a(n94),.q0(n94_0),.q1(_w_11837));
  spl2 g1814_s_0(.a(n1814),.q0(n1814_0),.q1(n1814_1));
  bfr _b_8916(.a(_w_10818),.q(n601));
  bfr _b_9143(.a(_w_11045),.q(_w_11046));
  bfr _b_8918(.a(_w_10820),.q(n1008));
  and_bb g1167(.a(N494_9),.b(N86_17),.q(_w_12930));
  bfr _b_8920(.a(_w_10822),.q(_w_10823));
  bfr _b_13783(.a(_w_15685),.q(_w_15686));
  bfr _b_8833(.a(_w_10735),.q(_w_10736));
  bfr _b_8924(.a(_w_10826),.q(_w_10827));
  bfr _b_8927(.a(_w_10829),.q(_w_10830));
  bfr _b_8928(.a(_w_10830),.q(_w_10831));
  bfr _b_12319(.a(_w_14221),.q(_w_14222));
  bfr _b_8929(.a(_w_10831),.q(_w_10832));
  bfr _b_8934(.a(_w_10836),.q(_w_10837));
  bfr _b_5480(.a(_w_7382),.q(_w_7383));
  bfr _b_8935(.a(_w_10837),.q(n728));
  bfr _b_7803(.a(_w_9705),.q(_w_9706));
  bfr _b_8939(.a(_w_10841),.q(_w_10842));
  bfr _b_8941(.a(_w_10843),.q(_w_10844));
  spl4L N35_s_1(.a(N35_0),.q0(N35_4),.q1(N35_5),.q2(_w_7259),.q3(_w_7261));
  bfr _b_10184(.a(_w_12086),.q(_w_12087));
  bfr _b_8943(.a(_w_10845),.q(_w_10846));
  bfr _b_12076(.a(_w_13978),.q(n791));
  bfr _b_6145(.a(_w_8047),.q(_w_8048));
  bfr _b_8949(.a(_w_10851),.q(_w_10852));
  bfr _b_8954(.a(_w_10856),.q(_w_10857));
  spl2 g1320_s_0(.a(n1320),.q0(n1320_0),.q1(n1320_1));
  bfr _b_8965(.a(_w_10867),.q(_w_10868));
  bfr _b_8966(.a(_w_10868),.q(_w_10869));
  bfr _b_8968(.a(_w_10870),.q(_w_10871));
  bfr _b_8969(.a(_w_10871),.q(_w_10872));
  bfr _b_13812(.a(_w_15714),.q(_w_15715));
  bfr _b_9739(.a(_w_11641),.q(_w_11642));
  bfr _b_11894(.a(_w_13796),.q(_w_13797));
  bfr _b_11365(.a(_w_13267),.q(_w_13268));
  bfr _b_8971(.a(_w_10873),.q(_w_10874));
  bfr _b_8972(.a(_w_10874),.q(_w_10875));
  bfr _b_4885(.a(_w_6787),.q(_w_6788));
  bfr _b_7711(.a(_w_9613),.q(_w_9614));
  bfr _b_8973(.a(_w_10875),.q(_w_10876));
  bfr _b_8975(.a(_w_10877),.q(_w_10878));
  bfr _b_8976(.a(_w_10878),.q(_w_10879));
  bfr _b_8978(.a(_w_10880),.q(n553));
  bfr _b_8981(.a(_w_10883),.q(n38));
  bfr _b_10092(.a(_w_11994),.q(_w_11995));
  bfr _b_8984(.a(_w_10886),.q(_w_10887));
  bfr _b_11631(.a(_w_13533),.q(_w_13534));
  bfr _b_4028(.a(_w_5930),.q(_w_5931));
  bfr _b_8985(.a(_w_10887),.q(_w_10888));
  bfr _b_8986(.a(_w_10888),.q(n1647_1));
  bfr _b_8988(.a(_w_10890),.q(_w_10891));
  bfr _b_8990(.a(_w_10892),.q(n700_1));
  bfr _b_8992(.a(_w_10894),.q(n461));
  bfr _b_8995(.a(_w_10897),.q(_w_10898));
  bfr _b_9297(.a(_w_11199),.q(_w_11200));
  bfr _b_8996(.a(_w_10898),.q(_w_10899));
  bfr _b_8999(.a(_w_10901),.q(_w_10902));
  bfr _b_8993(.a(_w_10895),.q(_w_10896));
  bfr _b_9000(.a(_w_10902),.q(_w_10903));
  or_bb g1021(.a(n1019_0),.b(n1020),.q(n1021));
  spl2 g956_s_0(.a(n956),.q0(n956_0),.q1(n956_1));
  bfr _b_6875(.a(_w_8777),.q(n131));
  bfr _b_9001(.a(_w_10903),.q(_w_10904));
  bfr _b_11759(.a(_w_13661),.q(_w_13662));
  bfr _b_9002(.a(_w_10904),.q(_w_10905));
  spl2 g430_s_0(.a(n430),.q0(n430_0),.q1(_w_13952));
  bfr _b_9003(.a(_w_10905),.q(_w_10906));
  bfr _b_9005(.a(_w_10907),.q(_w_10908));
  bfr _b_13156(.a(_w_15058),.q(_w_15059));
  bfr _b_9006(.a(_w_10908),.q(n452));
  bfr _b_13339(.a(_w_15241),.q(_w_15242));
  bfr _b_9008(.a(_w_10910),.q(_w_10911));
  spl4L N341_s_2(.a(N341_1),.q0(N341_8),.q1(N341_9),.q2(N341_10),.q3(N341_11));
  bfr _b_9009(.a(_w_10911),.q(_w_10912));
  bfr _b_9010(.a(_w_10912),.q(_w_10913));
  bfr _b_9011(.a(_w_10913),.q(n66_1));
  bfr _b_9014(.a(_w_10916),.q(_w_10917));
  spl2 g1167_s_0(.a(n1167),.q0(n1167_0),.q1(n1167_1));
  bfr _b_7534(.a(_w_9436),.q(_w_9437));
  bfr _b_9015(.a(_w_10917),.q(_w_10918));
  bfr _b_9017(.a(_w_10919),.q(_w_10920));
  bfr _b_9023(.a(_w_10925),.q(_w_10926));
  bfr _b_6023(.a(_w_7925),.q(_w_7926));
  bfr _b_9025(.a(_w_10927),.q(_w_10928));
  bfr _b_9027(.a(_w_10929),.q(_w_10930));
  bfr _b_13359(.a(_w_15261),.q(_w_15262));
  bfr _b_11115(.a(_w_13017),.q(_w_13018));
  bfr _b_10574(.a(_w_12476),.q(_w_12477));
  spl2 g105_s_0(.a(n105),.q0(n105_0),.q1(n105_1));
  spl2 g475_s_0(.a(n475),.q0(n475_0),.q1(n475_1));
  and_bi g733(.a(n646_1),.b(n649_1),.q(n733));
  and_bb g1328(.a(n1277_1),.b(n1326_1),.q(_w_9252));
  bfr _b_9029(.a(_w_10931),.q(_w_10932));
  bfr _b_9031(.a(_w_10933),.q(_w_10934));
  bfr _b_9037(.a(_w_10939),.q(_w_10940));
  and_bi g1611(.a(n1582_1),.b(n1585_1),.q(n1611));
  bfr _b_9039(.a(_w_10941),.q(_w_10942));
  and_bi g386(.a(n376_1),.b(n384_1),.q(_w_9959));
  bfr _b_9044(.a(_w_10946),.q(_w_10947));
  bfr _b_13057(.a(_w_14959),.q(n1771_1));
  bfr _b_9057(.a(_w_10959),.q(_w_10960));
  bfr _b_13913(.a(_w_15815),.q(_w_15816));
  spl2 g1529_s_0(.a(n1529),.q0(n1529_0),.q1(n1529_1));
  bfr _b_9058(.a(_w_10960),.q(_w_10961));
  and_bi g105(.a(n82_1),.b(n85_1),.q(n105));
  bfr _b_7084(.a(_w_8986),.q(_w_8987));
  bfr _b_9059(.a(_w_10961),.q(_w_10962));
  bfr _b_7610(.a(_w_9512),.q(_w_9513));
  bfr _b_9060(.a(_w_10962),.q(_w_10963));
  and_bb g1282(.a(N188_12),.b(N409_15),.q(n1282));
  bfr _b_9073(.a(_w_10975),.q(_w_10976));
  bfr _b_6824(.a(_w_8726),.q(n1237));
  bfr _b_9151(.a(_w_11053),.q(_w_11054));
  bfr _b_9075(.a(_w_10977),.q(_w_10978));
  bfr _b_9077(.a(_w_10979),.q(n1446_1));
  or_bb g1200(.a(n1182_0),.b(n1199_0),.q(n1200));
  bfr _b_9080(.a(_w_10982),.q(n389));
  bfr _b_9082(.a(_w_10984),.q(_w_10985));
  bfr _b_9085(.a(_w_10987),.q(_w_10988));
  bfr _b_9086(.a(_w_10988),.q(_w_10989));
  bfr _b_9088(.a(_w_10990),.q(_w_10991));
  bfr _b_9089(.a(_w_10991),.q(_w_10992));
  bfr _b_9091(.a(_w_10993),.q(_w_10994));
  bfr _b_9094(.a(_w_10996),.q(_w_10997));
  bfr _b_9099(.a(_w_11001),.q(_w_11002));
  bfr _b_3410(.a(_w_5312),.q(_w_5313));
  bfr _b_9100(.a(_w_11002),.q(_w_11003));
  bfr _b_3783(.a(_w_5685),.q(_w_5686));
  bfr _b_4054(.a(_w_5956),.q(_w_5957));
  spl2 g499_s_0(.a(n499),.q0(n499_0),.q1(n499_1));
  bfr _b_10131(.a(_w_12033),.q(n1399));
  and_bi g50(.a(n40_1),.b(n48_1),.q(_w_11576));
  bfr _b_9103(.a(_w_11005),.q(_w_11006));
  bfr _b_6899(.a(_w_8801),.q(_w_8802));
  bfr _b_5979(.a(_w_7881),.q(_w_7882));
  bfr _b_9857(.a(_w_11759),.q(_w_11760));
  bfr _b_9202(.a(_w_11104),.q(_w_11105));
  bfr _b_7953(.a(_w_9855),.q(_w_9856));
  bfr _b_9106(.a(_w_11008),.q(_w_11009));
  bfr _b_9107(.a(_w_11009),.q(_w_11010));
  bfr _b_6550(.a(_w_8452),.q(_w_8453));
  bfr _b_9110(.a(_w_11012),.q(_w_11013));
  and_bi g1767(.a(n1765_0),.b(n1766),.q(n1767));
  bfr _b_9111(.a(_w_11013),.q(_w_11014));
  spl2 g411_s_0(.a(n411),.q0(n411_0),.q1(n411_1));
  bfr _b_9114(.a(_w_11016),.q(n70));
  bfr _b_13756(.a(_w_15658),.q(_w_15659));
  bfr _b_4164(.a(_w_6066),.q(_w_6067));
  bfr _b_9127(.a(_w_11029),.q(_w_11030));
  bfr _b_9117(.a(_w_11019),.q(_w_11020));
  bfr _b_11399(.a(_w_13301),.q(_w_13302));
  bfr _b_9118(.a(_w_11020),.q(_w_11021));
  bfr _b_9119(.a(_w_11021),.q(n946));
  bfr _b_9122(.a(_w_11024),.q(n122));
  bfr _b_9125(.a(_w_11027),.q(n610));
  bfr _b_13814(.a(_w_15716),.q(_w_15717));
  bfr _b_7111(.a(_w_9013),.q(_w_9014));
  and_bi g1657(.a(n1610_1),.b(n1655_1),.q(_w_13984));
  bfr _b_9126(.a(_w_11028),.q(_w_11029));
  bfr _b_12135(.a(_w_14037),.q(N6220));
  bfr _b_9128(.a(_w_11030),.q(_w_11031));
  bfr _b_4078(.a(_w_5980),.q(_w_5981));
  bfr _b_9132(.a(_w_11034),.q(_w_11035));
  bfr _b_9134(.a(_w_11036),.q(_w_11037));
  bfr _b_8119(.a(_w_10021),.q(_w_10022));
  bfr _b_9135(.a(_w_11037),.q(_w_11038));
  bfr _b_6033(.a(_w_7935),.q(_w_7936));
  bfr _b_9136(.a(_w_11038),.q(_w_11039));
  bfr _b_6692(.a(_w_8594),.q(n938));
  bfr _b_9138(.a(_w_11040),.q(_w_11041));
  bfr _b_7743(.a(_w_9645),.q(_w_9646));
  bfr _b_9139(.a(_w_11041),.q(_w_11042));
  and_bi g598(.a(n524_1),.b(n596_1),.q(_w_9582));
  bfr _b_8516(.a(_w_10418),.q(_w_10419));
  bfr _b_9140(.a(_w_11042),.q(_w_11043));
  bfr _b_9141(.a(_w_11043),.q(_w_11044));
  bfr _b_12078(.a(_w_13980),.q(_w_13981));
  bfr _b_10117(.a(_w_12019),.q(_w_12020));
  bfr _b_9142(.a(_w_11044),.q(_w_11045));
  bfr _b_10218(.a(_w_12120),.q(_w_12121));
  bfr _b_9144(.a(_w_11046),.q(_w_11047));
  bfr _b_9146(.a(_w_11048),.q(_w_11049));
  bfr _b_11633(.a(_w_13535),.q(_w_13536));
  bfr _b_3759(.a(_w_5661),.q(_w_5662));
  bfr _b_9852(.a(_w_11754),.q(_w_11755));
  bfr _b_9149(.a(_w_11051),.q(n1535));
  bfr _b_9153(.a(_w_11055),.q(_w_11056));
  spl2 g889_s_0(.a(n889),.q0(n889_0),.q1(n889_1));
  bfr _b_9158(.a(_w_11060),.q(n125));
  bfr _b_9163(.a(_w_11065),.q(_w_11066));
  bfr _b_12526(.a(_w_14428),.q(_w_14429));
  bfr _b_9167(.a(_w_11069),.q(_w_11070));
  bfr _b_9168(.a(_w_11070),.q(_w_11071));
  bfr _b_14286(.a(_w_16188),.q(_w_16189));
  bfr _b_5705(.a(_w_7607),.q(N222_18));
  and_bi g1743(.a(n1741_0),.b(n1742),.q(n1743));
  bfr _b_10084(.a(_w_11986),.q(_w_11987));
  bfr _b_10213(.a(_w_12115),.q(_w_12116));
  bfr _b_9169(.a(_w_11071),.q(_w_11072));
  bfr _b_12415(.a(_w_14317),.q(_w_14318));
  spl2 g369_s_0(.a(n369),.q0(n369_0),.q1(n369_1));
  bfr _b_9171(.a(_w_11073),.q(_w_11074));
  spl2 g1549_s_0(.a(n1549),.q0(n1549_0),.q1(n1549_1));
  bfr _b_9173(.a(_w_11075),.q(_w_11076));
  bfr _b_9174(.a(_w_11076),.q(_w_11077));
  bfr _b_4010(.a(_w_5912),.q(N239_7));
  bfr _b_9314(.a(_w_11216),.q(_w_11217));
  bfr _b_9177(.a(_w_11079),.q(_w_11080));
  bfr _b_9182(.a(_w_11084),.q(_w_11085));
  bfr _b_11626(.a(_w_13528),.q(_w_13529));
  bfr _b_9187(.a(_w_11089),.q(_w_11090));
  bfr _b_5245(.a(_w_7147),.q(_w_7148));
  bfr _b_9192(.a(_w_11094),.q(_w_11095));
  bfr _b_9193(.a(_w_11095),.q(_w_11096));
  bfr _b_11268(.a(_w_13170),.q(_w_13171));
  or_bb g1083(.a(n1073_0),.b(n1082_0),.q(n1083));
  bfr _b_5258(.a(_w_7160),.q(_w_7161));
  bfr _b_8183(.a(_w_10085),.q(_w_10086));
  bfr _b_9195(.a(_w_11097),.q(_w_11098));
  bfr _b_9197(.a(_w_11099),.q(_w_11100));
  bfr _b_9200(.a(_w_11102),.q(_w_11103));
  bfr _b_7456(.a(_w_9358),.q(_w_9359));
  bfr _b_9201(.a(_w_11103),.q(_w_11104));
  bfr _b_7983(.a(_w_9885),.q(_w_9886));
  bfr _b_9208(.a(_w_11110),.q(_w_11111));
  bfr _b_9209(.a(_w_11111),.q(_w_11112));
  bfr _b_7458(.a(_w_9360),.q(_w_9361));
  bfr _b_9211(.a(_w_11113),.q(_w_11114));
  bfr _b_4238(.a(_w_6140),.q(_w_6141));
  bfr _b_9212(.a(_w_11114),.q(_w_11115));
  bfr _b_9414(.a(_w_11316),.q(_w_11317));
  bfr _b_9213(.a(_w_11115),.q(_w_11116));
  bfr _b_9222(.a(_w_11124),.q(_w_11125));
  bfr _b_10589(.a(_w_12491),.q(_w_12492));
  bfr _b_9224(.a(_w_11126),.q(_w_11127));
  bfr _b_13565(.a(_w_15467),.q(_w_15468));
  bfr _b_9225(.a(_w_11127),.q(_w_11128));
  bfr _b_9227(.a(_w_11129),.q(_w_11130));
  bfr _b_9228(.a(_w_11130),.q(_w_11131));
  bfr _b_4321(.a(_w_6223),.q(_w_6224));
  bfr _b_9230(.a(_w_11132),.q(n1610));
  bfr _b_9232(.a(_w_11134),.q(_w_11135));
  bfr _b_9234(.a(_w_11136),.q(_w_11137));
  bfr _b_10069(.a(_w_11971),.q(_w_11972));
  bfr _b_9235(.a(_w_11137),.q(_w_11138));
  bfr _b_9236(.a(_w_11138),.q(_w_11139));
  bfr _b_12674(.a(_w_14576),.q(_w_14577));
  bfr _b_9238(.a(_w_11140),.q(_w_11141));
  bfr _b_5244(.a(_w_7146),.q(_w_7147));
  bfr _b_5568(.a(_w_7470),.q(n382_1));
  bfr _b_9239(.a(_w_11141),.q(_w_11142));
  bfr _b_9242(.a(_w_11144),.q(_w_11145));
  bfr _b_9243(.a(_w_11145),.q(n944));
  spl2 g548_s_0(.a(n548),.q0(n548_0),.q1(n548_1));
  bfr _b_9244(.a(_w_11146),.q(_w_11147));
  bfr _b_10790(.a(_w_12692),.q(_w_12693));
  bfr _b_5274(.a(_w_7176),.q(_w_7177));
  bfr _b_5691(.a(_w_7593),.q(_w_7594));
  bfr _b_9247(.a(_w_11149),.q(_w_11150));
  bfr _b_9250(.a(_w_11152),.q(_w_11153));
  bfr _b_4857(.a(_w_6759),.q(_w_6760));
  bfr _b_7679(.a(_w_9581),.q(n558_1));
  bfr _b_9251(.a(_w_11153),.q(_w_11154));
  bfr _b_9252(.a(_w_11154),.q(_w_11155));
  bfr _b_9253(.a(_w_11155),.q(_w_11156));
  bfr _b_9261(.a(_w_11163),.q(_w_11164));
  bfr _b_9265(.a(_w_11167),.q(_w_11168));
  bfr _b_9266(.a(_w_11168),.q(_w_11169));
  spl2 g93_s_0(.a(n93),.q0(n93_0),.q1(n93_1));
  bfr _b_9270(.a(_w_11172),.q(_w_11173));
  bfr _b_9271(.a(_w_11173),.q(n822));
  bfr _b_9272(.a(_w_11174),.q(_w_11175));
  bfr _b_9277(.a(_w_11179),.q(_w_11180));
  spl2 g1309_s_0(.a(n1309),.q0(n1309_0),.q1(_w_15093));
  bfr _b_9279(.a(_w_11181),.q(_w_11182));
  bfr _b_14294(.a(_w_16196),.q(_w_16108));
  bfr _b_9283(.a(_w_11185),.q(_w_11186));
  bfr _b_9284(.a(_w_11186),.q(_w_11187));
  and_bb g1272(.a(N103_17),.b(N494_10),.q(_w_13079));
  bfr _b_9286(.a(_w_11188),.q(_w_11189));
  bfr _b_3687(.a(_w_5589),.q(_w_5590));
  and_bi g1413(.a(n1412_0),.b(n1375_0),.q(n1413));
  bfr _b_9288(.a(_w_11190),.q(_w_11191));
  bfr _b_7700(.a(_w_9602),.q(_w_9603));
  bfr _b_9205(.a(_w_11107),.q(n1408));
  bfr _b_9289(.a(_w_11191),.q(_w_11192));
  bfr _b_9291(.a(_w_11193),.q(_w_11194));
  bfr _b_9294(.a(_w_11196),.q(_w_11197));
  bfr _b_13477(.a(_w_15379),.q(_w_15380));
  bfr _b_9295(.a(_w_11197),.q(_w_11198));
  bfr _b_9296(.a(_w_11198),.q(_w_11199));
  bfr _b_8837(.a(_w_10739),.q(_w_10740));
  bfr _b_9299(.a(_w_11201),.q(_w_11202));
  bfr _b_9300(.a(_w_11202),.q(_w_11203));
  spl2 g709_s_0(.a(n709),.q0(n709_0),.q1(n709_1));
  bfr _b_9301(.a(_w_11203),.q(_w_11204));
  spl2 g804_s_0(.a(n804),.q0(n804_0),.q1(n804_1));
  bfr _b_9302(.a(_w_11204),.q(_w_11205));
  bfr _b_6825(.a(_w_8727),.q(n927));
  bfr _b_9672(.a(_w_11574),.q(_w_11575));
  bfr _b_9303(.a(_w_11205),.q(_w_11206));
  bfr _b_10914(.a(_w_12816),.q(_w_12817));
  bfr _b_5351(.a(_w_7253),.q(_w_7254));
  bfr _b_9528(.a(_w_11430),.q(_w_11431));
  bfr _b_7746(.a(_w_9648),.q(_w_9649));
  bfr _b_9304(.a(_w_11206),.q(_w_11207));
  bfr _b_12941(.a(_w_14843),.q(_w_14844));
  and_bi g178(.a(n136_1),.b(n176_1),.q(_w_12095));
  bfr _b_9306(.a(_w_11208),.q(_w_11209));
  spl2 g1617_s_0(.a(n1617),.q0(n1617_0),.q1(n1617_1));
  bfr _b_9307(.a(_w_11209),.q(_w_11210));
  bfr _b_9309(.a(_w_11211),.q(_w_11212));
  bfr _b_9974(.a(_w_11876),.q(_w_11877));
  bfr _b_9310(.a(_w_11212),.q(_w_11213));
  bfr _b_10933(.a(_w_12835),.q(_w_12836));
  bfr _b_10050(.a(_w_11952),.q(_w_11953));
  bfr _b_5741(.a(_w_7643),.q(_w_7644));
  bfr _b_9379(.a(_w_11281),.q(_w_11282));
  bfr _b_9313(.a(_w_11215),.q(_w_11216));
  bfr _b_9315(.a(_w_11217),.q(_w_11218));
  bfr _b_9320(.a(_w_11222),.q(_w_11223));
  bfr _b_9323(.a(_w_11225),.q(N6160));
  bfr _b_9326(.a(_w_11228),.q(_w_11229));
  bfr _b_9328(.a(_w_11230),.q(_w_11231));
  spl3L g456_s_0(.a(n456),.q0(n456_0),.q1(_w_7885),.q2(_w_7887));
  bfr _b_6586(.a(_w_8488),.q(_w_8489));
  bfr _b_6578(.a(_w_8480),.q(_w_8481));
  bfr _b_9329(.a(_w_11231),.q(_w_11232));
  bfr _b_9330(.a(_w_11232),.q(_w_11233));
  bfr _b_9331(.a(_w_11233),.q(_w_11234));
  bfr _b_9333(.a(_w_11235),.q(_w_11236));
  and_bi g1196(.a(n1194_0),.b(n1195),.q(n1196));
  bfr _b_9334(.a(_w_11236),.q(_w_11237));
  bfr _b_9335(.a(_w_11237),.q(_w_11238));
  bfr _b_9338(.a(_w_11240),.q(_w_11241));
  bfr _b_9848(.a(_w_11750),.q(_w_11751));
  bfr _b_9777(.a(_w_11679),.q(_w_11680));
  bfr _b_9342(.a(_w_11244),.q(_w_11245));
  bfr _b_13509(.a(_w_15411),.q(_w_15412));
  bfr _b_9345(.a(_w_11247),.q(_w_11248));
  bfr _b_9346(.a(_w_11248),.q(_w_11249));
  bfr _b_9352(.a(_w_11254),.q(_w_11255));
  bfr _b_10699(.a(_w_12601),.q(_w_12602));
  bfr _b_9354(.a(_w_11256),.q(_w_11257));
  bfr _b_10915(.a(_w_12817),.q(_w_12818));
  bfr _b_9357(.a(_w_11259),.q(_w_11260));
  bfr _b_9364(.a(_w_11266),.q(_w_11267));
  bfr _b_8138(.a(_w_10040),.q(_w_10041));
  bfr _b_9367(.a(_w_11269),.q(_w_11270));
  bfr _b_9369(.a(_w_11271),.q(_w_11272));
  bfr _b_9371(.a(_w_11273),.q(_w_11274));
  bfr _b_11488(.a(_w_13390),.q(_w_13391));
  bfr _b_9372(.a(_w_11274),.q(_w_11275));
  bfr _b_9374(.a(_w_11276),.q(_w_11277));
  and_bi g200(.a(n190_1),.b(n198_1),.q(_w_14290));
  bfr _b_9383(.a(_w_11285),.q(_w_11286));
  bfr _b_9385(.a(_w_11287),.q(_w_11288));
  bfr _b_6382(.a(_w_8284),.q(_w_8285));
  bfr _b_9387(.a(_w_11289),.q(_w_11290));
  bfr _b_9456(.a(_w_11358),.q(_w_11359));
  bfr _b_7237(.a(_w_9139),.q(n818));
  bfr _b_9389(.a(_w_11291),.q(_w_11292));
  bfr _b_9390(.a(_w_11292),.q(_w_11293));
  bfr _b_9392(.a(_w_11294),.q(_w_11295));
  bfr _b_12622(.a(_w_14524),.q(_w_14525));
  bfr _b_9394(.a(_w_11296),.q(_w_11297));
  bfr _b_9395(.a(_w_11297),.q(_w_11298));
  bfr _b_9396(.a(_w_11298),.q(_w_11299));
  bfr _b_12818(.a(_w_14720),.q(_w_14721));
  bfr _b_9575(.a(_w_11477),.q(_w_11478));
  bfr _b_9402(.a(_w_11304),.q(_w_11305));
  bfr _b_9403(.a(_w_11305),.q(_w_11306));
  bfr _b_13138(.a(_w_15040),.q(_w_15041));
  bfr _b_9406(.a(_w_11308),.q(_w_11309));
  bfr _b_9416(.a(_w_11318),.q(_w_11319));
  bfr _b_9418(.a(_w_11320),.q(_w_11321));
  bfr _b_9419(.a(_w_11321),.q(_w_11322));
  spl2 g40_s_0(.a(n40),.q0(n40_0),.q1(n40_1));
  bfr _b_9421(.a(_w_11323),.q(_w_11324));
  bfr _b_4749(.a(_w_6651),.q(_w_6652));
  bfr _b_5550(.a(_w_7452),.q(_w_7453));
  bfr _b_8491(.a(_w_10393),.q(_w_10394));
  bfr _b_9422(.a(_w_11324),.q(_w_11325));
  bfr _b_13548(.a(_w_15450),.q(_w_15451));
  bfr _b_8037(.a(_w_9939),.q(_w_9940));
  bfr _b_9423(.a(_w_11325),.q(_w_11326));
  bfr _b_9424(.a(_w_11326),.q(_w_11327));
  bfr _b_9425(.a(_w_11327),.q(_w_11328));
  bfr _b_9429(.a(_w_11331),.q(_w_11332));
  bfr _b_9431(.a(_w_11333),.q(_w_11334));
  bfr _b_9432(.a(_w_11334),.q(_w_11335));
  bfr _b_9435(.a(_w_11337),.q(_w_11338));
  bfr _b_9439(.a(_w_11341),.q(_w_11342));
  bfr _b_9440(.a(_w_11342),.q(_w_11343));
  bfr _b_9442(.a(_w_11344),.q(_w_11345));
  bfr _b_9547(.a(_w_11449),.q(_w_11450));
  bfr _b_9444(.a(_w_11346),.q(_w_11347));
  bfr _b_11209(.a(_w_13111),.q(_w_13112));
  bfr _b_9446(.a(_w_11348),.q(_w_11349));
  bfr _b_9447(.a(_w_11349),.q(_w_11350));
  bfr _b_9448(.a(_w_11350),.q(_w_11351));
  bfr _b_8701(.a(_w_10603),.q(_w_10604));
  bfr _b_9449(.a(_w_11351),.q(_w_11352));
  bfr _b_9450(.a(_w_11352),.q(_w_11353));
  or_bb g317(.a(n315_0),.b(n316),.q(n317));
  bfr _b_9453(.a(_w_11355),.q(_w_11356));
  bfr _b_9458(.a(_w_11360),.q(_w_11361));
  bfr _b_10874(.a(_w_12776),.q(_w_12777));
  bfr _b_4549(.a(_w_6451),.q(_w_6452));
  bfr _b_10087(.a(_w_11989),.q(_w_11990));
  bfr _b_9459(.a(_w_11361),.q(_w_11362));
  bfr _b_9460(.a(_w_11362),.q(_w_11363));
  and_bb g1610(.a(N154_18),.b(N511_13),.q(_w_11117));
  bfr _b_9461(.a(_w_11363),.q(_w_11364));
  bfr _b_10537(.a(_w_12439),.q(_w_12440));
  bfr _b_9465(.a(_w_11367),.q(_w_11368));
  bfr _b_12122(.a(_w_14024),.q(_w_14025));
  bfr _b_9466(.a(_w_11368),.q(_w_11369));
  bfr _b_9478(.a(_w_11380),.q(_w_11381));
  bfr _b_9467(.a(_w_11369),.q(_w_11370));
  bfr _b_9469(.a(_w_11371),.q(_w_11372));
  bfr _b_9470(.a(_w_11372),.q(_w_11373));
  spl2 g1809_s_0(.a(n1809),.q0(n1809_0),.q1(n1809_1));
  bfr _b_5783(.a(_w_7685),.q(_w_7686));
  bfr _b_7825(.a(_w_9727),.q(_w_9728));
  bfr _b_7961(.a(_w_9863),.q(_w_9864));
  bfr _b_9473(.a(_w_11375),.q(_w_11376));
  bfr _b_9474(.a(_w_11376),.q(_w_11377));
  bfr _b_9476(.a(_w_11378),.q(_w_11379));
  bfr _b_4278(.a(_w_6180),.q(n748_1));
  bfr _b_4810(.a(_w_6712),.q(_w_6713));
  bfr _b_5734(.a(_w_7636),.q(_w_7637));
  bfr _b_9477(.a(_w_11379),.q(_w_11380));
  bfr _b_9067(.a(_w_10969),.q(_w_10970));
  bfr _b_9481(.a(_w_11383),.q(_w_11384));
  bfr _b_10717(.a(_w_12619),.q(_w_12620));
  and_bb g444(.a(N392_8),.b(N69_11),.q(n444));
  bfr _b_9487(.a(_w_11389),.q(_w_11390));
  bfr _b_10214(.a(_w_12116),.q(_w_12117));
  bfr _b_9490(.a(_w_11392),.q(_w_11393));
  bfr _b_9780(.a(_w_11682),.q(_w_11683));
  bfr _b_9491(.a(_w_11393),.q(_w_11394));
  bfr _b_9497(.a(_w_11399),.q(n1398_1));
  and_bi g890(.a(n889_0),.b(n834_0),.q(n890));
  bfr _b_6140(.a(_w_8042),.q(_w_8043));
  bfr _b_9498(.a(_w_11400),.q(n1313));
  bfr _b_5872(.a(_w_7774),.q(_w_7775));
  spl2 g370_s_0(.a(n370),.q0(n370_0),.q1(n370_1));
  bfr _b_9499(.a(_w_11401),.q(_w_11402));
  bfr _b_9501(.a(_w_11403),.q(_w_11404));
  bfr _b_3538(.a(_w_5440),.q(_w_5441));
  bfr _b_9502(.a(_w_11404),.q(n1315_1));
  bfr _b_10716(.a(_w_12618),.q(_w_12619));
  bfr _b_9504(.a(_w_11406),.q(_w_11407));
  and_bi g525(.a(n502_1),.b(n505_1),.q(n525));
  bfr _b_9505(.a(_w_11407),.q(_w_11408));
  bfr _b_9510(.a(_w_11412),.q(_w_11413));
  spl2 g908_s_0(.a(n908),.q0(n908_0),.q1(n908_1));
  bfr _b_9514(.a(_w_11416),.q(_w_11417));
  bfr _b_13557(.a(_w_15459),.q(_w_15460));
  bfr _b_9515(.a(_w_11417),.q(_w_11418));
  bfr _b_4618(.a(_w_6520),.q(_w_6521));
  bfr _b_4025(.a(_w_5927),.q(_w_5928));
  bfr _b_10256(.a(_w_12158),.q(_w_12159));
  bfr _b_7835(.a(_w_9737),.q(n1813));
  bfr _b_9521(.a(_w_11423),.q(_w_11424));
  bfr _b_14193(.a(_w_16095),.q(_w_16096));
  bfr _b_9522(.a(_w_11424),.q(_w_11425));
  bfr _b_9523(.a(_w_11425),.q(_w_11426));
  or_bb g1698(.a(n1680_0),.b(n1697_0),.q(n1698));
  bfr _b_9525(.a(_w_11427),.q(_w_11428));
  bfr _b_9526(.a(_w_11428),.q(_w_11429));
  bfr _b_9530(.a(_w_11432),.q(_w_11433));
  bfr _b_10561(.a(_w_12463),.q(_w_12464));
  bfr _b_6855(.a(_w_8757),.q(_w_8758));
  bfr _b_9531(.a(_w_11433),.q(_w_11434));
  bfr _b_9533(.a(_w_11435),.q(_w_11436));
  and_bi g697(.a(n696_0),.b(n616_0),.q(n697));
  bfr _b_6629(.a(_w_8531),.q(_w_8532));
  bfr _b_9534(.a(_w_11436),.q(_w_11437));
  bfr _b_3802(.a(_w_5704),.q(_w_5705));
  bfr _b_9538(.a(_w_11440),.q(_w_11441));
  bfr _b_9539(.a(_w_11441),.q(_w_11442));
  bfr _b_14049(.a(_w_15951),.q(_w_15952));
  bfr _b_9541(.a(_w_11443),.q(_w_11444));
  bfr _b_9543(.a(_w_11445),.q(_w_11446));
  bfr _b_9544(.a(_w_11446),.q(_w_11447));
  bfr _b_9549(.a(_w_11451),.q(_w_11452));
  bfr _b_13459(.a(_w_15361),.q(_w_15362));
  bfr _b_6635(.a(_w_8537),.q(_w_8538));
  bfr _b_9550(.a(_w_11452),.q(_w_11453));
  spl2 g1686_s_0(.a(n1686),.q0(n1686_0),.q1(_w_6153));
  or_bb g341(.a(n339_0),.b(n340),.q(n341));
  bfr _b_9553(.a(_w_11455),.q(_w_11456));
  bfr _b_9977(.a(_w_11879),.q(_w_11880));
  bfr _b_7894(.a(_w_9796),.q(_w_9797));
  bfr _b_9555(.a(_w_11457),.q(_w_11458));
  bfr _b_12433(.a(_w_14335),.q(_w_14336));
  bfr _b_9556(.a(_w_11458),.q(_w_11459));
  bfr _b_5154(.a(_w_7056),.q(_w_7057));
  bfr _b_3504(.a(_w_5406),.q(_w_5407));
  bfr _b_9012(.a(_w_10914),.q(_w_10915));
  bfr _b_9558(.a(_w_11460),.q(_w_11461));
  bfr _b_13520(.a(_w_15422),.q(_w_15423));
  bfr _b_10201(.a(_w_12103),.q(_w_12104));
  bfr _b_9560(.a(_w_11462),.q(_w_11463));
  bfr _b_4002(.a(_w_5904),.q(_w_5905));
  bfr _b_9568(.a(_w_11470),.q(_w_11471));
  spl2 g103_s_0(.a(n103),.q0(n103_0),.q1(n103_1));
  bfr _b_9570(.a(_w_11472),.q(_w_11473));
  bfr _b_9214(.a(_w_11116),.q(n138));
  bfr _b_9571(.a(_w_11473),.q(_w_11474));
  bfr _b_11049(.a(_w_12951),.q(n304));
  spl4L N205_s_0(.a(_w_15532),.q0(N205_0),.q1(_w_8391),.q2(_w_8415),.q3(_w_8471));
  bfr _b_9572(.a(_w_11474),.q(_w_11475));
  bfr _b_9524(.a(_w_11426),.q(_w_11427));
  or_bb g167(.a(n165_0),.b(n166),.q(n167));
  bfr _b_9573(.a(_w_11475),.q(_w_11476));
  bfr _b_4446(.a(_w_6348),.q(_w_6349));
  bfr _b_4564(.a(_w_6466),.q(_w_6467));
  bfr _b_9578(.a(_w_11480),.q(_w_11481));
  bfr _b_9579(.a(_w_11481),.q(_w_11482));
  bfr _b_3731(.a(_w_5633),.q(_w_5634));
  bfr _b_9580(.a(_w_11482),.q(_w_11483));
  bfr _b_10064(.a(_w_11966),.q(_w_11967));
  bfr _b_9585(.a(_w_11487),.q(_w_11488));
  bfr _b_9586(.a(_w_11488),.q(_w_11489));
  bfr _b_9554(.a(_w_11456),.q(_w_11457));
  bfr _b_7869(.a(_w_9771),.q(_w_9772));
  bfr _b_9587(.a(_w_11489),.q(_w_11490));
  and_bi g1694(.a(n1692_0),.b(n1693),.q(n1694));
  bfr _b_9588(.a(_w_11490),.q(_w_11491));
  bfr _b_13754(.a(_w_15656),.q(_w_15657));
  bfr _b_9600(.a(_w_11502),.q(_w_11503));
  bfr _b_9602(.a(_w_11504),.q(_w_11505));
  bfr _b_9604(.a(_w_11506),.q(_w_11507));
  and_bi g361(.a(n354_1),.b(n357_1),.q(n361));
  bfr _b_9605(.a(_w_11507),.q(_w_11508));
  and_bi g1487(.a(n1485_0),.b(n1486),.q(n1487));
  bfr _b_9606(.a(_w_11508),.q(_w_11509));
  bfr _b_5873(.a(_w_7775),.q(_w_7776));
  bfr _b_9609(.a(_w_11511),.q(_w_11512));
  bfr _b_12051(.a(_w_13953),.q(_w_13954));
  bfr _b_9612(.a(_w_11514),.q(_w_11515));
  and_bi g674(.a(n624_1),.b(n672_1),.q(_w_9638));
  bfr _b_9613(.a(_w_11515),.q(_w_11516));
  bfr _b_10928(.a(_w_12830),.q(_w_12831));
  spl2 g1640_s_0(.a(n1640),.q0(n1640_0),.q1(n1640_1));
  bfr _b_9614(.a(_w_11516),.q(_w_11517));
  bfr _b_13256(.a(_w_15158),.q(_w_15159));
  or_bb g1658(.a(n1656_0),.b(n1657),.q(n1658));
  bfr _b_9616(.a(_w_11518),.q(_w_11519));
  and_bb g395(.a(n373_1),.b(n393_1),.q(_w_12059));
  bfr _b_9617(.a(_w_11519),.q(_w_11520));
  bfr _b_11758(.a(_w_13660),.q(_w_13661));
  and_bi g957(.a(n863_1),.b(n866_1),.q(n957));
  bfr _b_9619(.a(_w_11521),.q(_w_11522));
  bfr _b_9620(.a(_w_11522),.q(_w_11523));
  bfr _b_9624(.a(_w_11526),.q(_w_11527));
  and_bi g365(.a(n342_1),.b(n345_1),.q(n365));
  bfr _b_9627(.a(_w_11529),.q(_w_11530));
  bfr _b_9630(.a(_w_11532),.q(_w_11533));
  bfr _b_6823(.a(_w_8725),.q(n930));
  bfr _b_10122(.a(_w_12024),.q(_w_12025));
  bfr _b_9634(.a(_w_11536),.q(_w_11537));
  bfr _b_9636(.a(_w_11538),.q(_w_11539));
  bfr _b_9495(.a(_w_11397),.q(_w_11398));
  bfr _b_9640(.a(_w_11542),.q(_w_11543));
  bfr _b_13393(.a(_w_15295),.q(n331));
  bfr _b_9641(.a(_w_11543),.q(_w_11544));
  bfr _b_9603(.a(_w_11505),.q(_w_11506));
  bfr _b_9643(.a(_w_11545),.q(_w_11546));
  bfr _b_9645(.a(_w_11547),.q(_w_11548));
  bfr _b_9648(.a(_w_11550),.q(_w_11551));
  bfr _b_9649(.a(_w_11551),.q(_w_11552));
  bfr _b_8942(.a(_w_10844),.q(_w_10845));
  bfr _b_9650(.a(_w_11552),.q(_w_11553));
  bfr _b_9651(.a(_w_11553),.q(_w_11554));
  bfr _b_3560(.a(_w_5462),.q(_w_5463));
  bfr _b_9652(.a(_w_11554),.q(_w_11555));
  spl2 g81_s_0(.a(n81),.q0(n81_0),.q1(n81_1));
  bfr _b_9653(.a(_w_11555),.q(_w_11556));
  bfr _b_7214(.a(_w_9116),.q(_w_9117));
  bfr _b_9657(.a(_w_11559),.q(_w_11560));
  bfr _b_11774(.a(_w_13676),.q(_w_13677));
  and_bi g1667(.a(n1665_0),.b(n1666),.q(n1667));
  bfr _b_9953(.a(_w_11855),.q(_w_11856));
  bfr _b_9658(.a(_w_11560),.q(_w_11561));
  bfr _b_9659(.a(_w_11561),.q(_w_11562));
  bfr _b_9662(.a(_w_11564),.q(_w_11565));
  bfr _b_13685(.a(_w_15587),.q(_w_15588));
  bfr _b_9663(.a(_w_11565),.q(_w_11566));
  bfr _b_5429(.a(_w_7331),.q(_w_7332));
  bfr _b_9664(.a(_w_11566),.q(_w_11567));
  bfr _b_3595(.a(_w_5497),.q(_w_5498));
  or_bb g862(.a(n860_0),.b(n861),.q(n862));
  bfr _b_9668(.a(_w_11570),.q(_w_11571));
  bfr _b_9673(.a(_w_11575),.q(N1581));
  bfr _b_9674(.a(_w_11576),.q(n50));
  bfr _b_4540(.a(_w_6442),.q(_w_6443));
  bfr _b_9676(.a(_w_11578),.q(n1477));
  bfr _b_9677(.a(_w_11579),.q(n1513));
  bfr _b_11383(.a(_w_13285),.q(_w_13286));
  bfr _b_9678(.a(_w_11580),.q(n1559));
  bfr _b_9679(.a(_w_11581),.q(_w_11582));
  bfr _b_13289(.a(_w_15191),.q(_w_15192));
  bfr _b_9682(.a(_w_11584),.q(_w_11585));
  bfr _b_13580(.a(_w_15482),.q(_w_15483));
  bfr _b_4504(.a(_w_6406),.q(_w_6407));
  bfr _b_9692(.a(_w_11594),.q(_w_11595));
  bfr _b_9694(.a(_w_11596),.q(n1218_1));
  bfr _b_9698(.a(_w_11600),.q(n1035));
  bfr _b_7203(.a(_w_9105),.q(_w_9106));
  bfr _b_9700(.a(_w_11602),.q(_w_11603));
  bfr _b_9702(.a(_w_11604),.q(_w_11605));
  bfr _b_9703(.a(_w_11605),.q(n646_1));
  bfr _b_9704(.a(_w_11606),.q(n870));
  bfr _b_9705(.a(_w_11607),.q(_w_11608));
  bfr _b_9707(.a(_w_11609),.q(_w_11610));
  bfr _b_5515(.a(_w_7417),.q(_w_7418));
  bfr _b_9709(.a(_w_11611),.q(_w_11612));
  bfr _b_11546(.a(_w_13448),.q(_w_13449));
  bfr _b_9710(.a(_w_11612),.q(_w_11613));
  bfr _b_9711(.a(_w_11613),.q(_w_11614));
  spl2 g262_s_0(.a(n262),.q0(n262_0),.q1(_w_8560));
  bfr _b_9712(.a(_w_11614),.q(_w_11615));
  bfr _b_13583(.a(_w_15485),.q(_w_15486));
  bfr _b_10072(.a(_w_11974),.q(_w_11975));
  bfr _b_9715(.a(_w_11617),.q(_w_11618));
  bfr _b_10007(.a(_w_11909),.q(_w_11910));
  bfr _b_9725(.a(_w_11627),.q(n1845_1));
  bfr _b_9726(.a(_w_11628),.q(n1571));
  spl2 g1242_s_0(.a(n1242),.q0(n1242_0),.q1(_w_8224));
  bfr _b_4808(.a(_w_6710),.q(_w_6711));
  bfr _b_9732(.a(_w_11634),.q(_w_11635));
  bfr _b_11900(.a(_w_13802),.q(_w_13803));
  bfr _b_9733(.a(_w_11635),.q(_w_11636));
  spl2 g1270_s_0(.a(n1270),.q0(n1270_0),.q1(n1270_1));
  bfr _b_9734(.a(_w_11636),.q(n190));
  bfr _b_9735(.a(_w_11637),.q(_w_11638));
  and_bi g909(.a(n828_1),.b(n907_1),.q(_w_12839));
  bfr _b_9736(.a(_w_11638),.q(_w_11639));
  bfr _b_11941(.a(_w_13843),.q(_w_13844));
  bfr _b_9809(.a(_w_11711),.q(_w_11712));
  bfr _b_9740(.a(_w_11642),.q(_w_11643));
  bfr _b_9742(.a(_w_11644),.q(_w_11645));
  bfr _b_9745(.a(_w_11647),.q(_w_11648));
  bfr _b_10051(.a(_w_11953),.q(_w_11954));
  bfr _b_10452(.a(_w_12354),.q(n956));
  bfr _b_4225(.a(_w_6127),.q(_w_6128));
  bfr _b_9748(.a(_w_11650),.q(_w_11651));
  bfr _b_9749(.a(_w_11651),.q(_w_11652));
  bfr _b_9758(.a(_w_11660),.q(N171_1));
  bfr _b_8732(.a(_w_10634),.q(_w_10635));
  bfr _b_9760(.a(_w_11662),.q(_w_11663));
  bfr _b_9764(.a(_w_11666),.q(_w_11667));
  bfr _b_14148(.a(_w_16050),.q(_w_16051));
  bfr _b_7255(.a(_w_9157),.q(_w_9158));
  bfr _b_9765(.a(_w_11667),.q(_w_11668));
  bfr _b_6856(.a(_w_8758),.q(_w_8759));
  bfr _b_9773(.a(_w_11675),.q(_w_11676));
  bfr _b_9774(.a(_w_11676),.q(_w_11677));
  spl2 g539_s_0(.a(n539),.q0(n539_0),.q1(n539_1));
  and_bi g320(.a(n318_0),.b(n319),.q(n320));
  bfr _b_9779(.a(_w_11681),.q(_w_11682));
  bfr _b_9781(.a(_w_11683),.q(_w_11684));
  bfr _b_6241(.a(_w_8143),.q(_w_8144));
  bfr _b_9784(.a(_w_11686),.q(_w_11687));
  spl4L N18_s_2(.a(N18_1),.q0(N18_8),.q1(N18_9),.q2(N18_10),.q3(_w_12035));
  and_bi g1324(.a(n1323_0),.b(n1278_0),.q(n1324));
  bfr _b_9785(.a(_w_11687),.q(_w_11688));
  bfr _b_11697(.a(_w_13599),.q(_w_13600));
  bfr _b_9787(.a(_w_11689),.q(_w_11690));
  bfr _b_14238(.a(_w_16140),.q(_w_16141));
  bfr _b_9788(.a(_w_11690),.q(_w_11691));
  bfr _b_11282(.a(_w_13184),.q(_w_13185));
  bfr _b_9790(.a(_w_11692),.q(_w_11693));
  bfr _b_12976(.a(_w_14878),.q(_w_14879));
  bfr _b_9794(.a(_w_11696),.q(_w_11697));
  bfr _b_4985(.a(_w_6887),.q(_w_6888));
  bfr _b_9796(.a(_w_11698),.q(_w_11699));
  bfr _b_9801(.a(_w_11703),.q(_w_11704));
  bfr _b_9804(.a(_w_11706),.q(_w_11707));
  bfr _b_9805(.a(_w_11707),.q(_w_11708));
  bfr _b_8277(.a(_w_10179),.q(_w_10180));
  bfr _b_9806(.a(_w_11708),.q(_w_11709));
  bfr _b_9807(.a(_w_11709),.q(_w_11710));
  bfr _b_9812(.a(_w_11714),.q(_w_11715));
  and_bb g1255(.a(n1164_1),.b(n1253_1),.q(_w_13037));
  and_bi g1538(.a(n1509_1),.b(n1512_1),.q(n1538));
  bfr _b_9814(.a(_w_11716),.q(N171_2));
  bfr _b_9815(.a(_w_11717),.q(_w_11718));
  bfr _b_9817(.a(_w_11719),.q(_w_11720));
  bfr _b_5509(.a(_w_7411),.q(_w_7412));
  bfr _b_9820(.a(_w_11722),.q(_w_11723));
  bfr _b_8301(.a(_w_10203),.q(_w_10204));
  bfr _b_9822(.a(_w_11724),.q(_w_11725));
  bfr _b_4455(.a(_w_6357),.q(n1594_1));
  or_bb g886(.a(n884_0),.b(n885),.q(n886));
  bfr _b_9823(.a(_w_11725),.q(_w_11726));
  bfr _b_9824(.a(_w_11726),.q(_w_11727));
  bfr _b_9826(.a(_w_11728),.q(_w_11729));
  bfr _b_9829(.a(_w_11731),.q(_w_11732));
  bfr _b_12156(.a(_w_14058),.q(_w_14059));
  bfr _b_3477(.a(_w_5379),.q(_w_5380));
  and_bb g1046(.a(n1045_0),.b(n935_0),.q(n1046));
  bfr _b_9831(.a(_w_11733),.q(_w_11734));
  bfr _b_9264(.a(_w_11166),.q(_w_11167));
  bfr _b_9833(.a(_w_11735),.q(_w_11736));
  bfr _b_4347(.a(_w_6249),.q(_w_6250));
  bfr _b_9836(.a(_w_11738),.q(_w_11739));
  bfr _b_9837(.a(_w_11739),.q(_w_11740));
  bfr _b_9841(.a(_w_11743),.q(_w_11744));
  bfr _b_9843(.a(_w_11745),.q(_w_11746));
  bfr _b_8622(.a(_w_10524),.q(_w_10525));
  bfr _b_9845(.a(_w_11747),.q(_w_11748));
  bfr _b_9851(.a(_w_11753),.q(_w_11754));
  bfr _b_9856(.a(_w_11758),.q(_w_11759));
  bfr _b_9859(.a(_w_11761),.q(_w_11762));
  bfr _b_9864(.a(_w_11766),.q(_w_11767));
  bfr _b_9865(.a(_w_11767),.q(_w_11768));
  bfr _b_9866(.a(_w_11768),.q(_w_11769));
  bfr _b_9869(.a(_w_11771),.q(_w_11772));
  bfr _b_10197(.a(_w_12099),.q(_w_12100));
  bfr _b_5634(.a(_w_7536),.q(_w_7537));
  bfr _b_9655(.a(_w_11557),.q(_w_11558));
  bfr _b_9870(.a(_w_11772),.q(_w_11773));
  bfr _b_9872(.a(_w_11774),.q(_w_11775));
  bfr _b_9873(.a(_w_11775),.q(_w_11776));
  or_bb g968(.a(n961_0),.b(n967_0),.q(n968));
  bfr _b_9876(.a(_w_11778),.q(_w_11779));
  bfr _b_13025(.a(_w_14927),.q(_w_14928));
  bfr _b_6005(.a(_w_7907),.q(_w_7908));
  bfr _b_9883(.a(_w_11785),.q(_w_11786));
  and_bb g1346(.a(n1271_1),.b(n1344_1),.q(_w_13432));
  bfr _b_9884(.a(_w_11786),.q(_w_11787));
  bfr _b_9886(.a(_w_11788),.q(_w_11789));
  bfr _b_9887(.a(_w_11789),.q(_w_11790));
  and_bb g1699(.a(n1680_1),.b(n1697_1),.q(_w_12356));
  spl4L N273_s_4(.a(N273_3),.q0(N273_16),.q1(N273_17),.q2(N273_18),.q3(_w_12733));
  bfr _b_9888(.a(_w_11790),.q(_w_11791));
  bfr _b_9889(.a(_w_11791),.q(_w_11792));
  bfr _b_11777(.a(_w_13679),.q(_w_13680));
  bfr _b_8632(.a(_w_10534),.q(_w_10535));
  and_bi g1525(.a(n1454_1),.b(n1523_1),.q(_w_13885));
  bfr _b_8861(.a(_w_10763),.q(_w_10764));
  bfr _b_9890(.a(_w_11792),.q(_w_11793));
  bfr _b_9891(.a(_w_11793),.q(_w_11794));
  bfr _b_9893(.a(_w_11795),.q(_w_11796));
  bfr _b_6209(.a(_w_8111),.q(_w_8112));
  bfr _b_9898(.a(_w_11800),.q(_w_11801));
  bfr _b_9904(.a(_w_11806),.q(n1228));
  bfr _b_10979(.a(_w_12881),.q(_w_12882));
  bfr _b_5933(.a(_w_7835),.q(_w_7836));
  bfr _b_9905(.a(_w_11807),.q(_w_11808));
  bfr _b_9907(.a(_w_11809),.q(_w_11810));
  bfr _b_9908(.a(_w_11810),.q(_w_11811));
  bfr _b_4313(.a(_w_6215),.q(_w_6216));
  bfr _b_9909(.a(_w_11811),.q(_w_11812));
  bfr _b_6964(.a(_w_8866),.q(_w_8867));
  bfr _b_9916(.a(_w_11818),.q(_w_11819));
  bfr _b_11215(.a(_w_13117),.q(_w_13118));
  bfr _b_9917(.a(_w_11819),.q(_w_11820));
  bfr _b_9919(.a(_w_11821),.q(_w_11822));
  bfr _b_10076(.a(_w_11978),.q(_w_11979));
  bfr _b_7160(.a(_w_9062),.q(_w_9063));
  bfr _b_9920(.a(_w_11822),.q(_w_11823));
  bfr _b_3948(.a(_w_5850),.q(_w_5851));
  bfr _b_9924(.a(_w_11826),.q(_w_11827));
  bfr _b_8774(.a(_w_10676),.q(_w_10677));
  bfr _b_9927(.a(_w_11829),.q(_w_11830));
  bfr _b_9931(.a(_w_11833),.q(_w_11834));
  bfr _b_10649(.a(_w_12551),.q(_w_12552));
  bfr _b_9818(.a(_w_11720),.q(_w_11721));
  bfr _b_9932(.a(_w_11834),.q(_w_11835));
  bfr _b_3968(.a(_w_5870),.q(_w_5871));
  bfr _b_9937(.a(_w_11839),.q(_w_11840));
  bfr _b_13278(.a(_w_15180),.q(_w_15181));
  or_bb g179(.a(n177_0),.b(n178),.q(_w_10307));
  and_bb g1878(.a(N239_19),.b(N528_18),.q(_w_14737));
  bfr _b_9943(.a(_w_11845),.q(n576_1));
  bfr _b_9945(.a(_w_11847),.q(_w_11848));
  bfr _b_9946(.a(_w_11848),.q(_w_11849));
  bfr _b_9950(.a(_w_11852),.q(_w_11853));
  and_bi g1012(.a(n1010_0),.b(n1011),.q(n1012));
  bfr _b_6415(.a(_w_8317),.q(_w_8318));
  bfr _b_9951(.a(_w_11853),.q(_w_11854));
  bfr _b_9959(.a(_w_11861),.q(_w_11862));
  bfr _b_9511(.a(_w_11413),.q(_w_11414));
  bfr _b_9269(.a(_w_11171),.q(_w_11172));
  bfr _b_9978(.a(_w_11880),.q(_w_11881));
  bfr _b_9979(.a(_w_11881),.q(_w_11882));
  bfr _b_4545(.a(_w_6447),.q(_w_6448));
  bfr _b_9981(.a(_w_11883),.q(_w_11884));
  bfr _b_9983(.a(_w_11885),.q(_w_11886));
  bfr _b_6397(.a(_w_8299),.q(n1190));
  bfr _b_8036(.a(_w_9938),.q(_w_9939));
  bfr _b_9986(.a(_w_11888),.q(_w_11889));
  bfr _b_9992(.a(_w_11894),.q(_w_11895));
  bfr _b_6919(.a(_w_8821),.q(_w_8822));
  bfr _b_9993(.a(_w_11895),.q(_w_11896));
  bfr _b_10793(.a(_w_12695),.q(_w_12696));
  or_bb g46(.a(n35_1),.b(n45_0),.q(n46));
  bfr _b_9996(.a(_w_11898),.q(_w_11899));
  bfr _b_10002(.a(_w_11904),.q(_w_11905));
  bfr _b_10008(.a(_w_11910),.q(_w_11911));
  bfr _b_10009(.a(_w_11911),.q(_w_11912));
  spl4L N239_s_1(.a(N239_0),.q0(N239_4),.q1(N239_5),.q2(_w_5909),.q3(_w_5911));
  bfr _b_9381(.a(_w_11283),.q(_w_11284));
  bfr _b_10013(.a(_w_11915),.q(_w_11916));
  bfr _b_10014(.a(_w_11916),.q(_w_11917));
  bfr _b_13820(.a(_w_15722),.q(_w_15723));
  bfr _b_10015(.a(_w_11917),.q(_w_11918));
  bfr _b_10017(.a(_w_11919),.q(_w_11920));
  bfr _b_4691(.a(_w_6593),.q(_w_6594));
  bfr _b_7754(.a(_w_9656),.q(_w_9657));
  bfr _b_10019(.a(_w_11921),.q(_w_11922));
  bfr _b_13767(.a(_w_15669),.q(_w_15621));
  bfr _b_11482(.a(_w_13384),.q(_w_13385));
  bfr _b_3503(.a(_w_5405),.q(_w_5406));
  bfr _b_10023(.a(_w_11925),.q(_w_11926));
  spl2 g1855_s_0(.a(n1855),.q0(n1855_0),.q1(n1855_1));
  bfr _b_3565(.a(_w_5467),.q(_w_5468));
  bfr _b_10112(.a(_w_12014),.q(_w_12015));
  bfr _b_9828(.a(_w_11730),.q(_w_11731));
  spl2 g88_s_0(.a(n88),.q0(n88_0),.q1(_w_8785));
  bfr _b_10024(.a(_w_11926),.q(_w_11927));
  bfr _b_10026(.a(_w_11928),.q(_w_11929));
  bfr _b_10029(.a(_w_11931),.q(_w_11932));
  bfr _b_10030(.a(_w_11932),.q(_w_11933));
  and_bi g799(.a(n798_0),.b(n718_0),.q(n799));
  bfr _b_10032(.a(_w_11934),.q(_w_11935));
  bfr _b_10033(.a(_w_11935),.q(_w_11936));
  bfr _b_10035(.a(_w_11937),.q(_w_11938));
  bfr _b_4331(.a(_w_6233),.q(_w_6234));
  bfr _b_10037(.a(_w_11939),.q(_w_11940));
  bfr _b_13864(.a(_w_15766),.q(_w_15767));
  spl2 g1287_s_0(.a(n1287),.q0(n1287_0),.q1(n1287_1));
  bfr _b_10038(.a(_w_11940),.q(_w_11941));
  bfr _b_10044(.a(_w_11946),.q(_w_11947));
  bfr _b_11006(.a(_w_12908),.q(_w_12909));
  bfr _b_10045(.a(_w_11947),.q(_w_11948));
  bfr _b_10049(.a(_w_11951),.q(_w_11952));
  bfr _b_10052(.a(_w_11954),.q(_w_11955));
  bfr _b_10056(.a(_w_11958),.q(_w_11959));
  spl2 g445_s_0(.a(n445),.q0(n445_0),.q1(n445_1));
  spl2 g1629_s_0(.a(n1629),.q0(n1629_0),.q1(_w_13902));
  bfr _b_10062(.a(_w_11964),.q(_w_11965));
  bfr _b_10070(.a(_w_11972),.q(_w_11973));
  and_bb g626(.a(N120_10),.b(N375_11),.q(_w_9347));
  bfr _b_10073(.a(_w_11975),.q(_w_11976));
  bfr _b_10074(.a(_w_11976),.q(_w_11977));
  bfr _b_10236(.a(_w_12138),.q(_w_12139));
  or_bb g688(.a(n619_0),.b(n687_0),.q(n688));
  bfr _b_10077(.a(_w_11979),.q(_w_11980));
  bfr _b_3927(.a(_w_5829),.q(_w_5830));
  bfr _b_6351(.a(_w_8253),.q(_w_8254));
  bfr _b_10080(.a(_w_11982),.q(_w_11983));
  and_bi g908(.a(n907_0),.b(n828_0),.q(n908));
  bfr _b_5300(.a(_w_7202),.q(_w_7203));
  bfr _b_8688(.a(_w_10590),.q(_w_10591));
  bfr _b_10082(.a(_w_11984),.q(_w_11985));
  bfr _b_10083(.a(_w_11985),.q(_w_11986));
  bfr _b_10091(.a(_w_11993),.q(_w_11994));
  or_bb g1870(.a(n1852_0),.b(n1869_0),.q(n1870));
  bfr _b_10093(.a(_w_11995),.q(_w_11996));
  bfr _b_10094(.a(_w_11996),.q(_w_11997));
  bfr _b_10095(.a(_w_11997),.q(_w_11998));
  bfr _b_4277(.a(_w_6179),.q(_w_6180));
  or_bb g213(.a(n211_0),.b(n212),.q(n213));
  bfr _b_10098(.a(_w_12000),.q(_w_12001));
  bfr _b_4261(.a(_w_6163),.q(_w_6164));
  bfr _b_5667(.a(_w_7569),.q(_w_7570));
  bfr _b_10099(.a(_w_12001),.q(_w_12002));
  bfr _b_11259(.a(_w_13161),.q(_w_13162));
  bfr _b_10103(.a(_w_12005),.q(_w_12006));
  bfr _b_10108(.a(_w_12010),.q(N1901));
  bfr _b_10109(.a(_w_12011),.q(n1195));
  bfr _b_10110(.a(_w_12012),.q(_w_12013));
  bfr _b_10111(.a(_w_12013),.q(_w_12014));
  bfr _b_6631(.a(_w_8533),.q(_w_8534));
  bfr _b_10127(.a(_w_12029),.q(_w_12030));
  bfr _b_10128(.a(_w_12030),.q(n1351_1));
  bfr _b_10130(.a(_w_12032),.q(n1495));
  bfr _b_10133(.a(_w_12035),.q(_w_12036));
  bfr _b_10138(.a(_w_12040),.q(_w_12041));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  bfr _b_10144(.a(_w_12046),.q(_w_12047));
  bfr _b_6456(.a(_w_8358),.q(n1865));
  bfr _b_10145(.a(_w_12047),.q(_w_12048));
  bfr _b_10147(.a(_w_12049),.q(_w_12050));
  bfr _b_10148(.a(_w_12050),.q(_w_12051));
  bfr _b_5639(.a(_w_7541),.q(_w_7542));
  bfr _b_10150(.a(_w_12052),.q(_w_12053));
  bfr _b_3652(.a(_w_5554),.q(n923_1));
  bfr _b_10151(.a(_w_12053),.q(_w_12054));
  bfr _b_9623(.a(_w_11525),.q(_w_11526));
  bfr _b_10152(.a(_w_12054),.q(_w_12055));
  bfr _b_11982(.a(_w_13884),.q(n1074));
  bfr _b_10153(.a(_w_12055),.q(_w_12056));
  bfr _b_10155(.a(_w_12057),.q(_w_12058));
  spl2 g1812_s_0(.a(n1812),.q0(n1812_0),.q1(_w_13097));
  bfr _b_10156(.a(_w_12058),.q(N18_11));
  bfr _b_10157(.a(_w_12059),.q(n395));
  bfr _b_10160(.a(_w_12062),.q(_w_12063));
  spl2 g1784_s_0(.a(n1784),.q0(n1784_0),.q1(n1784_1));
  and_bi g1063(.a(n998_1),.b(n1001_1),.q(n1063));
  or_bb g1291(.a(n1289_0),.b(n1290_0),.q(n1291));
  bfr _b_10161(.a(_w_12063),.q(_w_12064));
  spl4L N290_s_3(.a(N290_2),.q0(N290_12),.q1(N290_13),.q2(N290_14),.q3(N290_15));
  bfr _b_10165(.a(_w_12067),.q(_w_12068));
  bfr _b_10167(.a(_w_12069),.q(_w_12070));
  bfr _b_11010(.a(_w_12912),.q(n1163));
  bfr _b_10168(.a(_w_12070),.q(_w_12071));
  bfr _b_9552(.a(_w_11454),.q(_w_11455));
  bfr _b_10169(.a(_w_12071),.q(_w_12072));
  bfr _b_10170(.a(_w_12072),.q(n54));
  bfr _b_14047(.a(_w_15949),.q(_w_15950));
  and_bb g993(.a(n953_1),.b(n991_1),.q(_w_10661));
  bfr _b_10171(.a(_w_12073),.q(n906));
  bfr _b_14378(.a(_w_16280),.q(_w_16281));
  bfr _b_10016(.a(_w_11918),.q(_w_11919));
  bfr _b_10172(.a(_w_12074),.q(n343));
  bfr _b_10123(.a(_w_12025),.q(n104));
  bfr _b_10175(.a(_w_12077),.q(n349));
  bfr _b_5618(.a(_w_7520),.q(_w_7521));
  bfr _b_10178(.a(_w_12080),.q(_w_12081));
  bfr _b_12243(.a(_w_14145),.q(_w_14146));
  and_bi g1467(.a(n1398_1),.b(n1401_1),.q(n1467));
  bfr _b_10179(.a(_w_12081),.q(_w_12082));
  and_bi g839(.a(n760_1),.b(n763_1),.q(n839));
  bfr _b_6502(.a(_w_8404),.q(_w_8405));
  bfr _b_10180(.a(_w_12082),.q(_w_12083));
  bfr _b_10182(.a(_w_12084),.q(_w_12085));
  bfr _b_10186(.a(_w_12088),.q(_w_12089));
  and_bi g1602(.a(n1600_0),.b(n1601),.q(n1602));
  bfr _b_7793(.a(_w_9695),.q(_w_9696));
  bfr _b_10188(.a(_w_12090),.q(_w_12091));
  bfr _b_10191(.a(_w_12093),.q(n1423));
  bfr _b_5952(.a(_w_7854),.q(_w_7855));
  bfr _b_10196(.a(_w_12098),.q(_w_12099));
  spl2 g1196_s_0(.a(n1196),.q0(n1196_0),.q1(n1196_1));
  bfr _b_10199(.a(_w_12101),.q(_w_12102));
  bfr _b_12141(.a(_w_14043),.q(_w_14044));
  and_bi g1395(.a(n1394_0),.b(n1381_0),.q(n1395));
  bfr _b_10202(.a(_w_12104),.q(_w_12105));
  bfr _b_13258(.a(_w_15160),.q(_w_15161));
  bfr _b_3674(.a(_w_5576),.q(_w_5577));
  bfr _b_10205(.a(_w_12107),.q(_w_12108));
  and_bb g1278(.a(N154_14),.b(N443_13),.q(_w_9222));
  bfr _b_7979(.a(_w_9881),.q(_w_9882));
  bfr _b_10209(.a(_w_12111),.q(_w_12112));
  bfr _b_6971(.a(_w_8873),.q(_w_8874));
  bfr _b_10212(.a(_w_12114),.q(_w_12115));
  bfr _b_10215(.a(_w_12117),.q(_w_12118));
  bfr _b_5039(.a(_w_6941),.q(_w_6942));
  bfr _b_4111(.a(_w_6013),.q(_w_6014));
  bfr _b_10217(.a(_w_12119),.q(_w_12120));
  bfr _b_12574(.a(_w_14476),.q(_w_14477));
  bfr _b_6221(.a(_w_8123),.q(_w_8124));
  bfr _b_7481(.a(_w_9383),.q(_w_9384));
  bfr _b_10220(.a(_w_12122),.q(_w_12123));
  and_bi g1751(.a(n1736_1),.b(n1749_1),.q(_w_11067));
  bfr _b_10224(.a(_w_12126),.q(_w_12127));
  bfr _b_5948(.a(_w_7850),.q(_w_7851));
  bfr _b_10226(.a(_w_12128),.q(_w_12129));
  bfr _b_5852(.a(_w_7754),.q(_w_7755));
  bfr _b_10232(.a(_w_12134),.q(_w_12135));
  bfr _b_10233(.a(_w_12135),.q(_w_12136));
  bfr _b_13033(.a(_w_14935),.q(_w_14936));
  bfr _b_10238(.a(_w_12140),.q(_w_12141));
  bfr _b_10239(.a(_w_12141),.q(_w_12142));
  bfr _b_10243(.a(_w_12145),.q(_w_12146));
  bfr _b_10247(.a(_w_12149),.q(_w_12150));
  bfr _b_10255(.a(_w_12157),.q(_w_12158));
  bfr _b_12542(.a(_w_14444),.q(_w_14445));
  bfr _b_7858(.a(_w_9760),.q(_w_9761));
  bfr _b_10259(.a(_w_12161),.q(_w_12162));
  bfr _b_3700(.a(_w_5602),.q(_w_5603));
  bfr _b_10261(.a(_w_12163),.q(_w_12164));
  bfr _b_10263(.a(_w_12165),.q(_w_12166));
  bfr _b_10265(.a(_w_12167),.q(_w_12168));
  bfr _b_10266(.a(_w_12168),.q(_w_12169));
  bfr _b_10267(.a(_w_12169),.q(_w_12170));
  bfr _b_10268(.a(_w_12170),.q(_w_12171));
  bfr _b_10269(.a(_w_12171),.q(_w_12172));
endmodule
