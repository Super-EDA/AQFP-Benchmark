module counter_128 (in_18_,in_1_,in_7_,in_109_,in_13_,in_106_,in_54_,in_118_,in_101_,in_3_,in_0_,in_113_,in_56_,in_30_,in_89_,in_35_,in_70_,in_38_,in_100_,in_105_,in_28_,in_10_,in_9_,in_78_,in_29_,in_60_,in_94_,in_108_,in_117_,in_103_,in_67_,in_44_,in_57_,in_76_,in_47_,in_20_,in_84_,in_17_,in_72_,in_116_,in_16_,in_120_,in_104_,in_64_,in_125_,in_58_,in_42_,in_40_,in_81_,in_115_,in_88_,in_24_,in_33_,in_123_,in_61_,in_79_,in_31_,in_36_,in_82_,in_111_,in_68_,in_2_,in_87_,in_74_,in_114_,in_53_,in_83_,in_86_,in_65_,in_102_,in_6_,in_75_,in_4_,in_93_,in_45_,in_90_,in_80_,in_73_,in_46_,in_25_,in_107_,in_37_,in_85_,in_49_,in_39_,in_63_,in_12_,in_112_,in_32_,in_119_,in_77_,in_34_,in_41_,in_122_,in_124_,in_48_,in_92_,in_15_,in_55_,in_50_,in_5_,in_127_,in_96_,in_22_,in_43_,in_52_,in_51_,in_21_,in_95_,in_59_,in_69_,in_121_,in_97_,in_11_,in_98_,in_126_,in_14_,in_91_,in_26_,in_99_,in_27_,in_71_,in_8_,in_23_,in_110_,in_62_,in_66_,in_19_,out_3_,out_2_,out_5_,out_1_,out_0_,out_7_,out_4_,out_6_);
  input in_18_,in_1_,in_7_,in_109_,in_13_,in_106_,in_54_,in_118_,in_101_,in_3_,in_0_,in_113_,in_56_,in_30_,in_89_,in_35_,in_70_,in_38_,in_100_,in_105_,in_28_,in_10_,in_9_,in_78_,in_29_,in_60_,in_94_,in_108_,in_117_,in_103_,in_67_,in_44_,in_57_,in_76_,in_47_,in_20_,in_84_,in_17_,in_72_,in_116_,in_16_,in_120_,in_104_,in_64_,in_125_,in_58_,in_42_,in_40_,in_81_,in_115_,in_88_,in_24_,in_33_,in_123_,in_61_,in_79_,in_31_,in_36_,in_82_,in_111_,in_68_,in_2_,in_87_,in_74_,in_114_,in_53_,in_83_,in_86_,in_65_,in_102_,in_6_,in_75_,in_4_,in_93_,in_45_,in_90_,in_80_,in_73_,in_46_,in_25_,in_107_,in_37_,in_85_,in_49_,in_39_,in_63_,in_12_,in_112_,in_32_,in_119_,in_77_,in_34_,in_41_,in_122_,in_124_,in_48_,in_92_,in_15_,in_55_,in_50_,in_5_,in_127_,in_96_,in_22_,in_43_,in_52_,in_51_,in_21_,in_95_,in_59_,in_69_,in_121_,in_97_,in_11_,in_98_,in_126_,in_14_,in_91_,in_26_,in_99_,in_27_,in_71_,in_8_,in_23_,in_110_,in_62_,in_66_,in_19_;
  output out_3_,out_2_,out_5_,out_1_,out_0_,out_7_,out_4_,out_6_;
  wire _w_1737,_w_1733,_w_1731,_w_1727,_w_1722,_w_1721,_w_1720,_w_1716,_w_1715,_w_1711,_w_1710,_w_1709,_w_1707,_w_1704,_w_1702,_w_1701,_w_1697,_w_1696,_w_1695,_w_1694,_w_1691,_w_1689,_w_1688,_w_1687,_w_1686,_w_1685,_w_1681,_w_1679,_w_1676,_w_1675,_w_1665,_w_1664,_w_1662,_w_1660,_w_1657,_w_1654,_w_1652,_w_1647,_w_1644,_w_1642,_w_1639,_w_1637,_w_1636,_w_1634,_w_1633,_w_1632,_w_1631,_w_1630,_w_1629,_w_1626,_w_1621,_w_1618,_w_1615,_w_1614,_w_1613,_w_1612,_w_1611,_w_1627,_w_1610,_w_1609,_w_1608,_w_1606,_w_1605,_w_1604,_w_1601,_w_1599,_w_1597,_w_1594,_w_1590,_w_1588,_w_1587,_w_1585,_w_1584,_w_1582,_w_1581,_w_1580,_w_1576,_w_1575,_w_1568,_w_1565,_w_1645,_w_1563,_w_1562,_w_1561,_w_1559,_w_1558,_w_1556,_w_1551,_w_1550,_w_1546,_w_1542,_w_1541,_w_1538,_w_1555,_w_1537,_w_1536,_w_1535,_w_1544,_w_1533,_w_1532,_w_1529,_w_1528,_w_1683,_w_1526,_w_1524,_w_1521,_w_1520,_w_1518,_w_1640,_w_1512,_w_1511,_w_1510,_w_1509,_w_1504,_w_1503,_w_1502,_w_1692,_w_1500,_w_1499,_w_1494,_w_1493,_w_1492,_w_1491,_w_1490,_w_1486,_w_1485,_w_1484,_w_1481,_w_1480,_w_1478,_w_1476,_w_1472,_w_1471,_w_1470,_w_1469,_w_1467,_w_1600,_w_1466,_w_1463,_w_1458,_w_1456,_w_1453,_w_1451,_w_1448,_w_1447,_w_1445,_w_1444,_w_1443,_w_1441,_w_1439,_w_1648,_w_1438,_w_1436,_w_1435,_w_1434,_w_1433,_w_1432,_w_1428,_w_1427,_w_1425,_w_1423,_w_1496,_w_1420,_w_1656,_w_1419,_w_1415,_w_1414,_w_1413,_w_1410,_w_1409,_w_1517,_w_1408,_w_1407,_w_1406,_w_1399,_w_1398,_w_1396,_w_1395,_w_1393,_w_1616,_w_1392,_w_1515,_w_1391,_w_1390,_w_1387,_w_1386,_w_1384,_w_1383,_w_1382,_w_1379,_w_1375,_w_1374,_w_1373,_w_1371,_w_1705,_w_1454,_w_1370,_w_1369,_w_1367,_w_1366,_w_1365,_w_1364,_w_1362,_w_1361,_w_1355,_w_1351,_w_1350,_w_1736,_w_1347,_w_1346,_w_1345,_w_1343,_w_1342,_w_1340,_w_1430,_w_1339,_w_1337,_w_1334,_w_1598,_w_1344,_w_1333,_w_1332,_w_1331,_w_1330,_w_1699,_w_1329,_w_1324,_w_1322,_w_1321,_w_1319,_w_1317,_w_1315,_w_1312,_w_1311,_w_1308,_w_1305,_w_1303,_w_1301,n525_1,_w_1666,n525_0,n415_1,n415_0,n215_5,n215_4,n215_2,n215_1,n215_0,n514_2,_w_1673,n514_1,n514_0,n510_2,n510_0,n398_4,n398_3,n398_2,n398_1,n398_0,n503_2,_w_1378,n503_1,n503_0,n349_5,n349_4,n349_2,_w_1641,n349_1,n422_1,n422_0,n143_4,n143_2,_w_1684,n143_0,n492_1,n482_1,n311_0,n267_0,n478_2,_w_1519,n478_1,n478_0,n367_2,n367_1,_w_1678,_w_1376,n516_1,n471_2,n471_1,n471_0,n467_1,n166_2,n166_1,n166_0,n496_2,n496_1,n452_1,n449_0,n443_1,n443_0,n440_2,_w_1482,n440_0,n146_2,n146_1,n146_0,n439_1,n234_3,_w_1452,n234_2,_w_1531,n234_0,n491_0,n441_4,n441_3,n441_2,n441_1,n441_0,n506_0,n436_1,n433_2,n433_1,n428_4,n428_2,n428_0,n426_3,n426_0,_w_1356,n491_2,n474_1,n474_0,n425_1,n412_2,n412_1,_w_1402,n409_2,n485_2,n426_1,n485_1,n395_3,n395_2,_w_1522,n395_1,_w_1653,n395_0,n391_2,n391_0,n513_2,n513_1,n218_1,_w_1623,n218_0,n444_3,n444_1,n385_2,n440_1,n385_1,n385_0,_w_1431,n177_2,_w_1651,n177_1,n509_0,n382_1,n237_0,_w_1442,n444_2,n379_2,n379_0,n345_1,n345_0,n364_1,n359_2,_w_1583,n359_1,n356_2,_w_1360,n356_1,n248_1,n248_0,n354_1,n354_0,n534,n525,_w_1553,n415,_w_1671,n300_0,n521,n292,_w_1564,_w_1380,n512,_w_1643,n510,n398,_w_1325,n507,n504,n271_3,n529_1,n503,n500,_w_1578,n349,n422,n143,_w_1358,n328_0,n494,n282_1,n492,n490,n400_1,n487,n532_0,n482,n311,n480,n479,_w_1514,n267,n516,n469,_w_1497,n468,n467,n243_2,n466,n476,n496,n163_0,n425_2,n475_1,n239_0,n453,n451,n449,n447,n440,n146,n281_2,n339_0,n361_1,n492_2,n438,n234,_w_1495,n441,n436,_w_1498,n435,n224_0,n486,_w_1505,n183_0,n183_3,n429,n236_1,n221_0,n428,_w_1596,n284_1,n474,n546,n346_2,n412,n306_0,n514,n409,_w_1507,n393_3,_w_1628,_w_1465,n405,_w_1335,n437,_w_1650,n404,n400,_w_1638,n399,n391,n155_1,n508,n387,_w_1506,n318,n386,n444,n385,_w_1706,n383,_w_1426,n177,n240_0,n311_1,n225_1,n308_3,n380,n379,_w_1714,n266,n237_1,n370,_w_1693,_w_1560,_w_1527,n366,n364,n186_4,n444_4,n138,_w_1700,n233_2,_w_1545,n360,n196_0,n434,n513_0,n488_0,n359,n207,n424,n541_2,n357,n356,n211_1,n355,n248,n222_0,_w_1738,n410,n352,n452_0,n351,n376,n348,n369,n343,n340,n356_3,n413,n339,n373_0,n420,n212,n335,n155_3,n274_2,n166,n289_1,n334,n192_0,n332,_w_1732,_w_1437,_w_1412,n148_0,n290_1,n331,n526,_w_1488,n330,n186,n471,n329,n152_0,n328,_w_1459,n519,n327,n325,n319,n457,n478,n358,n316,n257_2,n417,_w_1708,n315,n312,n159_0,n491,n310,n239,n308,_w_1659,n142,n293_1,n306,n199,n328_3,n341,n193_0,n301,n300,n299,n501,n192,_w_1304,n211,_w_1487,n297,_w_1310,n377_2,n458_2,n241,n267_1,n286,n427_0,_w_1416,n373_1,n285,n452,n244,n473,n371_2,n511,n237_2,n284,n234_1,n226,n317_2,n167,n155_0,n448,n446,n282,n277,n324,n281,n392_1,n278,n233,n276,_w_1477,n407,_w_1348,n467_0,n212_2,n313,n272,n269,_w_1677,_w_1353,n129_0,n421,n265,n317,n312_1,n277_1,n263,n489,n261,n523_1,n260,n259,n160_1,n215,n194_1,n258,n257,_w_1450,n253,_w_1513,n403,n370_1,n251,n530,n250,n178,n522,n154,n261_0,n359_0,n243,_w_1723,n302,n279,n182,_w_1674,n395_4,n291_2,n488,n136,_w_1543,n239_2,n322,n280,_w_1617,n433,_w_1462,n245,n130_2,n350_1,n516_0,n465,n206_2,_w_1682,n463,n212_4,_w_1421,n523,_w_1357,n240_2,n298,n354_2,n414,n345,n425_0,n275,_w_1646,n389,n293,n295,n221,n206,n305_0,n491_1,n425,n535_1,n348_1,_w_1489,n542_0,_w_1461,n307,n181,n305,n212_3,_w_1728,n137,n533,_w_1440,n475_0,_w_1622,n393,n402,n323,n428_3,_w_1540,_w_1309,n177_0,n372,n209_2,_w_1483,n270,n439,n339_1,n213,n230_1,n344_2,_w_1719,n285_0,n224,n367_0,n326_1,_w_1501,n294_3,n367,n320_2,n397_1,n370_0,n377_0,n147,n361,n371,n218,n294,n406_0,_w_1655,n365,_w_1349,n153_1,_w_1607,n442,n289_0,n197,n535,n174,n344,n195,n515,n532_1,n255,n374,n482_0,n265_0,n139,n291_0,n211_0,n288,n158,n344_4,_w_1328,n240,_w_1318,_w_1554,n246,n450,n431_3,n317_1,n209,_w_1460,n336,n325_0,_w_1475,_w_1417,n458_1,n377_1,_w_1530,n352_0,_w_1567,n527,n231,n240_1,n325_2,n168,n430,n326,n204,n283,n172,n373,n520,n208_0,n205,n131_1,n382,n254,n216_0,_w_1635,n296,n423,n407_3,n303,n313_1,n460,n257_0,n186_3,n355_1,n176,n528,n337,_w_1359,n149,n199_1,n381,_w_1372,n379_1,n406,n517_2,n537,_w_1341,n273,n307_0,n461,n548,n135,n542,n440_3,n403_1,n182_1,n290,n133,n163,n554,n150,n342,n162_0,n347,_w_1602,n173_1,n475,n427,_w_1658,n431_4,n257_1,n446_2,n232,n262_1,n256,n449_1,n185_1,n194_0,n535_0,n188,n400_0,n200,n222,_w_1620,n138_1,n549,_w_1516,n452_2,_w_1549,n274,n541_1,n350_3,n446_1,n181_1,n520_1,n288_0,n179,n485_0,n304,n543_0,_w_1570,n529,n141,n196,n132,n481_0,n317_0,_w_1300,n297_0,n130,_w_1690,n395,n368_0,n493,n502_0,n394,n169_2,n175,_w_1566,n131,n444_0,n271,n172_0,n240_3,n300_4,_w_1338,n140,n144,n443_2,n346_0,n265_1,n194,n517,n145,_w_1552,n410_2,_w_1403,n419,n350,n411,n143_3,_w_1591,_w_1508,n382_0,n202,n137_2,n148,n186_2,n384,n151,n280_0,n455,n268,n407_2,_w_1397,n152,n153,n236,_w_1539,n162_1,n374_2,n309,n156,n188_1,n157,n136_1,n184,n396,_w_1385,n193,n159,n179_1,_w_1326,n443,n185,n495,n160,n161,n162,n392,n165,n531,n169,_w_1302,n206_0,_w_1313,n354,n171,n312_0,_w_1525,n210,n524_0,n155,n180,n183,n377,n187,n320,n390,_w_1405,n481_1,n189,n419_1,n190,_w_1577,n228,n524,n513,n342_0,_w_1314,n191,n242,_w_1725,n432,n203,n477,n353,n217,n219,n506,n220,n225,n496_0,n299_0,n375,_w_1574,n416_3,_w_1523,n230,n215_3,n433_0,n235,n454,n198,n553,n362,n505,n368_1,n273_0,_w_1548,n409_1,n287_1,_w_1474,n536,_w_1668,n206_4,n539,n388_1,_w_1457,n368,n541,n543,n545,n547,_w_1388,n551,n552,_w_1336,n171_1,n555,n543_1,n543_2,_w_1735,n541_0,n498,n230_0,n203_0,n458_0,n142_1,n227_0,n227_1,n174_1,_w_1547,_w_1381,n293_0,n334_0,n176_1,n227_2,n225_0,n233_0,n337_4,_w_1698,n225_2,n151_1,n219_0,n143_1,n219_1,n268_2,n219_2,n394_0,n528_1,n203_2,n203_3,n242_0,_w_1717,n242_1,n191_0,n191_1,n431,n330_0,n209_1,n331_2,n524_1,n175_1,n524_2,n249,n321,n189_0,_w_1667,_w_1422,n282_0,n283_0,n189_1,_w_1739,n149_1,_w_1718,n189_2,_w_1411,n502_1,n183_1,n183_2,n247,n320_1,n523_0,n180_1,n180_0,n328_2,n439_0,n180_2,n455_1,n171_0,n216_1,n532,n169_0,n407_0,_w_1669,n169_1,n229,n169_3,n302_0,_w_1624,n165_0,_w_1670,n165_1,_w_1449,n287,n392_0,n436_0,n400_2,n277_0,n392_2,n294_1,n392_3,n160_0,_w_1680,n160_2,n227,n160_3,n306_1,n495_1,n344_1,_w_1730,n185_0,n324_2,n193_1,n201,n287_0,_w_1569,n458,n193_2,n157_0,n199_0,n374_3,n349_3,n157_1,n427_1,n314_1,n157_2,_w_1661,_w_1429,n349_0,n192_1,n330_1,_w_1595,n156_0,n177_3,n374_0,n236_0,n156_1,n155_2,n153_0,n455_0,n333_0,n333_1,n259_0,n151_0,n412_0,n363,n151_2,n346_5,n532_2,n243_0,n148_1,_w_1713,_w_1368,n150_2,n202_0,n394_1,_w_1424,n356_0,n294_4,n516_2,n208,n296_0,_w_1571,n202_1,n509_1,n350_0,_w_1377,n350_2,n419_0,_w_1464,n169_4,n145_0,n145_1,n263_1,n319_1,n129,n517_0,n140_0,n142_0,_w_1400,n140_2,n134_0,n134_1,n280_1,n262,n393_0,n134_3,n173,n131_0,n406_1,n131_2,n175_0,n462,n431_0,n431_1,n407_4,n431_2,n394_2,_w_1592,n394_3,n325_1,n310_1,n130_0,n129_1,_w_1649,n456,n502,n132_0,n132_1,n251_0,_w_1307,n264_0,n196_1,n179_0,n291,n368_2,n368_3,_w_1663,n297_2,n274_0,n427_2,n274_1,n410_4,n274_4,n222_2,n553_0,n200_0,n200_1,n200_2,n427_3,_w_1603,n475_2,n342_1,n222_3,n150_0,n150_1,n163_1,n163_2,n252,n212_1,n482_2,n163_3,n163_4,_w_1394,n203_1,n133_0,n133_1,n290_0,n439_2,n340_1,n497,n542_1,n397_2,n265_3,n214,n542_2,n338,n461_0,n206_1,n378,n461_1,n320_0,n237,n149_0,n337_0,_w_1354,n337_1,n337_2,n337_3,n176_0,n303_0,n303_1,_w_1401,n254_0,n254_1,_w_1323,n416,n528_0,n388,n214_0,n152_1,n376_0,n214_1,n205_0,n525_2,n484,n205_1,n333,n520_0,n134,n201_0,n373_2,n428_1,n518,n172_1,n509,n296_1,n499,n388_0,_w_1404,n326_0,_w_1455,n245_1,n553_1,n409_0,n430_0,n206_3,n327_0,n314,n430_2,_w_1363,n168_0,n364_0,n282_2,n194_2,n445,n324_1,n139_1,n336_0,n336_1,n517_1,n291_1,n355_2,n201_1,n291_3,n158_0,n317_3,n499_1,n346_4,n158_1,n304_2,n297_1,n430_1,n139_0,_w_1619,n374_1,n515_0,n238,n515_1,n311_2,n547_1,n134_2,n515_2,_w_1726,n197_2,_w_1389,n195_0,n344_0,n344_3,n174_0,n170,n174_2,_w_1418,n197_0,n197_1,n197_3,n499_0,_w_1573,n294_0,_w_1712,n294_2,n159_1,n371_0,n186_1,n371_1,n361_0,n419_2,n140_3,n361_2,n173_2,n459,n271_0,n271_1,_w_1703,n224_1,n270_0,n410_1,n270_1,_w_1306,n208_1,n271_2,n323_0,_w_1589,n393_1,n328_1,n418,n340_2,n393_2,n416_0,n168_1,n416_1,n188_0,n137_0,n529_0,n305_1,_w_1479,n305_2,n288_2,n307_1,n506_1,n426_2,n483,n221_1,n221_2,n376_1,n523_2,n346,n245_2,n481,n136_0,n279_0,n216_2,n216_3,n488_1,n485,n300_3,n182_0,n406_2,n407_1,n209_0,n279_1,n260_1,n302_1,n472,n313_0,n274_3,n243_1,n137_1,n251_1,n251_2,n492_0,n264,n403_0,n239_1,_w_1625,n140_1,n259_1,n260_0,n316_1,_w_1327,n261_2,n130_1,n262_2,_w_1586,n263_0,n276_0,_w_1468,n317_4,_w_1724,n323_1,n346_1,n397,n289,n416_2,n264_1,n173_0,n265_2,n269_0,n304_0,n269_1,_w_1320,n510_1,n273_1,n276_1,n391_1,n261_1,n281_0,n281_1,_w_1572,n277_2,n334_1,n426,n268_0,_w_1534,n547_0,n288_1,_w_1729,n268_1,_w_1593,n283_1,n223,n499_2,n314_2,n284_0,n285_1,n355_0,n285_2,n285_3,n446_0,n506_2,n408,n299_1,n300_1,n300_2,_w_1473,n304_1,_w_1672,n245_0,n308_0,n308_1,n308_2,n310_0,n216,n314_0,_w_1557,n314_3,n401,n316_0,n358_0,n358_1,n529_2,_w_1579,n319_0,n322_0,n322_1,n397_0,_w_1316,n164,n327_1,n186_0,n233_1,n331_0,n331_1,n332_0,_w_1446,n195_1,n332_1,n495_0,n334_2,n324_0,n334_3,n340_0,n410_0,n262_0,n212_0,n222_1,n181_0,n346_3,n138_0,n348_0,_w_1734,_w_1352,n352_1,n410_3;

  bfr _b_1183(.a(_w_1739),.q(n374_1));
  bfr _b_1179(.a(_w_1735),.q(_w_1736));
  bfr _b_1178(.a(_w_1734),.q(_w_1735));
  bfr _b_1177(.a(_w_1733),.q(_w_1734));
  bfr _b_1176(.a(_w_1732),.q(n240_1));
  bfr _b_1175(.a(_w_1731),.q(_w_1732));
  bfr _b_1174(.a(_w_1730),.q(_w_1731));
  bfr _b_1173(.a(_w_1729),.q(n215_1));
  bfr _b_1171(.a(_w_1727),.q(n325_2));
  bfr _b_1170(.a(_w_1726),.q(_w_1727));
  bfr _b_1169(.a(_w_1725),.q(n140_1));
  bfr _b_1168(.a(_w_1724),.q(_w_1725));
  bfr _b_1166(.a(_w_1722),.q(n266));
  bfr _b_1164(.a(_w_1720),.q(n368_1));
  bfr _b_1163(.a(_w_1719),.q(_w_1720));
  bfr _b_1162(.a(_w_1718),.q(_w_1719));
  bfr _b_1161(.a(_w_1717),.q(n222_1));
  bfr _b_1159(.a(_w_1715),.q(_w_1716));
  bfr _b_1158(.a(_w_1714),.q(n394_1));
  bfr _b_1157(.a(_w_1713),.q(_w_1714));
  bfr _b_1156(.a(_w_1712),.q(n134_1));
  bfr _b_1154(.a(_w_1710),.q(_w_1711));
  bfr _b_1153(.a(_w_1709),.q(n517_2));
  bfr _b_1152(.a(_w_1708),.q(_w_1709));
  bfr _b_1148(.a(_w_1704),.q(_w_1705));
  bfr _b_1147(.a(_w_1703),.q(_w_1704));
  bfr _b_1146(.a(_w_1702),.q(n151_2));
  bfr _b_1144(.a(_w_1700),.q(n130));
  bfr _b_1141(.a(_w_1697),.q(_w_1698));
  bfr _b_1140(.a(_w_1696),.q(n155_3));
  bfr _b_1138(.a(_w_1694),.q(_w_1695));
  bfr _b_1137(.a(_w_1693),.q(n160_3));
  bfr _b_1136(.a(_w_1692),.q(n392_1));
  bfr _b_1135(.a(_w_1691),.q(_w_1692));
  bfr _b_1133(.a(_w_1689),.q(n180_2));
  bfr _b_1131(.a(_w_1687),.q(n183_1));
  bfr _b_1129(.a(_w_1685),.q(_w_1686));
  bfr _b_1128(.a(_w_1684),.q(n328_1));
  bfr _b_1127(.a(_w_1683),.q(_w_1684));
  bfr _b_1126(.a(_w_1682),.q(_w_1683));
  bfr _b_1125(.a(_w_1681),.q(n524_2));
  bfr _b_1124(.a(_w_1680),.q(_w_1681));
  bfr _b_1160(.a(_w_1716),.q(_w_1717));
  bfr _b_1122(.a(_w_1678),.q(n427_1));
  bfr _b_1120(.a(_w_1676),.q(n203_3));
  bfr _b_1119(.a(_w_1675),.q(n428_4));
  bfr _b_1118(.a(_w_1674),.q(_w_1675));
  bfr _b_1116(.a(_w_1672),.q(n398_4));
  bfr _b_1114(.a(_w_1670),.q(_w_1671));
  bfr _b_1113(.a(_w_1669),.q(n337_4));
  bfr _b_1111(.a(_w_1667),.q(_w_1668));
  bfr _b_1110(.a(_w_1666),.q(_w_1667));
  or_bb g537(.a(n514_1),.b(n535_1),.q(n537));
  or_bb g150(.a(in_108_),.b(in_109_),.q(_w_1733));
  spl2 g240_s_0(.a(n240),.q0(n240_0),.q1(_w_1730));
  spl2 g215_s_0(.a(n215),.q0(n215_0),.q1(_w_1729));
  spl2 g291_s_1(.a(n291_1),.q0(n291_2),.q1(_w_1728));
  spl2 g336_s_0(.a(n336),.q0(n336_0),.q1(n336_1));
  bfr _b_813(.a(_w_1369),.q(_w_1370));
  and_bb g325(.a(in_58_),.b(in_59_),.q(n325));
  and_bb g349(.a(n259_0),.b(n348_0),.q(n349));
  spl2 g310_s_0(.a(n310),.q0(n310_0),.q1(n310_1));
  spl2 g388_s_0(.a(n388),.q0(n388_0),.q1(n388_1));
  spl2 g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(_w_1723));
  spl2 g201_s_0(.a(n201),.q0(n201_0),.q1(n201_1));
  spl2 g520_s_0(.a(n520),.q0(n520_0),.q1(n520_1));
  spl2 g528_s_0(.a(n528),.q0(n528_0),.q1(n528_1));
  and_bb g252(.a(n233_0),.b(n251_0),.q(n252));
  spl2 g303_s_0(.a(n303),.q0(n303_0),.q1(n303_1));
  bfr _b_1121(.a(_w_1677),.q(_w_1678));
  spl2 g176_s_0(.a(n176),.q0(n176_0),.q1(n176_1));
  bfr _b_1085(.a(_w_1641),.q(n177_3));
  spl2 g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1));
  bfr _b_1151(.a(_w_1707),.q(_w_1708));
  bfr _b_1139(.a(_w_1695),.q(n157_2));
  and_bb g219(.a(n146_1),.b(n218_0),.q(n219));
  and_bb g307(.a(in_34_),.b(in_35_),.q(n307));
  bfr _b_1063(.a(_w_1619),.q(n378));
  spl3L g406_s_0(.a(n406),.q0(n406_0),.q1(n406_1),.q2(n406_2));
  maj_bbb g317(.a(n304_0),.b(n310_0),.c(n316_0),.q(n317));
  spl2 g273_s_0(.a(n273),.q0(n273_0),.q1(n273_1));
  bfr _b_824(.a(_w_1380),.q(_w_1381));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  maj_bbi g188(.a(n173_2),.b(n187),.c(n186_0),.q(n188));
  spl2 g222_s_1(.a(n222_1),.q0(n222_2),.q1(n222_3));
  bfr _b_918(.a(_w_1474),.q(n215_3));
  spl3L g209_s_0(.a(n209),.q0(n209_0),.q1(n209_1),.q2(n209_2));
  bfr _b_974(.a(_w_1530),.q(n192));
  spl2 g368_s_0(.a(n368),.q0(n368_0),.q1(_w_1718));
  bfr _b_1084(.a(_w_1640),.q(n543_2));
  spl2 g502_s_0(.a(n502),.q0(n502_0),.q1(n502_1));
  spl2 g394_s_1(.a(n394_1),.q0(n394_2),.q1(n394_3));
  spl3L g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1),.q2(n361_2));
  spl2 g158_s_0(.a(n158),.q0(n158_0),.q1(n158_1));
  spl2 g394_s_0(.a(n394),.q0(n394_0),.q1(_w_1713));
  spl2 g134_s_0(.a(n134),.q0(n134_0),.q1(_w_1710));
  or_bb g466(.a(n257_2),.b(n391_2),.q(n466));
  spl2 g145_s_0(.a(n145),.q0(n145_0),.q1(n145_1));
  spl2 g346_s_0(.a(n346),.q0(n346_0),.q1(_w_1706));
  spl2 g350_s_1(.a(n350_1),.q0(n350_2),.q1(n350_3));
  or_bb g130(.a(in_124_),.b(in_125_),.q(_w_1697));
  bfr _b_967(.a(_w_1523),.q(_w_1524));
  bfr _b_855(.a(_w_1411),.q(n431_4));
  spl2 g175_s_0(.a(n175),.q0(n175_0),.q1(n175_1));
  spl2 g495_s_0(.a(n495),.q0(n495_0),.q1(n495_1));
  maj_bbi g273(.a(n268_2),.b(n272),.c(n271_0),.q(n273));
  spl2 g392_s_0(.a(n392),.q0(n392_0),.q1(_w_1691));
  bfr _b_833(.a(_w_1389),.q(n206_4));
  bfr _b_1167(.a(_w_1723),.q(_w_1724));
  spl3L g180_s_0(.a(n180),.q0(n180_0),.q1(n180_1),.q2(_w_1688));
  spl2 g328_s_0(.a(n328),.q0(n328_0),.q1(_w_1682));
  bfr _b_1037(.a(_w_1593),.q(_w_1594));
  spl3L g524_s_0(.a(n524),.q0(n524_0),.q1(n524_1),.q2(_w_1679));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  and_bi g367(.a(n366),.b(n365),.q(n367));
  spl2 g427_s_0(.a(n427),.q0(n427_0),.q1(_w_1677));
  spl2 g346_s_2(.a(n346_3),.q0(n346_4),.q1(n346_5));
  spl2 g203_s_1(.a(n203_1),.q0(n203_2),.q1(_w_1676));
  spl3L g221_s_0(.a(n221),.q0(n221_0),.q1(n221_1),.q2(n221_2));
  spl3L g225_s_0(.a(n225),.q0(n225_0),.q1(n225_1),.q2(n225_2));
  or_bb g546(.a(n491_1),.b(n513_1),.q(n546));
  spl3L g398_s_1(.a(n398_1),.q0(n398_2),.q1(n398_3),.q2(_w_1670));
  spl3L g227_s_0(.a(n227),.q0(n227_0),.q1(n227_1),.q2(n227_2));
  spl2 g337_s_1(.a(n337_2),.q0(n337_3),.q1(_w_1669));
  spl2 g160_s_0(.a(n160),.q0(n160_0),.q1(_w_1666));
  spl3L g541_s_0(.a(n541),.q0(n541_0),.q1(n541_1),.q2(_w_1663));
  spl3L g458_s_0(.a(n458),.q0(n458_0),.q1(n458_1),.q2(n458_2));
  maj_bbi g275(.a(n267_1),.b(n273_1),.c(n261_1),.q(_w_1662));
  and_bi g556(.a(n555),.b(n554),.q(out_6_));
  bfr _b_1078(.a(_w_1634),.q(n429));
  bfr _b_1172(.a(_w_1728),.q(n291_3));
  and_bi g553(.a(n552),.b(n551),.q(n553));
  and_bb g255(.a(n215_4),.b(n254_0),.q(n255));
  and_bb g176(.a(in_82_),.b(in_83_),.q(n176));
  and_bi g550(.a(n549),.b(n548),.q(_w_1657));
  and_bb g300(.a(n279_0),.b(n299_0),.q(n300));
  and_bi g540(.a(n539),.b(n349_0),.q(_w_1644));
  and_bb g297(.a(n280_0),.b(n296_0),.q(n297));
  bfr _b_758(.a(_w_1314),.q(_w_1315));
  and_bb g536(.a(n514_0),.b(n535_0),.q(n536));
  spl3L g430_s_0(.a(n430),.q0(n430_0),.q1(n430_1),.q2(n430_2));
  and_bi g535(.a(n534),.b(n533),.q(n535));
  or_bb g534(.a(n523_1),.b(n532_1),.q(n534));
  spl3L g543_s_0(.a(n543),.q0(n543_0),.q1(n543_1),.q2(_w_1638));
  spl2 g202_s_0(.a(n202),.q0(n202_0),.q1(n202_1));
  and_bb g533(.a(n523_0),.b(n532_0),.q(n533));
  spl2 g203_s_0(.a(n203),.q0(n203_0),.q1(_w_1635));
  and_bi g532(.a(n531),.b(n530),.q(n532));
  bfr _b_870(.a(_w_1426),.q(n329));
  or_bb g531(.a(n528_1),.b(n529_1),.q(n531));
  maj_bbb g529(.a(n499_2),.b(n506_2),.c(n510_2),.q(n529));
  or_bb g429(.a(n216_3),.b(n219_2),.q(_w_1634));
  and_bi g528(.a(n527),.b(n526),.q(n528));
  bfr _b_1027(.a(_w_1583),.q(_w_1584));
  spl2 g140_s_1(.a(n140_1),.q0(n140_2),.q1(_w_1630));
  and_bb g526(.a(n524_0),.b(n525_0),.q(n526));
  and_bb g288(.a(in_10_),.b(in_11_),.q(n288));
  maj_bbi g295(.a(n287_1),.b(n293_1),.c(n281_1),.q(_w_1629));
  spl2 g169_s_1(.a(n169_2),.q0(n169_3),.q1(n169_4));
  bfr _b_1083(.a(_w_1639),.q(_w_1640));
  and_bi g523(.a(n522),.b(n521),.q(n523));
  or_bb g522(.a(n515_1),.b(n520_1),.q(n522));
  bfr _b_1082(.a(_w_1638),.q(_w_1639));
  or_bb g519(.a(n516_1),.b(n517_1),.q(n519));
  and_bb g518(.a(n516_0),.b(n517_0),.q(n518));
  spl2 g403_s_0(.a(n403),.q0(n403_0),.q1(n403_1));
  bfr _b_1076(.a(_w_1632),.q(_w_1633));
  maj_bbb g516(.a(n395_4),.b(n398_4),.c(n475_2),.q(_w_1626));
  maj_bbb g510(.a(n426_0),.b(n439_2),.c(n452_2),.q(n510));
  or_bb g508(.a(n499_1),.b(n506_1),.q(n508));
  or_bb g555(.a(n542_1),.b(n553_1),.q(n555));
  spl3L g130_s_0(.a(n130),.q0(n130_0),.q1(n130_1),.q2(_w_1624));
  and_bb g507(.a(n499_0),.b(n506_0),.q(n507));
  or_bb g505(.a(n502_1),.b(n503_1),.q(n505));
  and_bb g497(.a(n495_0),.b(n496_0),.q(n497));
  bfr _b_945(.a(_w_1501),.q(_w_1502));
  spl3L g337_s_0(.a(n337),.q0(n337_0),.q1(n337_1),.q2(n337_2));
  spl2 g323_s_0(.a(n323),.q0(n323_0),.q1(n323_1));
  maj_bbb g503(.a(n440_0),.b(n443_2),.c(n446_2),.q(n503));
  or_bb g501(.a(n441_3),.b(n444_3),.q(n501));
  bfr _b_1102(.a(_w_1658),.q(_w_1659));
  or_bb g387(.a(n367_1),.b(n385_1),.q(n387));
  and_bi g499(.a(n498),.b(n497),.q(n499));
  bfr _b_864(.a(_w_1420),.q(n301));
  bfr _b_1069(.a(_w_1625),.q(n130_2));
  and_bi g495(.a(n494),.b(n493),.q(n495));
  bfr _b_801(.a(_w_1357),.q(n304_2));
  and_bb g489(.a(n471_0),.b(n488_0),.q(n489));
  and_bi g488(.a(n487),.b(n486),.q(n488));
  and_bb g483(.a(n481_0),.b(n482_0),.q(n483));
  and_bi g446(.a(n445),.b(n444_0),.q(n446));
  or_bb g378(.a(n320_2),.b(n376_1),.q(_w_1619));
  and_bi g251(.a(n250),.b(n249),.q(n251));
  and_bb g476(.a(n474_0),.b(n475_0),.q(n476));
  and_bi g474(.a(n473),.b(n472),.q(n474));
  or_bb g477(.a(n474_1),.b(n475_1),.q(n477));
  spl3L g542_s_0(.a(n542),.q0(n542_0),.q1(n542_1),.q2(n542_2));
  or_bb g480(.a(n407_3),.b(n410_3),.q(n480));
  and_bb g493(.a(n428_2),.b(n431_2),.q(n493));
  and_bi g470(.a(n469),.b(n468),.q(_w_1614));
  or_bb g469(.a(n349_5),.b(n467_1),.q(n469));
  and_bi g230(.a(n229),.b(n228),.q(n230));
  maj_bbb g160(.a(n157_0),.b(n158_0),.c(n159_0),.q(n160));
  and_bi g467(.a(n466),.b(n465),.q(n467));
  or_bb g305(.a(in_36_),.b(in_37_),.q(n305));
  and_bi g464(.a(n463),.b(n462),.q(_w_1611));
  bfr _b_1029(.a(_w_1585),.q(_w_1586));
  spl2 g240_s_1(.a(n240_1),.q0(n240_2),.q1(n240_3));
  or_bb g460(.a(n425_1),.b(n458_1),.q(n460));
  and_bi g458(.a(n457),.b(n456),.q(n458));
  maj_bbi g184(.a(n181_1),.b(n182_1),.c(n180_1),.q(_w_1610));
  and_bb g333(.a(in_50_),.b(in_51_),.q(n333));
  bfr _b_1040(.a(_w_1596),.q(_w_1597));
  bfr _b_917(.a(_w_1473),.q(_w_1474));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(n153_1));
  or_bb g264(.a(in_24_),.b(in_25_),.q(n264));
  and_bb g346(.a(n302_0),.b(n345_0),.q(n346));
  and_bi g455(.a(n454),.b(n453),.q(n455));
  or_bb g473(.a(n395_3),.b(n398_3),.q(n473));
  spl2 g553_s_0(.a(n553),.q0(n553_0),.q1(n553_1));
  bfr _b_873(.a(_w_1429),.q(_w_1430));
  and_bi g452(.a(n451),.b(n450),.q(n452));
  and_bi g461(.a(n460),.b(n459),.q(n461));
  spl3L g297_s_0(.a(n297),.q0(n297_0),.q1(n297_1),.q2(n297_2));
  spl2 g199_s_0(.a(n199),.q0(n199_0),.q1(n199_1));
  spl2 g455_s_0(.a(n455),.q0(n455_0),.q1(n455_1));
  spl2 g212_s_1(.a(n212_2),.q0(n212_3),.q1(n212_4));
  bfr _b_905(.a(_w_1461),.q(_w_1462));
  maj_bbb g183(.a(n180_0),.b(n181_0),.c(n182_0),.q(n183));
  and_bi g373(.a(n372),.b(n371_0),.q(n373));
  spl2 g326_s_0(.a(n326),.q0(n326_0),.q1(n326_1));
  and_bb g311(.a(in_42_),.b(in_43_),.q(n311));
  or_bb g448(.a(n443_1),.b(n446_1),.q(n448));
  spl3L g385_s_0(.a(n385),.q0(n385_0),.q1(n385_1),.q2(n385_2));
  and_bb g444(.a(n240_2),.b(n243_1),.q(n444));
  maj_bbb g240(.a(n197_2),.b(n203_2),.c(n206_1),.q(n240));
  spl2 g461_s_0(.a(n461),.q0(n461_0),.q1(n461_1));
  maj_bbb g440(.a(n212_1),.b(n239_2),.c(n245_2),.q(n440));
  and_bi g439(.a(n438),.b(n437),.q(n439));
  and_bi g409(.a(n408),.b(n407_0),.q(n409));
  and_bb g166(.a(n149_0),.b(n165_0),.q(n166));
  maj_bbb g482(.a(n409_2),.b(n412_2),.c(n416_0),.q(n482));
  bfr _b_803(.a(_w_1359),.q(n300_2));
  or_bb g438(.a(n427_3),.b(n436_1),.q(n438));
  and_bi g302(.a(n301),.b(n300_0),.q(n302));
  and_bb g437(.a(n427_2),.b(n436_0),.q(n437));
  and_bb g468(.a(n349_4),.b(n467_0),.q(n468));
  bfr _b_951(.a(_w_1507),.q(_w_1508));
  maj_bbb g525(.a(n441_4),.b(n444_4),.c(n503_2),.q(_w_1604));
  bfr _b_768(.a(_w_1324),.q(n485_2));
  or_bb g190(.a(n172_1),.b(n188_1),.q(_w_1609));
  and_bb g431(.a(n222_2),.b(n225_1),.q(n431));
  and_bi g430(.a(n429),.b(n428_0),.q(n430));
  or_bb g490(.a(n471_1),.b(n488_1),.q(n490));
  maj_bbb g427(.a(n169_1),.b(n221_2),.c(n227_2),.q(n427));
  and_bb g511(.a(n509_0),.b(n510_0),.q(n511));
  or_bb g152(.a(in_96_),.b(in_97_),.q(n152));
  and_bi g425(.a(n424),.b(n423),.q(n425));
  or_bb g424(.a(n393_3),.b(n422_1),.q(n424));
  bfr _b_1068(.a(_w_1624),.q(_w_1625));
  spl2 g427_s_1(.a(n427_1),.q0(n427_2),.q1(n427_3));
  and_bb g420(.a(n406_0),.b(n419_0),.q(n420));
  or_bb g418(.a(n415_1),.b(n416_3),.q(n418));
  spl2 g155_s_0(.a(n155),.q0(n155_0),.q1(_w_1600));
  bfr _b_942(.a(_w_1498),.q(_w_1499));
  and_bi g415(.a(n414),.b(n413),.q(n415));
  or_bb g414(.a(n409_1),.b(n412_1),.q(n414));
  spl2 g274_s_1(.a(n274_2),.q0(n274_3),.q1(_w_1721));
  and_bi g491(.a(n490),.b(n489),.q(n491));
  and_bi g443(.a(n442),.b(n441_0),.q(n443));
  and_bb g413(.a(n409_0),.b(n412_0),.q(n413));
  or_bb g261(.a(in_28_),.b(in_29_),.q(_w_1596));
  and_bb g407(.a(n374_2),.b(n377_1),.q(n407));
  or_bb g527(.a(n524_1),.b(n525_1),.q(n527));
  bfr _b_1108(.a(_w_1664),.q(_w_1665));
  spl2 g333_s_0(.a(n333),.q0(n333_0),.q1(n333_1));
  bfr _b_789(.a(_w_1345),.q(n334_3));
  and_bi g403(.a(n402),.b(n401),.q(n403));
  bfr _b_783(.a(_w_1339),.q(n410_4));
  spl2 g185_s_0(.a(n185),.q0(n185_0),.q1(n185_1));
  bfr _b_1075(.a(_w_1631),.q(_w_1632));
  or_bb g552(.a(n541_1),.b(n543_1),.q(n552));
  spl3L g219_s_0(.a(n219),.q0(n219_0),.q1(n219_1),.q2(n219_2));
  and_bi g397(.a(n396),.b(n395_0),.q(n397));
  maj_bbb g394(.a(n300_1),.b(n355_2),.c(n361_2),.q(n394));
  or_bb g366(.a(n300_4),.b(n364_1),.q(n366));
  bfr _b_912(.a(_w_1468),.q(_w_1469));
  maj_bbb g392(.a(n257_0),.b(n349_2),.c(n391_0),.q(n392));
  and_bb g389(.a(n346_4),.b(n388_0),.q(n389));
  and_bi g388(.a(n387),.b(n386),.q(n388));
  and_bi g168(.a(n167),.b(n166_0),.q(n168));
  maj_bbi g296(.a(n281_2),.b(n295),.c(n294_0),.q(n296));
  and_bi g382(.a(n381),.b(n380),.q(n382));
  maj_bbb g426(.a(n215_2),.b(n233_2),.c(n251_2),.q(n426));
  bfr _b_882(.a(_w_1438),.q(n349_3));
  and_bi g406(.a(n405),.b(n404),.q(n406));
  spl2 g197_s_1(.a(n197_1),.q0(n197_2),.q1(_w_1690));
  spl2 g234_s_1(.a(n234_1),.q0(n234_2),.q1(n234_3));
  spl2 g196_s_0(.a(n196),.q0(n196_0),.q1(n196_1));
  and_bi g509(.a(n508),.b(n507),.q(n509));
  bfr _b_1145(.a(_w_1701),.q(_w_1702));
  spl2 g269_s_0(.a(n269),.q0(n269_0),.q1(n269_1));
  or_bb g151(.a(in_100_),.b(in_101_),.q(n151));
  and_bi g436(.a(n435),.b(n434),.q(n436));
  and_bi g148(.a(n147),.b(n146_0),.q(n148));
  and_bb g249(.a(n212_3),.b(n248_0),.q(n249));
  and_bb g246(.a(n239_0),.b(n245_0),.q(n246));
  maj_bbb g542(.a(n514_2),.b(n523_2),.c(n532_2),.q(n542));
  bfr _b_778(.a(_w_1334),.q(_w_1335));
  and_bb g551(.a(n541_0),.b(n543_0),.q(n551));
  or_bb g232(.a(n169_4),.b(n230_1),.q(n232));
  and_bi g449(.a(n448),.b(n447),.q(n449));
  and_bb g231(.a(n169_3),.b(n230_0),.q(n231));
  bfr _b_1067(.a(_w_1623),.q(n131_2));
  or_bb g229(.a(n221_1),.b(n227_1),.q(n229));
  and_bi g221(.a(n220),.b(n219_0),.q(n221));
  or_bb g247(.a(n239_1),.b(n245_1),.q(n247));
  and_bi g248(.a(n247),.b(n246),.q(n248));
  and_bi g245(.a(n244),.b(n243_0),.q(n245));
  or_bb g408(.a(n374_3),.b(n377_2),.q(_w_1591));
  maj_bbb g222(.a(n155_2),.b(n160_2),.c(n163_1),.q(n222));
  or_bb g220(.a(n146_2),.b(n218_1),.q(_w_1590));
  and_bb g521(.a(n515_0),.b(n520_0),.q(n521));
  or_bb g549(.a(n492_2),.b(n547_1),.q(n549));
  bfr _b_787(.a(_w_1343),.q(_w_1344));
  spl3L g282_s_0(.a(n282),.q0(n282_0),.q1(n282_1),.q2(_w_1588));
  spl3L g157_s_0(.a(n157),.q0(n157_0),.q1(n157_1),.q2(_w_1694));
  and_bi g400(.a(n399),.b(n398_0),.q(n400));
  bfr _b_867(.a(_w_1423),.q(n314_1));
  bfr _b_1023(.a(_w_1579),.q(_w_1580));
  and_bi g385(.a(n384),.b(n383),.q(n385));
  bfr _b_875(.a(_w_1431),.q(n324));
  bfr _b_1025(.a(_w_1581),.q(_w_1582));
  bfr _b_863(.a(_w_1419),.q(n174_2));
  and_bb g371(.a(n340_1),.b(n370_0),.q(n371));
  maj_bbi g242(.a(n206_4),.b(n241),.c(n240_0),.q(n242));
  bfr _b_957(.a(_w_1513),.q(n172));
  and_bb g359(.a(n297_1),.b(n358_0),.q(n359));
  or_bb g213(.a(n191_1),.b(n211_1),.q(_w_1578));
  spl2 g293_s_0(.a(n293),.q0(n293_0),.q1(n293_1));
  maj_bbi g208(.a(n193_2),.b(n207),.c(n206_0),.q(n208));
  spl2 g183_s_1(.a(n183_1),.q0(n183_2),.q1(_w_1577));
  or_bb g210(.a(n192_1),.b(n208_1),.q(_w_1575));
  or_bb g174(.a(in_84_),.b(in_85_),.q(n174));
  bfr _b_861(.a(_w_1417),.q(n372));
  and_bb g209(.a(n192_0),.b(n208_0),.q(n209));
  maj_bbb g163(.a(n150_0),.b(n156_0),.c(n162_0),.q(n163));
  or_bb g360(.a(n297_2),.b(n358_1),.q(_w_1587));
  bfr _b_769(.a(_w_1325),.q(_w_1326));
  spl3L g517_s_0(.a(n517),.q0(n517_0),.q1(n517_1),.q2(_w_1707));
  or_bb g147(.a(n129_1),.b(n145_1),.q(_w_1608));
  or_bb g421(.a(n406_1),.b(n419_1),.q(n421));
  and_bi g485(.a(n484),.b(n483),.q(n485));
  and_bi g322(.a(n321),.b(n320_0),.q(n322));
  spl2 g342_s_0(.a(n342),.q0(n342_0),.q1(n342_1));
  spl2 g302_s_0(.a(n302),.q0(n302_0),.q1(n302_1));
  and_bi g364(.a(n363),.b(n362),.q(n364));
  maj_bbi g272(.a(n269_1),.b(n270_1),.c(n268_1),.q(_w_1569));
  or_bb g258(.a(n171_1),.b(n214_1),.q(_w_1568));
  maj_bbi g204(.a(n201_1),.b(n202_1),.c(n200_1),.q(_w_1567));
  or_bb g226(.a(n166_2),.b(n224_1),.q(_w_1566));
  spl2 g162_s_0(.a(n162),.q0(n162_0),.q1(n162_1));
  spl2 g416_s_1(.a(n416_1),.q0(n416_2),.q1(n416_3));
  maj_bbi g217(.a(n134_3),.b(n140_3),.c(n143_3),.q(n217));
  spl2 g263_s_0(.a(n263),.q0(n263_0),.q1(n263_1));
  spl2 g222_s_0(.a(n222),.q0(n222_0),.q1(_w_1715));
  and_bb g225(.a(n166_1),.b(n224_0),.q(n225));
  spl2 g488_s_0(.a(n488),.q0(n488_0),.q1(n488_1));
  and_bi g481(.a(n480),.b(n479),.q(n481));
  bfr _b_1056(.a(_w_1612),.q(_w_1613));
  maj_bbb g274(.a(n261_0),.b(n267_0),.c(n273_0),.q(n274));
  and_bi g478(.a(n477),.b(n476),.q(n478));
  maj_bbb g203(.a(n200_0),.b(n201_0),.c(n202_0),.q(n203));
  spl3L g137_s_0(.a(n137),.q0(n137_0),.q1(n137_1),.q2(_w_1564));
  or_bb g457(.a(n426_3),.b(n455_1),.q(n457));
  and_bb g201(.a(in_70_),.b(in_71_),.q(n201));
  spl2 g133_s_0(.a(n133),.q0(n133_0),.q1(n133_1));
  maj_bbi g154(.a(n152_0),.b(n153_0),.c(n151_0),.q(_w_1563));
  spl3L g163_s_0(.a(n163),.q0(n163_0),.q1(n163_1),.q2(n163_2));
  maj_bbi g199(.a(n194_2),.b(n198),.c(n197_0),.q(n199));
  maj_bbi g292(.a(n289_1),.b(n290_1),.c(n288_1),.q(_w_1562));
  or_bb g343(.a(n322_0),.b(n342_0),.q(_w_1561));
  bfr _b_1112(.a(_w_1668),.q(n160_1));
  maj_bbb g206(.a(n193_0),.b(n199_0),.c(n205_0),.q(n206));
  spl2 g346_s_1(.a(n346_1),.q0(n346_2),.q1(_w_1559));
  and_bi g214(.a(n213),.b(n212_0),.q(n214));
  maj_bbi g198(.a(n195_1),.b(n196_1),.c(n194_1),.q(_w_1558));
  or_bb g175(.a(in_80_),.b(in_81_),.q(n175));
  maj_bbb g393(.a(n346_2),.b(n367_2),.c(n385_2),.q(n393));
  or_bb g396(.a(n350_3),.b(n354_2),.q(_w_1556));
  and_bi g191(.a(n190),.b(n189_0),.q(n191));
  or_bb g182(.a(in_88_),.b(in_89_),.q(n182));
  spl3L g397_s_0(.a(n397),.q0(n397_0),.q1(n397_1),.q2(n397_2));
  and_bi g520(.a(n519),.b(n518),.q(n520));
  bfr _b_998(.a(_w_1554),.q(n129));
  maj_bbi g241(.a(n197_3),.b(n203_3),.c(n206_3),.q(n241));
  spl3L g274_s_0(.a(n274),.q0(n274_0),.q1(n274_1),.q2(n274_2));
  spl2 g160_s_1(.a(n160_1),.q0(n160_2),.q1(_w_1693));
  maj_bbb g291(.a(n288_0),.b(n289_0),.c(n290_0),.q(n291));
  bfr _b_1117(.a(_w_1673),.q(_w_1674));
  maj_bbi g187(.a(n179_1),.b(n185_1),.c(n173_1),.q(_w_1555));
  and_bb g129(.a(in_126_),.b(in_127_),.q(_w_1547));
  spl2 g287_s_0(.a(n287),.q0(n287_0),.q1(n287_1));
  and_bb g423(.a(n393_2),.b(n422_0),.q(n423));
  bfr _b_1073(.a(_w_1629),.q(n295));
  maj_bbb g155(.a(n151_1),.b(n152_1),.c(n153_1),.q(n155));
  maj_bbi g338(.a(n330_1),.b(n336_1),.c(n324_1),.q(_w_1546));
  spl2 g242_s_0(.a(n242),.q0(n242_0),.q1(n242_1));
  bfr _b_1165(.a(_w_1721),.q(n274_4));
  maj_bbi g218(.a(n143_4),.b(n217),.c(n216_0),.q(n218));
  or_bb g487(.a(n478_1),.b(n485_1),.q(n487));
  bfr _b_1123(.a(_w_1679),.q(_w_1680));
  and_bb g196(.a(in_66_),.b(in_67_),.q(n196));
  maj_bbi g310(.a(n305_2),.b(n309),.c(n308_0),.q(n310));
  spl2 g294_s_1(.a(n294_2),.q0(n294_3),.q1(_w_1576));
  spl2 g368_s_1(.a(n368_1),.q0(n368_2),.q1(n368_3));
  spl2 g431_s_0(.a(n431),.q0(n431_0),.q1(n431_1));
  spl2 g205_s_0(.a(n205),.q0(n205_0),.q1(n205_1));
  bfr _b_1093(.a(_w_1649),.q(_w_1650));
  spl3L g325_s_0(.a(n325),.q0(n325_0),.q1(n325_1),.q2(_w_1726));
  or_bb g331(.a(in_52_),.b(in_53_),.q(n331));
  and_bb g380(.a(n373_0),.b(n379_0),.q(n380));
  bfr _b_772(.a(_w_1328),.q(_w_1329));
  or_bb g268(.a(in_20_),.b(in_21_),.q(n268));
  and_bb g459(.a(n425_0),.b(n458_0),.q(n459));
  or_bb g244(.a(n209_2),.b(n242_1),.q(_w_1545));
  maj_bbi g235(.a(n177_3),.b(n183_3),.c(n186_3),.q(n235));
  and_bb g149(.a(in_110_),.b(in_111_),.q(_w_1537));
  bfr _b_767(.a(_w_1323),.q(_w_1324));
  spl2 g474_s_0(.a(n474),.q0(n474_0),.q1(n474_1));
  or_bb g384(.a(n344_4),.b(n382_1),.q(n384));
  bfr _b_858(.a(_w_1414),.q(_w_1415));
  maj_bbi g318(.a(n310_1),.b(n316_1),.c(n304_1),.q(_w_1534));
  maj_bbb g515(.a(n471_2),.b(n478_2),.c(n485_2),.q(n515));
  bfr _b_880(.a(_w_1436),.q(out_7_));
  bfr _b_1130(.a(_w_1686),.q(_w_1687));
  bfr _b_890(.a(_w_1446),.q(_w_1447));
  maj_bbi g144(.a(n136_1),.b(n142_1),.c(n130_1),.q(_w_1533));
  spl2 g214_s_0(.a(n214),.q0(n214_0),.q1(n214_1));
  and_bb g158(.a(in_102_),.b(in_103_),.q(n158));
  spl2 g284_s_0(.a(n284),.q0(n284_0),.q1(n284_1));
  bfr _b_797(.a(_w_1353),.q(_w_1354));
  spl3L g131_s_0(.a(n131),.q0(n131_0),.q1(n131_1),.q2(_w_1622));
  spl2 g547_s_0(.a(n547),.q0(n547_0),.q1(n547_1));
  and_bb g312(.a(in_38_),.b(in_39_),.q(n312));
  maj_bbi g141(.a(n138_1),.b(n139_1),.c(n137_1),.q(_w_1532));
  maj_bbb g368(.a(n328_2),.b(n334_2),.c(n337_1),.q(n368));
  maj_bbi g179(.a(n174_2),.b(n178),.c(n177_0),.q(n179));
  maj_bbi g164(.a(n156_1),.b(n162_1),.c(n150_1),.q(_w_1531));
  maj_bbb g140(.a(n137_0),.b(n138_0),.c(n139_0),.q(n140));
  and_bb g479(.a(n407_2),.b(n410_2),.q(n479));
  and_bb g447(.a(n443_0),.b(n446_0),.q(n447));
  and_bi g506(.a(n505),.b(n504),.q(n506));
  bfr _b_1155(.a(_w_1711),.q(_w_1712));
  and_bb g192(.a(in_78_),.b(in_79_),.q(_w_1523));
  spl3L g492_s_0(.a(n492),.q0(n492_0),.q1(n492_1),.q2(n492_2));
  and_bb g530(.a(n528_0),.b(n529_0),.q(n530));
  maj_bbi g286(.a(n283_1),.b(n284_1),.c(n282_1),.q(_w_1522));
  spl2 g330_s_0(.a(n330),.q0(n330_0),.q1(n330_1));
  and_bb g243(.a(n209_1),.b(n242_0),.q(n243));
  spl2 g440_s_1(.a(n440_1),.q0(n440_2),.q1(n440_3));
  bfr _b_1180(.a(_w_1736),.q(n150));
  maj_bbb g496(.a(n427_0),.b(n430_2),.c(n433_2),.q(n496));
  maj_bbb g356(.a(n285_2),.b(n291_2),.c(n294_1),.q(n356));
  bfr _b_944(.a(_w_1500),.q(_w_1501));
  bfr _b_970(.a(_w_1526),.q(_w_1527));
  bfr _b_1079(.a(_w_1635),.q(_w_1636));
  spl2 g215_s_2(.a(n215_3),.q0(n215_4),.q1(n215_5));
  bfr _b_816(.a(_w_1372),.q(_w_1373));
  maj_bbi g207(.a(n199_1),.b(n205_1),.c(n193_1),.q(_w_1574));
  maj_bbb g265(.a(n262_0),.b(n263_0),.c(n264_0),.q(n265));
  bfr _b_1132(.a(_w_1688),.q(_w_1689));
  maj_bbb g517(.a(n407_4),.b(n410_4),.c(n482_2),.q(_w_1519));
  and_bb g289(.a(in_6_),.b(in_7_),.q(n289));
  bfr _b_814(.a(_w_1370),.q(n499_2));
  or_bb g321(.a(n303_1),.b(n319_1),.q(_w_1607));
  maj_bbi g161(.a(n158_1),.b(n159_1),.c(n157_1),.q(_w_1518));
  maj_bbb g294(.a(n281_0),.b(n287_0),.c(n293_0),.q(n294));
  maj_bbb g514(.a(n491_2),.b(n492_0),.c(n513_2),.q(n514));
  and_bb g137(.a(in_122_),.b(in_123_),.q(n137));
  spl2 g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1));
  spl2 g314_s_1(.a(n314_1),.q0(n314_2),.q1(_w_1603));
  and_bi g171(.a(n170),.b(n169_0),.q(n171));
  spl3L g377_s_0(.a(n377),.q0(n377_0),.q1(n377_1),.q2(n377_2));
  maj_bbi g185(.a(n180_2),.b(n184),.c(n183_0),.q(n185));
  and_bb g548(.a(n492_1),.b(n547_0),.q(n548));
  spl3L g452_s_0(.a(n452),.q0(n452_0),.q1(n452_1),.q2(n452_2));
  maj_bbi g162(.a(n157_2),.b(n161),.c(n160_0),.q(n162));
  and_bb g237(.a(n189_1),.b(n236_0),.q(n237));
  spl2 g395_s_0(.a(n395),.q0(n395_0),.q1(n395_1));
  and_bb g441(.a(n234_2),.b(n237_1),.q(n441));
  or_bb g250(.a(n212_4),.b(n248_1),.q(n250));
  spl2 g312_s_0(.a(n312),.q0(n312_0),.q1(n312_1));
  bfr _b_853(.a(_w_1409),.q(_w_1410));
  maj_bbi g135(.a(n132_1),.b(n133_1),.c(n131_1),.q(_w_1517));
  maj_bbb g543(.a(n524_2),.b(n525_2),.c(n529_2),.q(_w_1514));
  and_bb g354(.a(n277_1),.b(n352_0),.q(n354));
  or_bb g283(.a(in_0_),.b(in_1_),.q(n283));
  and_bb g326(.a(in_54_),.b(in_55_),.q(n326));
  bfr _b_938(.a(_w_1494),.q(n399));
  or_bb g484(.a(n481_1),.b(n482_1),.q(n484));
  and_bb g172(.a(in_94_),.b(in_95_),.q(_w_1506));
  spl2 g138_s_0(.a(n138),.q0(n138_0),.q1(n138_1));
  bfr _b_1000(.a(_w_1556),.q(n396));
  maj_bbb g492(.a(n392_0),.b(n425_2),.c(n458_2),.q(n492));
  maj_bbb g374(.a(n308_2),.b(n314_2),.c(n317_1),.q(n374));
  bfr _b_914(.a(_w_1470),.q(_w_1471));
  and_bb g138(.a(in_118_),.b(in_119_),.q(n138));
  maj_bbi g223(.a(n155_3),.b(n160_3),.c(n163_3),.q(n223));
  bfr _b_829(.a(_w_1385),.q(n216_1));
  bfr _b_1061(.a(_w_1617),.q(_w_1618));
  and_bb g434(.a(n430_0),.b(n433_0),.q(n434));
  bfr _b_983(.a(_w_1539),.q(_w_1540));
  spl2 g165_s_0(.a(n165),.q0(n165_0),.q1(n165_1));
  bfr _b_1051(.a(_w_1607),.q(n321));
  maj_bbi g224(.a(n163_4),.b(n223),.c(n222_0),.q(n224));
  or_bb g512(.a(n509_1),.b(n510_1),.q(n512));
  or_bb g445(.a(n240_3),.b(n243_2),.q(_w_1505));
  or_bb g256(.a(n215_5),.b(n254_1),.q(n256));
  bfr _b_791(.a(_w_1347),.q(_w_1348));
  maj_bbb g197(.a(n194_0),.b(n195_0),.c(n196_0),.q(n197));
  spl3L g166_s_0(.a(n166),.q0(n166_0),.q1(n166_1),.q2(n166_2));
  bfr _b_820(.a(_w_1376),.q(_w_1377));
  spl2 g290_s_0(.a(n290),.q0(n290_0),.q1(n290_1));
  spl3L g189_s_0(.a(n189),.q0(n189_0),.q1(n189_1),.q2(n189_2));
  spl3L g200_s_0(.a(n200),.q0(n200_0),.q1(n200_1),.q2(_w_1503));
  spl2 g358_s_0(.a(n358),.q0(n358_0),.q1(n358_1));
  and_bb g303(.a(in_46_),.b(in_47_),.q(_w_1495));
  bfr _b_874(.a(_w_1430),.q(_w_1431));
  and_bi g547(.a(n546),.b(n545),.q(n547));
  or_bb g399(.a(n356_3),.b(n359_2),.q(_w_1494));
  or_bb g381(.a(n373_1),.b(n379_1),.q(n381));
  spl3L g407_s_1(.a(n407_1),.q0(n407_2),.q1(n407_3),.q2(_w_1491));
  or_bb g435(.a(n430_1),.b(n433_1),.q(n435));
  or_bb g167(.a(n149_1),.b(n165_1),.q(_w_1490));
  spl3L g475_s_0(.a(n475),.q0(n475_0),.q1(n475_1),.q2(n475_2));
  and_bb g417(.a(n415_0),.b(n416_2),.q(n417));
  bfr _b_1045(.a(_w_1601),.q(_w_1602));
  or_bb g306(.a(in_32_),.b(in_33_),.q(n306));
  bfr _b_1091(.a(_w_1647),.q(_w_1648));
  or_bb g539(.a(n259_1),.b(n348_1),.q(_w_1489));
  bfr _b_1072(.a(_w_1628),.q(n516));
  bfr _b_1115(.a(_w_1671),.q(_w_1672));
  or_bb g454(.a(n439_1),.b(n452_1),.q(n454));
  and_bi g233(.a(n232),.b(n231),.q(n233));
  and_bb g465(.a(n257_1),.b(n391_1),.q(n465));
  or_bb g304(.a(in_44_),.b(in_45_),.q(_w_1570));
  bfr _b_1018(.a(_w_1574),.q(n207));
  maj_bbb g234(.a(n177_2),.b(n183_2),.c(n186_1),.q(n234));
  spl2 g129_s_0(.a(n129),.q0(n129_0),.q1(n129_1));
  or_bb g195(.a(in_64_),.b(in_65_),.q(n195));
  bfr _b_1049(.a(_w_1605),.q(_w_1606));
  spl2 g296_s_0(.a(n296),.q0(n296_0),.q1(n296_1));
  spl2 g279_s_0(.a(n279),.q0(n279_0),.q1(n279_1));
  bfr _b_795(.a(_w_1351),.q(n328_3));
  or_bb g170(.a(n148_1),.b(n168_1),.q(_w_1488));
  spl2 g291_s_0(.a(n291),.q0(n291_0),.q1(_w_1485));
  spl2 g155_s_1(.a(n155_1),.q0(n155_2),.q1(_w_1696));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(n179_1));
  maj_bbb g177(.a(n174_0),.b(n175_0),.c(n176_0),.q(n177));
  or_bb g193(.a(in_76_),.b(in_77_),.q(_w_1481));
  bfr _b_926(.a(_w_1482),.q(_w_1483));
  and_bb g428(.a(n216_2),.b(n219_1),.q(n428));
  maj_bbb g471(.a(n393_0),.b(n406_2),.c(n419_2),.q(n471));
  and_bi g257(.a(n256),.b(n255),.q(n257));
  and_bi g538(.a(n537),.b(n536),.q(_w_1642));
  and_bi g412(.a(n411),.b(n410_0),.q(n412));
  bfr _b_915(.a(_w_1471),.q(_w_1472));
  maj_bbb g216(.a(n134_2),.b(n140_2),.c(n143_1),.q(n216));
  and_bb g228(.a(n221_0),.b(n227_0),.q(n228));
  or_bb g131(.a(in_116_),.b(in_117_),.q(n131));
  or_bb g202(.a(in_72_),.b(in_73_),.q(n202));
  bfr _b_1150(.a(_w_1706),.q(n346_1));
  spl2 g283_s_0(.a(n283),.q0(n283_0),.q1(n283_1));
  maj_bbb g186(.a(n173_0),.b(n179_0),.c(n185_0),.q(n186));
  maj_bbi g178(.a(n175_1),.b(n176_1),.c(n174_1),.q(_w_1477));
  maj_bbb g134(.a(n131_0),.b(n132_0),.c(n133_0),.q(n134));
  bfr _b_1092(.a(_w_1648),.q(_w_1649));
  or_bb g327(.a(in_56_),.b(in_57_),.q(n327));
  spl3L g324_s_0(.a(n324),.q0(n324_0),.q1(n324_1),.q2(_w_1475));
  spl2 g215_s_1(.a(n215_1),.q0(n215_2),.q1(_w_1473));
  and_bb g410(.a(n368_2),.b(n371_1),.q(n410));
  bfr _b_807(.a(_w_1363),.q(n285_1));
  and_bb g260(.a(in_30_),.b(in_31_),.q(_w_1465));
  and_bi g419(.a(n418),.b(n417),.q(n419));
  and_bb g262(.a(in_26_),.b(in_27_),.q(n262));
  maj_bbi g236(.a(n186_4),.b(n235),.c(n234_0),.q(n236));
  or_bb g282(.a(in_4_),.b(in_5_),.q(n282));
  and_bb g263(.a(in_22_),.b(in_23_),.q(n263));
  or_bb g341(.a(n323_1),.b(n339_1),.q(_w_1661));
  bfr _b_1047(.a(_w_1603),.q(n314_3));
  maj_bbi g267(.a(n262_2),.b(n266),.c(n265_0),.q(n267));
  or_bb g269(.a(in_16_),.b(in_17_),.q(n269));
  maj_bbi g287(.a(n282_2),.b(n286),.c(n285_0),.q(n287));
  and_bb g404(.a(n394_2),.b(n403_0),.q(n404));
  maj_bbb g308(.a(n305_0),.b(n306_0),.c(n307_0),.q(n308));
  bfr _b_1134(.a(_w_1690),.q(n197_3));
  maj_bbb g524(.a(n428_4),.b(n431_4),.c(n496_2),.q(_w_1478));
  spl3L g317_s_0(.a(n317),.q0(n317_0),.q1(n317_1),.q2(n317_2));
  and_bb g270(.a(in_18_),.b(in_19_),.q(n270));
  spl3L g373_s_0(.a(n373),.q0(n373_0),.q1(n373_1),.q2(n373_2));
  spl2 g171_s_0(.a(n171),.q0(n171_0),.q1(n171_1));
  maj_bbi g315(.a(n312_1),.b(n313_1),.c(n311_1),.q(_w_1464));
  spl2 g230_s_0(.a(n230),.q0(n230_0),.q1(n230_1));
  or_bb g298(.a(n280_1),.b(n296_1),.q(_w_1463));
  and_bi g379(.a(n378),.b(n377_0),.q(n379));
  maj_bbi g276(.a(n261_2),.b(n275),.c(n274_0),.q(n276));
  and_bb g280(.a(in_14_),.b(in_15_),.q(_w_1451));
  maj_bbi g335(.a(n332_1),.b(n333_1),.c(n331_1),.q(_w_1450));
  spl2 g134_s_1(.a(n134_1),.q0(n134_2),.q1(_w_1557));
  spl3L g311_s_0(.a(n311),.q0(n311_0),.q1(n311_1),.q2(_w_1448));
  bfr _b_1087(.a(_w_1643),.q(out_5_));
  or_bb g281(.a(in_12_),.b(in_13_),.q(_w_1444));
  spl2 g349_s_2(.a(n349_3),.q0(n349_4),.q1(n349_5));
  bfr _b_1039(.a(_w_1595),.q(n411));
  bfr _b_859(.a(_w_1415),.q(_w_1416));
  or_bb g132(.a(in_112_),.b(in_113_),.q(n132));
  and_bb g277(.a(n260_0),.b(n276_0),.q(n277));
  spl3L g194_s_0(.a(n194),.q0(n194_0),.q1(n194_1),.q2(_w_1442));
  maj_bbb g285(.a(n282_0),.b(n283_0),.c(n284_0),.q(n285));
  or_bb g290(.a(in_8_),.b(in_9_),.q(n290));
  and_bb g200(.a(in_74_),.b(in_75_),.q(n200));
  or_bb g353(.a(n277_2),.b(n352_1),.q(_w_1441));
  bfr _b_794(.a(_w_1350),.q(n331_2));
  bfr _b_1095(.a(_w_1651),.q(_w_1652));
  bfr _b_819(.a(_w_1375),.q(n317_4));
  bfr _b_900(.a(_w_1456),.q(_w_1457));
  bfr _b_1028(.a(_w_1584),.q(_w_1585));
  maj_bbb g334(.a(n331_0),.b(n332_0),.c(n333_0),.q(n334));
  maj_bbi g330(.a(n325_2),.b(n329),.c(n328_0),.q(n330));
  bfr _b_898(.a(_w_1454),.q(_w_1455));
  or_bb g432(.a(n222_3),.b(n225_2),.q(_w_1440));
  and_bb g456(.a(n426_2),.b(n455_0),.q(n456));
  bfr _b_928(.a(_w_1484),.q(n193));
  or_bb g278(.a(n260_1),.b(n276_1),.q(_w_1459));
  spl2 g148_s_0(.a(n148),.q0(n148_0),.q1(n148_1));
  maj_bbi g309(.a(n306_1),.b(n307_1),.c(n305_1),.q(_w_1439));
  or_bb g390(.a(n346_5),.b(n388_1),.q(n390));
  maj_bbb g544(.a(n541_2),.b(n542_2),.c(n543_2),.q(_w_1436));
  spl3L g496_s_0(.a(n496),.q0(n496_0),.q1(n496_1),.q2(n496_2));
  bfr _b_757(.a(_w_1313),.q(n234_1));
  bfr _b_927(.a(_w_1483),.q(_w_1484));
  spl2 g186_s_1(.a(n186_2),.q0(n186_3),.q1(_w_1435));
  and_bb g395(.a(n350_2),.b(n354_1),.q(n395));
  and_bi g391(.a(n390),.b(n389),.q(n391));
  spl3L g173_s_0(.a(n173),.q0(n173_0),.q1(n173_1),.q2(_w_1433));
  bfr _b_891(.a(_w_1447),.q(n281));
  bfr _b_759(.a(_w_1315),.q(_w_1316));
  maj_bbi g357(.a(n285_3),.b(n291_3),.c(n294_3),.q(n357));
  bfr _b_818(.a(_w_1374),.q(n265_1));
  bfr _b_981(.a(_w_1537),.q(_w_1538));
  and_bi g433(.a(n432),.b(n431_0),.q(n433));
  bfr _b_1109(.a(_w_1665),.q(n541_2));
  spl2 g143_s_1(.a(n143_2),.q0(n143_3),.q1(_w_1432));
  bfr _b_809(.a(_w_1365),.q(n268_2));
  or_bb g324(.a(in_60_),.b(in_61_),.q(_w_1428));
  or_bb g442(.a(n234_3),.b(n237_2),.q(_w_1427));
  maj_bbb g328(.a(n325_0),.b(n326_0),.c(n327_0),.q(n328));
  maj_bbi g329(.a(n326_1),.b(n327_1),.c(n325_1),.q(_w_1426));
  maj_bbi g339(.a(n324_2),.b(n338),.c(n337_0),.q(n339));
  and_bi g211(.a(n210),.b(n209_0),.q(n211));
  spl2 g370_s_0(.a(n370),.q0(n370_0),.q1(n370_1));
  and_bi g345(.a(n343),.b(n344_0),.q(n345));
  maj_bbi g376(.a(n317_4),.b(n375),.c(n374_0),.q(n376));
  maj_bbi g165(.a(n150_2),.b(n164),.c(n163_0),.q(n165));
  bfr _b_999(.a(_w_1555),.q(n187));
  and_bb g365(.a(n300_3),.b(n364_0),.q(n365));
  maj_bbi g336(.a(n331_2),.b(n335),.c(n334_0),.q(n336));
  or_bb g405(.a(n394_3),.b(n403_1),.q(n405));
  maj_bbb g337(.a(n324_0),.b(n330_0),.c(n336_0),.q(n337));
  bfr _b_780(.a(_w_1336),.q(n356_1));
  spl2 g163_s_1(.a(n163_2),.q0(n163_3),.q1(_w_1425));
  bfr _b_856(.a(_w_1412),.q(_w_1413));
  bfr _b_849(.a(_w_1405),.q(_w_1406));
  and_bb g554(.a(n542_0),.b(n553_0),.q(n554));
  maj_bbb g143(.a(n130_0),.b(n136_0),.c(n142_0),.q(n143));
  bfr _b_1181(.a(_w_1737),.q(_w_1738));
  bfr _b_1103(.a(_w_1659),.q(_w_1660));
  spl2 g428_s_0(.a(n428),.q0(n428_0),.q1(n428_1));
  and_bb g340(.a(n323_0),.b(n339_0),.q(n340));
  bfr _b_964(.a(_w_1520),.q(_w_1521));
  and_bb g377(.a(n320_1),.b(n376_0),.q(n377));
  and_bi g342(.a(n341),.b(n340_0),.q(n342));
  spl2 g236_s_0(.a(n236),.q0(n236_0),.q1(n236_1));
  spl3L g239_s_0(.a(n239),.q0(n239_0),.q1(n239_1),.q2(n239_2));
  or_bb g238(.a(n189_2),.b(n236_1),.q(_w_1424));
  maj_bbi g316(.a(n311_2),.b(n315),.c(n314_0),.q(n316));
  spl2 g314_s_0(.a(n314),.q0(n314_0),.q1(_w_1421));
  and_bi g259(.a(n258),.b(n215_0),.q(n259));
  and_bb g344(.a(n322_1),.b(n342_1),.q(n344));
  and_bi g502(.a(n501),.b(n500),.q(n502));
  bfr _b_904(.a(_w_1460),.q(_w_1461));
  maj_bbb g350(.a(n265_2),.b(n271_2),.c(n274_1),.q(n350));
  bfr _b_770(.a(_w_1326),.q(_w_1327));
  bfr _b_940(.a(_w_1496),.q(_w_1497));
  bfr _b_781(.a(_w_1337),.q(_w_1338));
  bfr _b_1024(.a(_w_1580),.q(_w_1581));
  maj_bbi g352(.a(n274_4),.b(n351),.c(n350_0),.q(n352));
  and_bi g355(.a(n353),.b(n354_0),.q(n355));
  spl2 g168_s_0(.a(n168),.q0(n168_0),.q1(n168_1));
  spl3L g146_s_0(.a(n146),.q0(n146_0),.q1(n146_1),.q2(n146_2));
  spl2 g156_s_0(.a(n156),.q0(n156_0),.q1(n156_1));
  spl3L g174_s_0(.a(n174),.q0(n174_0),.q1(n174_1),.q2(_w_1418));
  maj_bbb g475(.a(n394_0),.b(n397_2),.c(n400_2),.q(n475));
  spl2 g393_s_1(.a(n393_1),.q0(n393_2),.q1(n393_3));
  and_bb g545(.a(n491_0),.b(n513_0),.q(n545));
  maj_bbi g358(.a(n294_4),.b(n357),.c(n356_0),.q(n358));
  bfr _b_1142(.a(_w_1698),.q(_w_1699));
  spl2 g449_s_0(.a(n449),.q0(n449_0),.q1(n449_1));
  spl2 g344_s_1(.a(n344_2),.q0(n344_3),.q1(n344_4));
  or_bb g498(.a(n495_1),.b(n496_1),.q(n498));
  spl2 g313_s_0(.a(n313),.q0(n313_0),.q1(n313_1));
  spl2 g218_s_0(.a(n218),.q0(n218_0),.q1(n218_1));
  and_bb g320(.a(n303_0),.b(n319_0),.q(n320));
  and_bi g361(.a(n360),.b(n359_0),.q(n361));
  or_bb g363(.a(n355_1),.b(n361_1),.q(n363));
  spl3L g169_s_0(.a(n169),.q0(n169_0),.q1(n169_1),.q2(_w_1412));
  spl2 g327_s_0(.a(n327),.q0(n327_0),.q1(n327_1));
  bfr _b_838(.a(_w_1394),.q(_w_1395));
  and_bi g254(.a(n253),.b(n252),.q(n254));
  maj_bbi g369(.a(n328_3),.b(n334_3),.c(n337_3),.q(n369));
  spl3L g431_s_1(.a(n431_1),.q0(n431_2),.q1(n431_3),.q2(_w_1409));
  maj_bbi g370(.a(n337_4),.b(n369),.c(n368_0),.q(n370));
  bfr _b_1033(.a(_w_1589),.q(n282_2));
  or_bb g332(.a(in_48_),.b(in_49_),.q(n332));
  spl2 g159_s_0(.a(n159),.q0(n159_0),.q1(n159_1));
  or_bb g194(.a(in_68_),.b(in_69_),.q(n194));
  maj_bbi g375(.a(n308_3),.b(n314_3),.c(n317_3),.q(n375));
  maj_bbb g541(.a(n515_2),.b(n516_2),.c(n517_2),.q(_w_1460));
  or_bb g494(.a(n428_3),.b(n431_3),.q(n494));
  and_bi g299(.a(n298),.b(n297_0),.q(n299));
  or_bb g173(.a(in_92_),.b(in_93_),.q(_w_1405));
  spl2 g195_s_0(.a(n195),.q0(n195_0),.q1(n195_1));
  and_bb g383(.a(n344_3),.b(n382_0),.q(n383));
  spl2 g374_s_1(.a(n374_1),.q0(n374_2),.q1(n374_3));
  bfr _b_1182(.a(_w_1738),.q(_w_1739));
  bfr _b_929(.a(_w_1485),.q(_w_1486));
  spl3L g515_s_0(.a(n515),.q0(n515_0),.q1(n515_1),.q2(n515_2));
  spl3L g344_s_0(.a(n344),.q0(n344_0),.q1(n344_1),.q2(_w_1403));
  spl2 g197_s_0(.a(n197),.q0(n197_0),.q1(_w_1400));
  spl3L g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1),.q2(n294_2));
  spl3L g371_s_0(.a(n371),.q0(n371_0),.q1(n371_1),.q2(n371_2));
  bfr _b_984(.a(_w_1540),.q(_w_1541));
  spl2 g271_s_0(.a(n271),.q0(n271_0),.q1(_w_1397));
  spl2 g270_s_0(.a(n270),.q0(n270_0),.q1(n270_1));
  bfr _b_865(.a(_w_1421),.q(_w_1422));
  spl2 g208_s_0(.a(n208),.q0(n208_0),.q1(n208_1));
  spl3L g305_s_0(.a(n305),.q0(n305_0),.q1(n305_1),.q2(_w_1390));
  bfr _b_810(.a(_w_1366),.q(_w_1367));
  spl2 g181_s_0(.a(n181),.q0(n181_0),.q1(n181_1));
  spl2 g350_s_0(.a(n350),.q0(n350_0),.q1(_w_1703));
  bfr _b_1062(.a(_w_1618),.q(out_2_));
  spl3L g428_s_1(.a(n428_1),.q0(n428_2),.q1(n428_3),.q2(_w_1673));
  spl2 g307_s_0(.a(n307),.q0(n307_0),.q1(n307_1));
  spl2 g132_s_0(.a(n132),.q0(n132_0),.q1(n132_1));
  spl3L g206_s_0(.a(n206),.q0(n206_0),.q1(n206_1),.q2(n206_2));
  bfr _b_932(.a(_w_1488),.q(n170));
  spl3L g359_s_0(.a(n359),.q0(n359_0),.q1(n359_1),.q2(n359_2));
  spl2 g206_s_1(.a(n206_2),.q0(n206_3),.q1(_w_1389));
  bfr _b_992(.a(_w_1548),.q(_w_1549));
  spl3L g523_s_0(.a(n523),.q0(n523_0),.q1(n523_1),.q2(_w_1386));
  spl3L g245_s_0(.a(n245),.q0(n245_0),.q1(n245_1),.q2(n245_2));
  spl3L g529_s_0(.a(n529),.q0(n529_0),.q1(n529_1),.q2(n529_2));
  spl2 g216_s_0(.a(n216),.q0(n216_0),.q1(_w_1383));
  bfr _b_1005(.a(_w_1561),.q(n343));
  spl2 g216_s_1(.a(n216_1),.q0(n216_2),.q1(n216_3));
  spl2 g254_s_0(.a(n254),.q0(n254_0),.q1(n254_1));
  spl2 g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1));
  spl3L g243_s_0(.a(n243),.q0(n243_0),.q1(n243_1),.q2(n243_2));
  bfr _b_1035(.a(_w_1591),.q(n408));
  spl3L g251_s_0(.a(n251),.q0(n251_0),.q1(n251_1),.q2(n251_2));
  spl2 g481_s_0(.a(n481),.q0(n481_0),.q1(n481_1));
  spl3L g532_s_0(.a(n532),.q0(n532_0),.q1(n532_1),.q2(_w_1380));
  spl3L g257_s_0(.a(n257),.q0(n257_0),.q1(n257_1),.q2(n257_2));
  spl2 g259_s_0(.a(n259),.q0(n259_0),.q1(n259_1));
  spl3L g320_s_0(.a(n320),.q0(n320_0),.q1(n320_1),.q2(n320_2));
  spl2 g260_s_0(.a(n260),.q0(n260_0),.q1(n260_1));
  spl3L g261_s_0(.a(n261),.q0(n261_0),.q1(n261_1),.q2(_w_1378));
  bfr _b_1004(.a(_w_1560),.q(n346_3));
  spl3L g262_s_0(.a(n262),.q0(n262_0),.q1(n262_1),.q2(_w_1376));
  and_bb g169(.a(n148_0),.b(n168_0),.q(n169));
  spl2 g317_s_1(.a(n317_2),.q0(n317_3),.q1(_w_1375));
  bfr _b_883(.a(_w_1439),.q(n309));
  spl2 g264_s_0(.a(n264),.q0(n264_0),.q1(n264_1));
  and_bb g472(.a(n395_2),.b(n398_2),.q(n472));
  spl2 g265_s_0(.a(n265),.q0(n265_0),.q1(_w_1372));
  spl2 g265_s_1(.a(n265_1),.q0(n265_2),.q1(_w_1371));
  spl3L g499_s_0(.a(n499),.q0(n499_0),.q1(n499_1),.q2(_w_1368));
  spl2 g407_s_0(.a(n407),.q0(n407_0),.q1(n407_1));
  or_bb g253(.a(n233_1),.b(n251_1),.q(n253));
  spl2 g276_s_0(.a(n276),.q0(n276_0),.q1(n276_1));
  spl3L g233_s_0(.a(n233),.q0(n233_0),.q1(n233_1),.q2(n233_2));
  bfr _b_972(.a(_w_1528),.q(_w_1529));
  bfr _b_910(.a(_w_1466),.q(_w_1467));
  spl3L g281_s_0(.a(n281),.q0(n281_0),.q1(n281_1),.q2(_w_1366));
  and_bb g453(.a(n439_0),.b(n452_0),.q(n453));
  spl3L g277_s_0(.a(n277),.q0(n277_0),.q1(n277_1),.q2(n277_2));
  spl3L g268_s_0(.a(n268),.q0(n268_0),.q1(n268_1),.q2(_w_1364));
  spl3L g367_s_0(.a(n367),.q0(n367_0),.q1(n367_1),.q2(n367_2));
  or_bb g402(.a(n397_1),.b(n400_1),.q(n402));
  spl2 g535_s_0(.a(n535),.q0(n535_0),.q1(n535_1));
  bfr _b_788(.a(_w_1344),.q(n212_2));
  spl2 g285_s_0(.a(n285),.q0(n285_0),.q1(_w_1361));
  bfr _b_922(.a(_w_1478),.q(_w_1479));
  or_bb g372(.a(n340_2),.b(n370_1),.q(_w_1417));
  bfr _b_760(.a(_w_1316),.q(n491_2));
  bfr _b_924(.a(_w_1480),.q(n524));
  spl2 g285_s_1(.a(n285_1),.q0(n285_2),.q1(_w_1360));
  spl2 g211_s_0(.a(n211),.q0(n211_0),.q1(n211_1));
  spl2 g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1));
  spl2 g339_s_0(.a(n339),.q0(n339_0),.q1(n339_1));
  spl2 g299_s_0(.a(n299),.q0(n299_0),.q1(n299_1));
  and_bb g212(.a(n191_0),.b(n211_0),.q(n212));
  spl3L g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1),.q2(_w_1358));
  spl3L g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1),.q2(_w_1356));
  spl2 g306_s_0(.a(n306),.q0(n306_0),.q1(n306_1));
  spl2 g308_s_0(.a(n308),.q0(n308_0),.q1(_w_1353));
  spl2 g308_s_1(.a(n308_1),.q0(n308_2),.q1(_w_1352));
  bfr _b_1106(.a(_w_1662),.q(n275));
  spl2 g316_s_0(.a(n316),.q0(n316_0),.q1(n316_1));
  bfr _b_990(.a(_w_1546),.q(n338));
  bfr _b_963(.a(_w_1519),.q(_w_1520));
  spl3L g186_s_0(.a(n186),.q0(n186_0),.q1(n186_1),.q2(n186_2));
  bfr _b_959(.a(_w_1515),.q(_w_1516));
  and_bi g422(.a(n421),.b(n420),.q(n422));
  spl3L g331_s_0(.a(n331),.q0(n331_0),.q1(n331_1),.q2(_w_1349));
  spl2 g334_s_0(.a(n334),.q0(n334_0),.q1(_w_1346));
  spl2 g334_s_1(.a(n334_1),.q0(n334_2),.q1(_w_1345));
  spl3L g212_s_0(.a(n212),.q0(n212_0),.q1(n212_1),.q2(_w_1343));
  and_bi g513(.a(n512),.b(n511),.q(n513));
  spl3L g444_s_1(.a(n444_1),.q0(n444_2),.q1(n444_3),.q2(_w_1340));
  spl3L g340_s_0(.a(n340),.q0(n340_0),.q1(n340_1),.q2(n340_2));
  bfr _b_934(.a(_w_1490),.q(n167));
  spl2 g348_s_0(.a(n348),.q0(n348_0),.q1(n348_1));
  bfr _b_836(.a(_w_1392),.q(_w_1393));
  spl3L g446_s_0(.a(n446),.q0(n446_0),.q1(n446_1),.q2(n446_2));
  spl2 g376_s_0(.a(n376),.q0(n376_0),.q1(n376_1));
  or_bb g313(.a(in_40_),.b(in_41_),.q(n313));
  maj_bbi g156(.a(n151_2),.b(n154),.c(n155_0),.q(n156));
  spl2 g410_s_0(.a(n410),.q0(n410_0),.q1(n410_1));
  spl2 g364_s_0(.a(n364),.q0(n364_0),.q1(n364_1));
  spl3L g410_s_1(.a(n410_1),.q0(n410_2),.q1(n410_3),.q2(_w_1337));
  spl3L g354_s_0(.a(n354),.q0(n354_0),.q1(n354_1),.q2(n354_2));
  spl2 g248_s_0(.a(n248),.q0(n248_0),.q1(n248_1));
  spl3L g355_s_0(.a(n355),.q0(n355_0),.q1(n355_1),.q2(n355_2));
  spl2 g356_s_0(.a(n356),.q0(n356_0),.q1(_w_1334));
  bfr _b_1064(.a(_w_1620),.q(_w_1621));
  spl2 g356_s_1(.a(n356_1),.q0(n356_2),.q1(n356_3));
  maj_bbb g314(.a(n311_0),.b(n312_0),.c(n313_0),.q(n314));
  spl2 g345_s_0(.a(n345),.q0(n345_0),.q1(n345_1));
  spl3L g379_s_0(.a(n379),.q0(n379_0),.q1(n379_1),.q2(n379_2));
  bfr _b_871(.a(_w_1427),.q(n442));
  or_bb g347(.a(n302_1),.b(n345_1),.q(_w_1592));
  spl3L g237_s_0(.a(n237),.q0(n237_0),.q1(n237_1),.q2(n237_2));
  and_bb g500(.a(n441_2),.b(n444_2),.q(n500));
  spl2 g509_s_0(.a(n509),.q0(n509_0),.q1(n509_1));
  spl2 g177_s_0(.a(n177),.q0(n177_0),.q1(_w_1331));
  bfr _b_811(.a(_w_1367),.q(n281_2));
  bfr _b_826(.a(_w_1382),.q(n532_2));
  spl3L g513_s_0(.a(n513),.q0(n513_0),.q1(n513_1),.q2(_w_1328));
  bfr _b_844(.a(_w_1400),.q(_w_1401));
  spl3L g391_s_0(.a(n391),.q0(n391_0),.q1(n391_1),.q2(n391_2));
  spl3L g400_s_0(.a(n400),.q0(n400_0),.q1(n400_1),.q2(n400_2));
  spl3L g485_s_0(.a(n485),.q0(n485_0),.q1(n485_1),.q2(_w_1322));
  and_bb g157(.a(in_106_),.b(in_107_),.q(n157));
  spl3L g412_s_0(.a(n412),.q0(n412_0),.q1(n412_1),.q2(n412_2));
  and_bb g189(.a(n172_0),.b(n188_0),.q(n189));
  bfr _b_884(.a(_w_1440),.q(n432));
  spl3L g425_s_0(.a(n425),.q0(n425_0),.q1(n425_1),.q2(n425_2));
  spl2 g426_s_0(.a(n426),.q0(n426_0),.q1(_w_1320));
  bfr _b_862(.a(_w_1418),.q(_w_1419));
  and_bb g398(.a(n356_2),.b(n359_1),.q(n398));
  spl2 g426_s_1(.a(n426_1),.q0(n426_2),.q1(n426_3));
  spl3L g433_s_0(.a(n433),.q0(n433_0),.q1(n433_1),.q2(n433_2));
  spl3L g506_s_0(.a(n506),.q0(n506_0),.q1(n506_1),.q2(_w_1317));
  bfr _b_933(.a(_w_1489),.q(n539));
  bfr _b_848(.a(_w_1404),.q(n344_2));
  bfr _b_1006(.a(_w_1562),.q(n292));
  spl3L g491_s_0(.a(n491),.q0(n491_0),.q1(n491_1),.q2(_w_1314));
  maj_bbi g142(.a(n137_2),.b(n141),.c(n140_0),.q(n142));
  bfr _b_764(.a(_w_1320),.q(_w_1321));
  bfr _b_828(.a(_w_1384),.q(_w_1385));
  spl2 g234_s_0(.a(n234),.q0(n234_0),.q1(_w_1311));
  bfr _b_1143(.a(_w_1699),.q(_w_1700));
  and_bb g504(.a(n502_0),.b(n503_0),.q(n504));
  maj_bbi g319(.a(n304_2),.b(n318),.c(n317_0),.q(n319));
  spl3L g439_s_0(.a(n439),.q0(n439_0),.q1(n439_1),.q2(n439_2));
  bfr _b_1030(.a(_w_1586),.q(n323));
  spl2 g440_s_0(.a(n440),.q0(n440_0),.q1(_w_1309));
  spl3L g443_s_0(.a(n443),.q0(n443_0),.q1(n443_1),.q2(n443_2));
  bfr _b_771(.a(_w_1327),.q(n395_4));
  bfr _b_792(.a(_w_1348),.q(n334_1));
  spl2 g467_s_0(.a(n467),.q0(n467_0),.q1(n467_1));
  spl3L g516_s_0(.a(n516),.q0(n516_0),.q1(n516_1),.q2(_w_1306));
  spl2 g267_s_0(.a(n267),.q0(n267_0),.q1(n267_1));
  spl3L g482_s_0(.a(n482),.q0(n482_0),.q1(n482_1),.q2(n482_2));
  maj_bbb g271(.a(n268_0),.b(n269_0),.c(n270_0),.q(n271));
  spl3L g143_s_0(.a(n143),.q0(n143_0),.q1(n143_1),.q2(n143_2));
  spl2 g422_s_0(.a(n422),.q0(n422_0),.q1(n422_1));
  spl3L g503_s_0(.a(n503),.q0(n503_0),.q1(n503_1),.q2(n503_2));
  spl2 g398_s_0(.a(n398),.q0(n398_0),.q1(n398_1));
  or_bb g411(.a(n368_3),.b(n371_2),.q(_w_1595));
  bfr _b_825(.a(_w_1381),.q(_w_1382));
  spl3L g510_s_0(.a(n510),.q0(n510_0),.q1(n510_1),.q2(n510_2));
  bfr _b_782(.a(_w_1338),.q(_w_1339));
  spl3L g514_s_0(.a(n514),.q0(n514_0),.q1(n514_1),.q2(n514_2));
  spl2 g392_s_1(.a(n392_1),.q0(n392_2),.q1(n392_3));
  spl2 g415_s_0(.a(n415),.q0(n415_0),.q1(n415_1));
  maj_bbi g351(.a(n265_3),.b(n271_3),.c(n274_3),.q(n351));
  bfr _b_835(.a(_w_1391),.q(n305_2));
  spl3L g525_s_0(.a(n525),.q0(n525_0),.q1(n525_1),.q2(_w_1300));
  bfr _b_989(.a(_w_1545),.q(n244));
  bfr _b_744(.a(_w_1300),.q(_w_1301));
  bfr _b_745(.a(_w_1301),.q(_w_1302));
  bfr _b_746(.a(_w_1302),.q(n525_2));
  bfr _b_747(.a(_w_1303),.q(_w_1304));
  and_bi g348(.a(n347),.b(n346_0),.q(n348));
  and_bb g153(.a(in_98_),.b(in_99_),.q(n153));
  spl2 g224_s_0(.a(n224),.q0(n224_0),.q1(n224_1));
  bfr _b_876(.a(_w_1432),.q(n143_4));
  bfr _b_748(.a(_w_1304),.q(_w_1305));
  bfr _b_749(.a(_w_1305),.q(n478_2));
  bfr _b_939(.a(_w_1495),.q(_w_1496));
  bfr _b_750(.a(_w_1306),.q(_w_1307));
  and_bb g146(.a(n129_0),.b(n145_0),.q(n146));
  bfr _b_751(.a(_w_1307),.q(_w_1308));
  bfr _b_785(.a(_w_1341),.q(_w_1342));
  and_bb g450(.a(n440_2),.b(n449_0),.q(n450));
  bfr _b_815(.a(_w_1371),.q(n265_3));
  bfr _b_1055(.a(_w_1611),.q(_w_1612));
  bfr _b_752(.a(_w_1308),.q(n516_2));
  bfr _b_753(.a(_w_1309),.q(_w_1310));
  bfr _b_779(.a(_w_1335),.q(_w_1336));
  bfr _b_754(.a(_w_1310),.q(n440_1));
  bfr _b_755(.a(_w_1311),.q(_w_1312));
  bfr _b_756(.a(_w_1312),.q(_w_1313));
  bfr _b_762(.a(_w_1318),.q(_w_1319));
  bfr _b_763(.a(_w_1319),.q(n506_2));
  bfr _b_765(.a(_w_1321),.q(n426_1));
  bfr _b_766(.a(_w_1322),.q(_w_1323));
  spl2 g300_s_1(.a(n300_2),.q0(n300_3),.q1(n300_4));
  bfr _b_896(.a(_w_1452),.q(_w_1453));
  and_bb g462(.a(n392_2),.b(n461_0),.q(n462));
  bfr _b_773(.a(_w_1329),.q(_w_1330));
  bfr _b_817(.a(_w_1373),.q(_w_1374));
  bfr _b_1009(.a(_w_1565),.q(n137_2));
  maj_bbi g145(.a(n130_2),.b(n144),.c(n143_0),.q(n145));
  bfr _b_774(.a(_w_1330),.q(n513_2));
  bfr _b_775(.a(_w_1331),.q(_w_1332));
  bfr _b_852(.a(_w_1408),.q(n173));
  bfr _b_776(.a(_w_1332),.q(_w_1333));
  bfr _b_1016(.a(_w_1572),.q(_w_1573));
  bfr _b_777(.a(_w_1333),.q(n177_1));
  bfr _b_784(.a(_w_1340),.q(_w_1341));
  and_bb g401(.a(n397_0),.b(n400_0),.q(n401));
  bfr _b_786(.a(_w_1342),.q(n444_4));
  and_bb g215(.a(n171_0),.b(n214_0),.q(n215));
  bfr _b_790(.a(_w_1346),.q(_w_1347));
  bfr _b_793(.a(_w_1349),.q(_w_1350));
  bfr _b_796(.a(_w_1352),.q(n308_3));
  and_bb g386(.a(n367_0),.b(n385_0),.q(n386));
  spl3L g409_s_0(.a(n409),.q0(n409_0),.q1(n409_1),.q2(n409_2));
  bfr _b_798(.a(_w_1354),.q(_w_1355));
  bfr _b_799(.a(_w_1355),.q(n308_1));
  spl2 g139_s_0(.a(n139),.q0(n139_0),.q1(n139_1));
  bfr _b_947(.a(_w_1503),.q(_w_1504));
  bfr _b_977(.a(_w_1533),.q(n144));
  bfr _b_1026(.a(_w_1582),.q(_w_1583));
  bfr _b_800(.a(_w_1356),.q(_w_1357));
  bfr _b_802(.a(_w_1358),.q(_w_1359));
  bfr _b_952(.a(_w_1508),.q(_w_1509));
  bfr _b_804(.a(_w_1360),.q(n285_3));
  bfr _b_806(.a(_w_1362),.q(_w_1363));
  maj_bbi g136(.a(n131_2),.b(n135),.c(n134_0),.q(n136));
  bfr _b_808(.a(_w_1364),.q(_w_1365));
  bfr _b_812(.a(_w_1368),.q(_w_1369));
  bfr _b_821(.a(_w_1377),.q(n262_2));
  bfr _b_823(.a(_w_1379),.q(n261_2));
  bfr _b_827(.a(_w_1383),.q(_w_1384));
  bfr _b_953(.a(_w_1509),.q(_w_1510));
  bfr _b_830(.a(_w_1386),.q(_w_1387));
  bfr _b_935(.a(_w_1491),.q(_w_1492));
  bfr _b_831(.a(_w_1387),.q(_w_1388));
  bfr _b_832(.a(_w_1388),.q(n523_2));
  bfr _b_834(.a(_w_1390),.q(_w_1391));
  bfr _b_837(.a(_w_1393),.q(n416_1));
  bfr _b_846(.a(_w_1402),.q(n197_1));
  bfr _b_968(.a(_w_1524),.q(_w_1525));
  bfr _b_839(.a(_w_1395),.q(n393_1));
  bfr _b_841(.a(_w_1397),.q(_w_1398));
  bfr _b_842(.a(_w_1398),.q(_w_1399));
  bfr _b_843(.a(_w_1399),.q(n271_1));
  spl3L g151_s_0(.a(n151),.q0(n151_0),.q1(n151_1),.q2(_w_1701));
  bfr _b_845(.a(_w_1401),.q(_w_1402));
  and_bb g181(.a(in_86_),.b(in_87_),.q(n181));
  bfr _b_847(.a(_w_1403),.q(_w_1404));
  bfr _b_850(.a(_w_1406),.q(_w_1407));
  bfr _b_851(.a(_w_1407),.q(_w_1408));
  bfr _b_1041(.a(_w_1597),.q(_w_1598));
  bfr _b_854(.a(_w_1410),.q(_w_1411));
  spl2 g328_s_1(.a(n328_1),.q0(n328_2),.q1(_w_1351));
  bfr _b_857(.a(_w_1413),.q(n169_2));
  bfr _b_860(.a(_w_1416),.q(n349_1));
  bfr _b_866(.a(_w_1422),.q(_w_1423));
  bfr _b_868(.a(_w_1424),.q(n238));
  maj_bbi g293(.a(n288_2),.b(n292),.c(n291_0),.q(n293));
  bfr _b_869(.a(_w_1425),.q(n163_4));
  bfr _b_872(.a(_w_1428),.q(_w_1429));
  spl3L g441_s_1(.a(n441_1),.q0(n441_2),.q1(n441_3),.q2(_w_1631));
  bfr _b_877(.a(_w_1433),.q(_w_1434));
  bfr _b_878(.a(_w_1434),.q(n173_2));
  bfr _b_879(.a(_w_1435),.q(n186_4));
  bfr _b_885(.a(_w_1441),.q(n353));
  bfr _b_886(.a(_w_1442),.q(_w_1443));
  bfr _b_887(.a(_w_1443),.q(n194_2));
  bfr _b_888(.a(_w_1444),.q(_w_1445));
  bfr _b_1031(.a(_w_1587),.q(n360));
  maj_bbb g416(.a(n344_1),.b(n373_2),.c(n379_2),.q(n416));
  bfr _b_892(.a(_w_1448),.q(_w_1449));
  bfr _b_925(.a(_w_1481),.q(_w_1482));
  bfr _b_1003(.a(_w_1559),.q(_w_1560));
  bfr _b_893(.a(_w_1449),.q(n311_2));
  spl2 g416_s_0(.a(n416),.q0(n416_0),.q1(_w_1392));
  spl2 g322_s_0(.a(n322),.q0(n322_0),.q1(n322_1));
  spl3L g395_s_1(.a(n395_1),.q0(n395_2),.q1(n395_3),.q2(_w_1325));
  bfr _b_894(.a(_w_1450),.q(n335));
  bfr _b_895(.a(_w_1451),.q(_w_1452));
  bfr _b_897(.a(_w_1453),.q(_w_1454));
  and_bb g180(.a(in_90_),.b(in_91_),.q(n180));
  or_bb g451(.a(n440_3),.b(n449_1),.q(n451));
  bfr _b_899(.a(_w_1455),.q(_w_1456));
  bfr _b_901(.a(_w_1457),.q(_w_1458));
  bfr _b_902(.a(_w_1458),.q(n280));
  bfr _b_903(.a(_w_1459),.q(n278));
  bfr _b_906(.a(_w_1462),.q(n541));
  spl3L g193_s_0(.a(n193),.q0(n193_0),.q1(n193_1),.q2(_w_1620));
  spl2 g349_s_0(.a(n349),.q0(n349_0),.q1(_w_1414));
  bfr _b_907(.a(_w_1463),.q(n298));
  bfr _b_908(.a(_w_1464),.q(n315));
  and_bi g227(.a(n226),.b(n225_0),.q(n227));
  bfr _b_1100(.a(_w_1656),.q(out_1_));
  spl2 g441_s_0(.a(n441),.q0(n441_0),.q1(n441_1));
  bfr _b_889(.a(_w_1445),.q(_w_1446));
  bfr _b_909(.a(_w_1465),.q(_w_1466));
  bfr _b_1105(.a(_w_1661),.q(n341));
  bfr _b_911(.a(_w_1467),.q(_w_1468));
  maj_bbi g266(.a(n263_1),.b(n264_1),.c(n262_1),.q(_w_1722));
  bfr _b_913(.a(_w_1469),.q(_w_1470));
  bfr _b_916(.a(_w_1472),.q(n260));
  bfr _b_919(.a(_w_1475),.q(_w_1476));
  bfr _b_920(.a(_w_1476),.q(n324_2));
  and_bi g279(.a(n278),.b(n277_0),.q(n279));
  spl2 g319_s_0(.a(n319),.q0(n319_0),.q1(n319_1));
  bfr _b_921(.a(_w_1477),.q(n178));
  bfr _b_923(.a(_w_1479),.q(_w_1480));
  bfr _b_930(.a(_w_1486),.q(_w_1487));
  and_bb g323(.a(in_62_),.b(in_63_),.q(_w_1579));
  bfr _b_931(.a(_w_1487),.q(n291_1));
  spl2 g289_s_0(.a(n289),.q0(n289_0),.q1(n289_1));
  bfr _b_937(.a(_w_1493),.q(n407_4));
  bfr _b_941(.a(_w_1497),.q(_w_1498));
  or_bb g301(.a(n279_1),.b(n299_1),.q(_w_1420));
  bfr _b_943(.a(_w_1499),.q(_w_1500));
  and_bi g239(.a(n238),.b(n237_0),.q(n239));
  bfr _b_1017(.a(_w_1573),.q(n304));
  spl3L g478_s_0(.a(n478),.q0(n478_0),.q1(n478_1),.q2(_w_1303));
  bfr _b_946(.a(_w_1502),.q(n303));
  spl2 g382_s_0(.a(n382),.q0(n382_0),.q1(n382_1));
  bfr _b_948(.a(_w_1504),.q(n200_2));
  spl2 g436_s_0(.a(n436),.q0(n436_0),.q1(n436_1));
  bfr _b_949(.a(_w_1505),.q(n445));
  spl2 g177_s_1(.a(n177_1),.q0(n177_2),.q1(_w_1641));
  bfr _b_950(.a(_w_1506),.q(_w_1507));
  bfr _b_973(.a(_w_1529),.q(_w_1530));
  spl2 g136_s_0(.a(n136),.q0(n136_0),.q1(n136_1));
  bfr _b_955(.a(_w_1511),.q(_w_1512));
  or_bb g463(.a(n392_3),.b(n461_1),.q(n463));
  bfr _b_761(.a(_w_1317),.q(_w_1318));
  bfr _b_975(.a(_w_1531),.q(n164));
  bfr _b_1015(.a(_w_1571),.q(_w_1572));
  bfr _b_956(.a(_w_1512),.q(_w_1513));
  spl2 g393_s_0(.a(n393),.q0(n393_0),.q1(_w_1394));
  bfr _b_958(.a(_w_1514),.q(_w_1515));
  spl2 g271_s_1(.a(n271_1),.q0(n271_2),.q1(_w_1396));
  bfr _b_960(.a(_w_1516),.q(n543));
  bfr _b_961(.a(_w_1517),.q(n135));
  spl2 g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1));
  bfr _b_962(.a(_w_1518),.q(n161));
  bfr _b_965(.a(_w_1521),.q(n517));
  bfr _b_971(.a(_w_1527),.q(_w_1528));
  maj_bbi g205(.a(n200_2),.b(n204),.c(n203_0),.q(n205));
  bfr _b_966(.a(_w_1522),.q(n286));
  spl2 g374_s_0(.a(n374),.q0(n374_0),.q1(_w_1737));
  bfr _b_969(.a(_w_1525),.q(_w_1526));
  bfr _b_976(.a(_w_1532),.q(n141));
  bfr _b_979(.a(_w_1535),.q(_w_1536));
  bfr _b_980(.a(_w_1536),.q(n288_2));
  spl3L g419_s_0(.a(n419),.q0(n419_0),.q1(n419_1),.q2(n419_2));
  bfr _b_982(.a(_w_1538),.q(_w_1539));
  spl2 g183_s_0(.a(n183),.q0(n183_0),.q1(_w_1685));
  and_bb g362(.a(n355_0),.b(n361_0),.q(n362));
  spl3L g471_s_0(.a(n471),.q0(n471_0),.q1(n471_1),.q2(n471_2));
  bfr _b_985(.a(_w_1541),.q(_w_1542));
  bfr _b_987(.a(_w_1543),.q(_w_1544));
  bfr _b_988(.a(_w_1544),.q(n149));
  spl2 g444_s_0(.a(n444),.q0(n444_0),.q1(n444_1));
  bfr _b_840(.a(_w_1396),.q(n271_3));
  bfr _b_991(.a(_w_1547),.q(_w_1548));
  bfr _b_993(.a(_w_1549),.q(_w_1550));
  spl2 g332_s_0(.a(n332),.q0(n332_0),.q1(n332_1));
  bfr _b_1001(.a(_w_1557),.q(n134_3));
  bfr _b_994(.a(_w_1550),.q(_w_1551));
  bfr _b_995(.a(_w_1551),.q(_w_1552));
  bfr _b_996(.a(_w_1552),.q(_w_1553));
  bfr _b_997(.a(_w_1553),.q(_w_1554));
  bfr _b_1002(.a(_w_1558),.q(n198));
  bfr _b_1007(.a(_w_1563),.q(n154));
  bfr _b_1008(.a(_w_1564),.q(_w_1565));
  bfr _b_1010(.a(_w_1566),.q(n226));
  bfr _b_986(.a(_w_1542),.q(_w_1543));
  bfr _b_1011(.a(_w_1567),.q(n204));
  bfr _b_1012(.a(_w_1568),.q(n258));
  bfr _b_1013(.a(_w_1569),.q(n272));
  and_bb g486(.a(n478_0),.b(n485_0),.q(n486));
  bfr _b_1014(.a(_w_1570),.q(_w_1571));
  bfr _b_1019(.a(_w_1575),.q(n210));
  bfr _b_1020(.a(_w_1576),.q(n294_4));
  bfr _b_1021(.a(_w_1577),.q(n183_3));
  bfr _b_1054(.a(_w_1610),.q(n184));
  or_bb g159(.a(in_104_),.b(in_105_),.q(n159));
  bfr _b_1022(.a(_w_1578),.q(n213));
  and_bb g284(.a(in_2_),.b(in_3_),.q(n284));
  bfr _b_1032(.a(_w_1588),.q(_w_1589));
  bfr _b_1034(.a(_w_1590),.q(n220));
  bfr _b_1036(.a(_w_1592),.q(n347));
  bfr _b_1038(.a(_w_1594),.q(n150_2));
  bfr _b_1042(.a(_w_1598),.q(_w_1599));
  bfr _b_1043(.a(_w_1599),.q(n261));
  spl2 g349_s_1(.a(n349_1),.q0(n349_2),.q1(_w_1437));
  bfr _b_1044(.a(_w_1600),.q(_w_1601));
  bfr _b_1046(.a(_w_1602),.q(n155_1));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(n280_1));
  bfr _b_1048(.a(_w_1604),.q(_w_1605));
  bfr _b_822(.a(_w_1378),.q(_w_1379));
  bfr _b_1050(.a(_w_1606),.q(n525));
  bfr _b_1052(.a(_w_1608),.q(n147));
  or_bb g139(.a(in_120_),.b(in_121_),.q(n139));
  bfr _b_954(.a(_w_1510),.q(_w_1511));
  bfr _b_936(.a(_w_1492),.q(_w_1493));
  bfr _b_1053(.a(_w_1609),.q(n190));
  spl3L g150_s_0(.a(n150),.q0(n150_0),.q1(n150_1),.q2(_w_1593));
  and_bb g133(.a(in_114_),.b(in_115_),.q(n133));
  spl3L g288_s_0(.a(n288),.q0(n288_0),.q1(n288_1),.q2(_w_1535));
  bfr _b_1057(.a(_w_1613),.q(out_3_));
  bfr _b_1058(.a(_w_1614),.q(_w_1615));
  bfr _b_1059(.a(_w_1615),.q(_w_1616));
  bfr _b_1060(.a(_w_1616),.q(_w_1617));
  bfr _b_1065(.a(_w_1621),.q(n193_2));
  bfr _b_978(.a(_w_1534),.q(n318));
  bfr _b_1107(.a(_w_1663),.q(_w_1664));
  bfr _b_1066(.a(_w_1622),.q(_w_1623));
  bfr _b_1070(.a(_w_1626),.q(_w_1627));
  bfr _b_1071(.a(_w_1627),.q(_w_1628));
  bfr _b_1074(.a(_w_1630),.q(n140_3));
  bfr _b_1077(.a(_w_1633),.q(n441_4));
  bfr _b_881(.a(_w_1437),.q(_w_1438));
  bfr _b_1080(.a(_w_1636),.q(_w_1637));
  bfr _b_1081(.a(_w_1637),.q(n203_1));
  bfr _b_1149(.a(_w_1705),.q(n350_1));
  bfr _b_1086(.a(_w_1642),.q(_w_1643));
  bfr _b_1088(.a(_w_1644),.q(_w_1645));
  bfr _b_805(.a(_w_1361),.q(_w_1362));
  spl2 g352_s_0(.a(n352),.q0(n352_0),.q1(n352_1));
  bfr _b_1089(.a(_w_1645),.q(_w_1646));
  bfr _b_1090(.a(_w_1646),.q(_w_1647));
  bfr _b_1094(.a(_w_1650),.q(_w_1651));
  bfr _b_1096(.a(_w_1652),.q(_w_1653));
  bfr _b_1097(.a(_w_1653),.q(_w_1654));
  bfr _b_1098(.a(_w_1654),.q(_w_1655));
  bfr _b_1099(.a(_w_1655),.q(_w_1656));
  bfr _b_1101(.a(_w_1657),.q(_w_1658));
  bfr _b_1104(.a(_w_1660),.q(out_4_));
  assign out_0_ = 1'b0;
endmodule
