module c5315( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G158 , G159 , G16 , G160 , G161 , G162 , G163 , G164 , G165 , G166 , G167 , G168 , G169 , G17 , G170 , G171 , G172 , G173 , G174 , G175 , G176 , G177 , G178 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G5193 , G5194 , G5195 , G5196 , G5197 , G5198 , G5199 , G5200 , G5201 , G5202 , G5203 , G5204 , G5205 , G5206 , G5207 , G5208 , G5209 , G5210 , G5211 , G5212 , G5213 , G5214 , G5215 , G5216 , G5217 , G5218 , G5219 , G5220 , G5221 , G5222 , G5223 , G5224 , G5225 , G5226 , G5227 , G5228 , G5229 , G5230 , G5231 , G5232 , G5233 , G5234 , G5235 , G5236 , G5237 , G5238 , G5239 , G5240 , G5241 , G5242 , G5243 , G5244 , G5245 , G5246 , G5247 , G5248 , G5249 , G5250 , G5251 , G5252 , G5253 , G5254 , G5255 , G5256 , G5257 , G5258 , G5259 , G5260 , G5261 , G5262 , G5263 , G5264 , G5265 , G5266 , G5267 , G5268 , G5269 , G5270 , G5271 , G5272 , G5273 , G5274 , G5275 , G5276 , G5277 , G5278 , G5279 , G5280 , G5281 , G5282 , G5283 , G5284 , G5285 , G5286 , G5287 , G5288 , G5289 , G5290 , G5291 , G5292 , G5293 , G5294 , G5295 , G5296 , G5297 , G5298 , G5299 , G5300 , G5301 , G5302 , G5303 , G5304 , G5305 , G5306 , G5307 , G5308 , G5309 , G5310 , G5311 , G5312 , G5313 , G5314 , G5315 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 ;
  assign n179 = G153 & G156 ;
  assign n180 = G66 & G67 ;
  assign n181 = G1 & G134 ;
  assign n182 = ~G165 & G63 ;
  assign n183 = ~G11 | G164 ;
  assign n184 = ~G136 | ~G154 ;
  assign n185 = ~G11 | ~G12 ;
  assign n186 = ~G65 | ~n185 ;
  assign n187 = G163 & G34 ;
  assign n188 = ~G163 & G33 ;
  assign n189 = n187 | n188 ;
  assign n190 = ~n185 | ~n189 ;
  assign n191 = G13 & G163 ;
  assign n192 = ~G163 & G35 ;
  assign n193 = n191 | n192 ;
  assign n194 = ~n185 | ~n193 ;
  assign n195 = ~G32 | ~n185 ;
  assign n196 = ~G163 & G9 ;
  assign n197 = G163 & G8 ;
  assign n198 = n185 & ~n197 ;
  assign n199 = ~n196 & n198 ;
  assign n200 = G66 & ~n199 ;
  assign n201 = ~G163 & G30 ;
  assign n202 = G10 & G163 ;
  assign n203 = n185 & ~n202 ;
  assign n204 = ~n201 & n203 ;
  assign n205 = G66 & ~n204 ;
  assign n206 = ~G163 & G7 ;
  assign n207 = G163 & G28 ;
  assign n208 = n185 & ~n207 ;
  assign n209 = ~n206 & n208 ;
  assign n210 = G66 & ~n209 ;
  assign n211 = ~G163 & G29 ;
  assign n212 = G163 & G31 ;
  assign n213 = n185 & ~n212 ;
  assign n214 = ~n211 & n213 ;
  assign n215 = G66 & ~n214 ;
  assign n216 = G100 | G117 ;
  assign n217 = ~G101 & G117 ;
  assign n218 = n216 & ~n217 ;
  assign n219 = G145 & ~n218 ;
  assign n220 = G102 & G117 ;
  assign n221 = ~G117 & G98 ;
  assign n222 = n220 | n221 ;
  assign n223 = ~G145 & n222 ;
  assign n224 = n219 | n223 ;
  assign n225 = G100 | G119 ;
  assign n226 = ~G101 & G119 ;
  assign n227 = n225 & ~n226 ;
  assign n228 = G146 & ~n227 ;
  assign n229 = G102 & G119 ;
  assign n230 = ~G119 & G98 ;
  assign n231 = n229 | n230 ;
  assign n232 = ~G146 & n231 ;
  assign n233 = n228 | n232 ;
  assign n234 = n224 & n233 ;
  assign n235 = G128 | G169 ;
  assign n236 = G128 & ~G168 ;
  assign n237 = n235 & ~n236 ;
  assign n238 = G150 & ~n237 ;
  assign n239 = G128 & G167 ;
  assign n240 = ~G128 & G166 ;
  assign n241 = n239 | n240 ;
  assign n242 = ~G150 & n241 ;
  assign n243 = n238 | n242 ;
  assign n244 = G113 | G98 ;
  assign n245 = ~G102 & G113 ;
  assign n246 = n244 & ~n245 ;
  assign n247 = G100 | G115 ;
  assign n248 = ~G101 & G115 ;
  assign n249 = n247 & ~n248 ;
  assign n250 = n246 & ~n249 ;
  assign n251 = G100 | G130 ;
  assign n252 = ~G101 & G130 ;
  assign n253 = n251 & ~n252 ;
  assign n254 = ~G148 & G166 ;
  assign n255 = G148 & ~G169 ;
  assign n256 = n254 | n255 ;
  assign n257 = ~n253 & n256 ;
  assign n258 = n250 & n257 ;
  assign n259 = n243 & n258 ;
  assign n260 = G121 | G169 ;
  assign n261 = G121 & ~G168 ;
  assign n262 = n260 & ~n261 ;
  assign n263 = G147 & ~n262 ;
  assign n264 = G121 & G167 ;
  assign n265 = ~G121 & G166 ;
  assign n266 = n264 | n265 ;
  assign n267 = ~G147 & n266 ;
  assign n268 = n263 | n267 ;
  assign n269 = G126 | G169 ;
  assign n270 = G126 & ~G168 ;
  assign n271 = n269 & ~n270 ;
  assign n272 = G149 & ~n271 ;
  assign n273 = G126 & G167 ;
  assign n274 = ~G126 & G166 ;
  assign n275 = n273 | n274 ;
  assign n276 = ~G149 & n275 ;
  assign n277 = n272 | n276 ;
  assign n278 = n268 & n277 ;
  assign n279 = n259 & n278 ;
  assign n280 = n234 & n279 ;
  assign n281 = G169 | G94 ;
  assign n282 = ~G168 & G94 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = G140 & ~n283 ;
  assign n285 = G167 & G94 ;
  assign n286 = G166 & ~G94 ;
  assign n287 = n285 | n286 ;
  assign n288 = ~G140 & n287 ;
  assign n289 = n284 | n288 ;
  assign n290 = G169 | G90 ;
  assign n291 = ~G168 & G90 ;
  assign n292 = n290 & ~n291 ;
  assign n293 = G143 & ~n292 ;
  assign n294 = G167 & G90 ;
  assign n295 = G166 & ~G90 ;
  assign n296 = n294 | n295 ;
  assign n297 = ~G143 & n296 ;
  assign n298 = n293 | n297 ;
  assign n299 = G169 | G92 ;
  assign n300 = ~G168 & G92 ;
  assign n301 = n299 & ~n300 ;
  assign n302 = G144 & ~n301 ;
  assign n303 = G167 & G92 ;
  assign n304 = G166 & ~G92 ;
  assign n305 = n303 | n304 ;
  assign n306 = ~G144 & n305 ;
  assign n307 = n302 | n306 ;
  assign n308 = n298 & n307 ;
  assign n309 = n289 & n308 ;
  assign n310 = G109 | G169 ;
  assign n311 = G109 & ~G168 ;
  assign n312 = n310 & ~n311 ;
  assign n313 = G135 & ~n312 ;
  assign n314 = G109 & G167 ;
  assign n315 = ~G109 & G166 ;
  assign n316 = n314 | n315 ;
  assign n317 = ~G135 & n316 ;
  assign n318 = n313 | n317 ;
  assign n319 = G169 | G96 ;
  assign n320 = ~G168 & G96 ;
  assign n321 = n319 & ~n320 ;
  assign n322 = G141 & ~n321 ;
  assign n323 = G167 & G96 ;
  assign n324 = G166 & ~G96 ;
  assign n325 = n323 | n324 ;
  assign n326 = ~G141 & n325 ;
  assign n327 = n322 | n326 ;
  assign n328 = n318 & n327 ;
  assign n329 = G107 | G169 ;
  assign n330 = G107 & ~G168 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = G139 & ~n331 ;
  assign n333 = G107 & G167 ;
  assign n334 = ~G107 & G166 ;
  assign n335 = n333 | n334 ;
  assign n336 = ~G139 & n335 ;
  assign n337 = n332 | n336 ;
  assign n338 = G101 | G88 ;
  assign n339 = ~G100 & G88 ;
  assign n340 = n338 & ~n339 ;
  assign n341 = G142 & ~n340 ;
  assign n342 = G88 & G98 ;
  assign n343 = G102 & ~G88 ;
  assign n344 = n342 | n343 ;
  assign n345 = ~G142 & n344 ;
  assign n346 = n341 | n345 ;
  assign n347 = n337 & n346 ;
  assign n348 = G103 | G169 ;
  assign n349 = G103 & ~G168 ;
  assign n350 = n348 & ~n349 ;
  assign n351 = G137 & ~n350 ;
  assign n352 = G103 & G167 ;
  assign n353 = ~G103 & G166 ;
  assign n354 = n352 | n353 ;
  assign n355 = ~G137 & n354 ;
  assign n356 = n351 | n355 ;
  assign n357 = G105 | G169 ;
  assign n358 = G105 & ~G168 ;
  assign n359 = n357 & ~n358 ;
  assign n360 = G138 & ~n359 ;
  assign n361 = G105 & G167 ;
  assign n362 = ~G105 & G166 ;
  assign n363 = n361 | n362 ;
  assign n364 = ~G138 & n363 ;
  assign n365 = n360 | n364 ;
  assign n366 = n356 & n365 ;
  assign n367 = n347 & n366 ;
  assign n368 = n328 & n367 ;
  assign n369 = n309 & n368 ;
  assign n370 = G124 & G96 ;
  assign n371 = ~G124 & G97 ;
  assign n372 = n370 | n371 ;
  assign n373 = G141 & n372 ;
  assign n374 = G141 | n372 ;
  assign n375 = ~n373 & n374 ;
  assign n376 = G109 & G124 ;
  assign n377 = G110 & ~G124 ;
  assign n378 = n376 | n377 ;
  assign n379 = G135 & n378 ;
  assign n380 = G135 | n378 ;
  assign n381 = ~n379 & n380 ;
  assign n382 = G107 & G124 ;
  assign n383 = G108 & ~G124 ;
  assign n384 = n382 | n383 ;
  assign n385 = G139 | n384 ;
  assign n386 = G139 & n384 ;
  assign n387 = n385 & ~n386 ;
  assign n388 = n381 & n387 ;
  assign n389 = G105 & G124 ;
  assign n390 = G106 & ~G124 ;
  assign n391 = n389 | n390 ;
  assign n392 = G138 & n391 ;
  assign n393 = G138 | n391 ;
  assign n394 = ~n392 & n393 ;
  assign n395 = G103 & G124 ;
  assign n396 = G104 & ~G124 ;
  assign n397 = n395 | n396 ;
  assign n398 = G137 | n397 ;
  assign n399 = G137 & n397 ;
  assign n400 = n398 & ~n399 ;
  assign n401 = n394 & n400 ;
  assign n402 = n388 & n401 ;
  assign n403 = n375 & n402 ;
  assign n404 = G124 & G88 ;
  assign n405 = ~G124 & G89 ;
  assign n406 = n404 | n405 ;
  assign n407 = G142 & n406 ;
  assign n408 = G142 | n406 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = G124 & G90 ;
  assign n411 = ~G124 & G91 ;
  assign n412 = n410 | n411 ;
  assign n413 = G143 & n412 ;
  assign n414 = G143 | n412 ;
  assign n415 = ~n413 & n414 ;
  assign n416 = G124 & G92 ;
  assign n417 = ~G124 & G93 ;
  assign n418 = n416 | n417 ;
  assign n419 = G144 & n418 ;
  assign n420 = G144 | n418 ;
  assign n421 = ~n419 & n420 ;
  assign n422 = G124 & G94 ;
  assign n423 = ~G124 & G95 ;
  assign n424 = n422 | n423 ;
  assign n425 = G140 & n424 ;
  assign n426 = G140 | n424 ;
  assign n427 = ~n425 & n426 ;
  assign n428 = n421 & n427 ;
  assign n429 = n415 & n428 ;
  assign n430 = n409 & n429 ;
  assign n431 = n403 & n430 ;
  assign n432 = G123 | G125 ;
  assign n433 = G148 & n432 ;
  assign n434 = G148 | n432 ;
  assign n435 = ~n433 & n434 ;
  assign n436 = G123 & G128 ;
  assign n437 = ~G123 & G129 ;
  assign n438 = n436 | n437 ;
  assign n439 = G150 | n438 ;
  assign n440 = G123 & G130 ;
  assign n441 = ~G123 & G131 ;
  assign n442 = n440 | n441 ;
  assign n443 = G150 & n438 ;
  assign n444 = n442 | n443 ;
  assign n445 = n439 & ~n444 ;
  assign n446 = G123 & G126 ;
  assign n447 = ~G123 & G127 ;
  assign n448 = n446 | n447 ;
  assign n449 = G149 & n448 ;
  assign n450 = G149 | n448 ;
  assign n451 = ~n449 & n450 ;
  assign n452 = n445 & n451 ;
  assign n453 = n435 & n452 ;
  assign n454 = G117 & G123 ;
  assign n455 = G118 & ~G123 ;
  assign n456 = n454 | n455 ;
  assign n457 = G145 & n456 ;
  assign n458 = G145 | n456 ;
  assign n459 = ~n457 & n458 ;
  assign n460 = G119 & G123 ;
  assign n461 = G120 & ~G123 ;
  assign n462 = n460 | n461 ;
  assign n463 = G146 & n462 ;
  assign n464 = G146 | n462 ;
  assign n465 = ~n463 & n464 ;
  assign n466 = n459 & n465 ;
  assign n467 = G113 & G123 ;
  assign n468 = G114 & ~G123 ;
  assign n469 = n467 | n468 ;
  assign n470 = G115 & G123 ;
  assign n471 = G116 & ~G123 ;
  assign n472 = n470 | n471 ;
  assign n473 = n469 | n472 ;
  assign n474 = G122 | G123 ;
  assign n475 = ~G121 & G123 ;
  assign n476 = n474 & ~n475 ;
  assign n477 = G147 & n476 ;
  assign n478 = G147 | n476 ;
  assign n479 = ~n477 & n478 ;
  assign n480 = ~n473 & n479 ;
  assign n481 = n466 & n480 ;
  assign n482 = n453 & n481 ;
  assign n483 = G113 | G115 ;
  assign n484 = G113 & G115 ;
  assign n485 = n483 & ~n484 ;
  assign n486 = G117 & ~G119 ;
  assign n487 = ~G117 & G119 ;
  assign n488 = n486 | n487 ;
  assign n489 = ~n485 & n488 ;
  assign n490 = n485 & ~n488 ;
  assign n491 = n489 | n490 ;
  assign n492 = G130 & ~G132 ;
  assign n493 = ~G130 & G132 ;
  assign n494 = n492 | n493 ;
  assign n495 = G121 & ~n494 ;
  assign n496 = ~G121 & n494 ;
  assign n497 = n495 | n496 ;
  assign n498 = G126 & ~G128 ;
  assign n499 = ~G126 & G128 ;
  assign n500 = n498 | n499 ;
  assign n501 = n497 & ~n500 ;
  assign n502 = ~n497 & n500 ;
  assign n503 = n501 | n502 ;
  assign n504 = n491 | n503 ;
  assign n505 = n491 & n503 ;
  assign n506 = ~n504 | n505 ;
  assign n507 = G88 | G90 ;
  assign n508 = G88 & G90 ;
  assign n509 = n507 & ~n508 ;
  assign n510 = G92 & ~G94 ;
  assign n511 = ~G92 & G94 ;
  assign n512 = n510 | n511 ;
  assign n513 = ~n509 & n512 ;
  assign n514 = n509 & ~n512 ;
  assign n515 = n513 | n514 ;
  assign n516 = G103 | G96 ;
  assign n517 = G103 & G96 ;
  assign n518 = n516 & ~n517 ;
  assign n519 = G109 & ~G111 ;
  assign n520 = ~G109 & G111 ;
  assign n521 = n519 | n520 ;
  assign n522 = n518 | n521 ;
  assign n523 = n518 & n521 ;
  assign n524 = n522 & ~n523 ;
  assign n525 = G105 & ~G107 ;
  assign n526 = ~G105 & G107 ;
  assign n527 = n525 | n526 ;
  assign n528 = n524 & ~n527 ;
  assign n529 = ~n524 & n527 ;
  assign n530 = n528 | n529 ;
  assign n531 = n515 & n530 ;
  assign n532 = n515 | n530 ;
  assign n533 = n531 | ~n532 ;
  assign n534 = n379 & n385 ;
  assign n535 = n386 | n392 ;
  assign n536 = n534 | n535 ;
  assign n537 = n393 & n536 ;
  assign n538 = n375 & n400 ;
  assign n539 = n537 & n538 ;
  assign n540 = n374 & n399 ;
  assign n541 = n373 | n540 ;
  assign n542 = n539 | n541 ;
  assign n543 = n430 & n542 ;
  assign n544 = n420 & n425 ;
  assign n545 = n419 | n544 ;
  assign n546 = n414 & n545 ;
  assign n547 = n413 | n546 ;
  assign n548 = n408 & n547 ;
  assign n549 = n407 | n548 ;
  assign n550 = n543 | n549 ;
  assign n551 = n469 | ~n472 ;
  assign n552 = G176 & ~G177 ;
  assign n553 = G60 & n552 ;
  assign n554 = ~G21 & n442 ;
  assign n555 = G21 & ~n442 ;
  assign n556 = n554 | n555 ;
  assign n557 = ~G176 & n556 ;
  assign n558 = G176 & ~n253 ;
  assign n559 = G177 & ~n558 ;
  assign n560 = ~n557 & n559 ;
  assign n561 = ~n553 & ~n560 ;
  assign n562 = G58 & n552 ;
  assign n563 = n439 & ~n443 ;
  assign n564 = n442 & ~n563 ;
  assign n565 = n445 | n564 ;
  assign n566 = G176 | n565 ;
  assign n567 = G176 & n243 ;
  assign n568 = G177 & ~n567 ;
  assign n569 = n566 & n568 ;
  assign n570 = ~n562 & ~n569 ;
  assign n571 = G48 & n552 ;
  assign n572 = G2 & n381 ;
  assign n573 = G2 | n381 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = G176 | n574 ;
  assign n576 = G176 & n318 ;
  assign n577 = G177 & ~n576 ;
  assign n578 = n575 & n577 ;
  assign n579 = ~n571 & ~n578 ;
  assign n580 = n469 & n472 ;
  assign n581 = n473 & ~n580 ;
  assign n582 = G173 | n579 ;
  assign n583 = G173 & ~n561 ;
  assign n584 = G172 & ~n583 ;
  assign n585 = n582 & n584 ;
  assign n586 = ~G172 & G173 ;
  assign n587 = G3 & n586 ;
  assign n588 = G172 | G173 ;
  assign n589 = G22 & ~n588 ;
  assign n590 = n587 | n589 ;
  assign n591 = n585 | n590 ;
  assign n592 = G19 & n552 ;
  assign n593 = n443 & n450 ;
  assign n594 = n449 | n593 ;
  assign n595 = n433 | n594 ;
  assign n596 = n434 & n595 ;
  assign n597 = n453 | n596 ;
  assign n598 = n479 | n597 ;
  assign n599 = n479 & n597 ;
  assign n600 = n598 & ~n599 ;
  assign n601 = ~G176 & n600 ;
  assign n602 = G176 & n268 ;
  assign n603 = G177 & ~n602 ;
  assign n604 = ~n601 & n603 ;
  assign n605 = ~n592 & ~n604 ;
  assign n606 = G59 & n552 ;
  assign n607 = n452 | n594 ;
  assign n608 = ~n435 & n607 ;
  assign n609 = n435 & ~n607 ;
  assign n610 = n608 | n609 ;
  assign n611 = ~G176 & n610 ;
  assign n612 = G176 & n256 ;
  assign n613 = G177 & ~n612 ;
  assign n614 = ~n611 & n613 ;
  assign n615 = ~n606 & ~n614 ;
  assign n616 = G50 & n552 ;
  assign n617 = n443 | n445 ;
  assign n618 = n451 | n617 ;
  assign n619 = n451 & n617 ;
  assign n620 = n618 & ~n619 ;
  assign n621 = ~G176 & n620 ;
  assign n622 = G176 & n277 ;
  assign n623 = G177 & ~n622 ;
  assign n624 = ~n621 & n623 ;
  assign n625 = ~n616 & ~n624 ;
  assign n626 = G174 | n579 ;
  assign n627 = G174 & ~n561 ;
  assign n628 = G175 & ~n627 ;
  assign n629 = n626 & n628 ;
  assign n630 = G174 & ~G175 ;
  assign n631 = G3 & n630 ;
  assign n632 = G174 | G175 ;
  assign n633 = G22 & ~n632 ;
  assign n634 = n631 | n633 ;
  assign n635 = n629 | n634 ;
  assign n636 = G53 & n552 ;
  assign n637 = G2 & n403 ;
  assign n638 = G2 & n402 ;
  assign n639 = n398 & n537 ;
  assign n640 = n399 | n639 ;
  assign n641 = ~n375 & n640 ;
  assign n642 = n375 & ~n640 ;
  assign n643 = n641 | n642 ;
  assign n644 = n638 | n643 ;
  assign n645 = ~n637 & n644 ;
  assign n646 = ~G176 & n645 ;
  assign n647 = G176 & n327 ;
  assign n648 = G177 & ~n647 ;
  assign n649 = ~n646 & n648 ;
  assign n650 = ~n636 & ~n649 ;
  assign n651 = G57 & n552 ;
  assign n652 = n388 & n394 ;
  assign n653 = n537 | n652 ;
  assign n654 = G2 | n537 ;
  assign n655 = n653 & n654 ;
  assign n656 = ~n400 & n655 ;
  assign n657 = n400 & ~n655 ;
  assign n658 = n656 | n657 ;
  assign n659 = ~G176 & n658 ;
  assign n660 = G176 & n356 ;
  assign n661 = G177 & ~n660 ;
  assign n662 = ~n659 & n661 ;
  assign n663 = ~n651 & ~n662 ;
  assign n664 = G56 & n552 ;
  assign n665 = n379 | n572 ;
  assign n666 = n387 & n665 ;
  assign n667 = n386 | n666 ;
  assign n668 = n394 | n667 ;
  assign n669 = n394 & n667 ;
  assign n670 = n668 & ~n669 ;
  assign n671 = ~G176 & n670 ;
  assign n672 = G176 & n365 ;
  assign n673 = G177 & ~n672 ;
  assign n674 = ~n671 & n673 ;
  assign n675 = ~n664 & ~n674 ;
  assign n676 = G55 & n552 ;
  assign n677 = n387 | n665 ;
  assign n678 = ~n666 & n677 ;
  assign n679 = ~G176 & n678 ;
  assign n680 = G176 & n337 ;
  assign n681 = G177 & ~n680 ;
  assign n682 = ~n679 & n681 ;
  assign n683 = ~n676 & ~n682 ;
  assign n684 = n456 & n469 ;
  assign n685 = n456 | n469 ;
  assign n686 = ~n684 & n685 ;
  assign n687 = n462 & n472 ;
  assign n688 = n462 | n472 ;
  assign n689 = ~n687 & n688 ;
  assign n690 = ~n686 & n689 ;
  assign n691 = n686 & ~n689 ;
  assign n692 = n690 | n691 ;
  assign n693 = G123 & G132 ;
  assign n694 = ~G123 & G133 ;
  assign n695 = n693 | n694 ;
  assign n696 = n438 | n448 ;
  assign n697 = n438 & n448 ;
  assign n698 = n696 & ~n697 ;
  assign n699 = n695 | n698 ;
  assign n700 = n695 & n698 ;
  assign n701 = n699 & ~n700 ;
  assign n702 = n432 & n476 ;
  assign n703 = G125 | n474 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = ~n442 & n704 ;
  assign n706 = n442 & ~n704 ;
  assign n707 = n705 | n706 ;
  assign n708 = n701 & ~n707 ;
  assign n709 = ~n701 & n707 ;
  assign n710 = n708 | n709 ;
  assign n711 = ~n692 & n710 ;
  assign n712 = n692 & ~n710 ;
  assign n713 = ~n711 & ~n712 ;
  assign n714 = n391 & n397 ;
  assign n715 = n391 | n397 ;
  assign n716 = ~n714 & n715 ;
  assign n717 = ~n378 & n384 ;
  assign n718 = n378 & ~n384 ;
  assign n719 = n717 | n718 ;
  assign n720 = n716 | n719 ;
  assign n721 = n716 & n719 ;
  assign n722 = n720 & ~n721 ;
  assign n723 = n412 & n418 ;
  assign n724 = n412 | n418 ;
  assign n725 = ~n723 & n724 ;
  assign n726 = G111 & G124 ;
  assign n727 = G112 & ~G124 ;
  assign n728 = n726 | n727 ;
  assign n729 = n424 & ~n728 ;
  assign n730 = ~n424 & n728 ;
  assign n731 = n729 | n730 ;
  assign n732 = ~n372 & n406 ;
  assign n733 = n372 & ~n406 ;
  assign n734 = n732 | n733 ;
  assign n735 = ~n731 & n734 ;
  assign n736 = n731 & ~n734 ;
  assign n737 = n735 | n736 ;
  assign n738 = ~n725 & n737 ;
  assign n739 = n725 & ~n737 ;
  assign n740 = n738 | n739 ;
  assign n741 = ~n722 & n740 ;
  assign n742 = n722 & ~n740 ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = n542 | n637 ;
  assign n745 = n429 & n744 ;
  assign n746 = n547 | n745 ;
  assign n747 = n409 | n746 ;
  assign n748 = n409 & n746 ;
  assign n749 = n747 & ~n748 ;
  assign n750 = n427 | n744 ;
  assign n751 = n427 & n744 ;
  assign n752 = n750 & ~n751 ;
  assign n753 = ~n574 & n678 ;
  assign n754 = n658 & n753 ;
  assign n755 = n670 & n754 ;
  assign n756 = n645 & n755 ;
  assign n757 = ~n752 & n756 ;
  assign n758 = n749 & n757 ;
  assign n759 = n428 & n744 ;
  assign n760 = n545 | n759 ;
  assign n761 = ~n415 & n760 ;
  assign n762 = n415 & ~n760 ;
  assign n763 = n761 | n762 ;
  assign n764 = n426 & n744 ;
  assign n765 = n425 | n744 ;
  assign n766 = ~n764 & n765 ;
  assign n767 = n421 | n766 ;
  assign n768 = n421 & n766 ;
  assign n769 = n767 & ~n768 ;
  assign n770 = n763 & ~n769 ;
  assign n771 = n758 & n770 ;
  assign n772 = n478 & n597 ;
  assign n773 = n477 | n772 ;
  assign n774 = n464 & n773 ;
  assign n775 = n463 | n773 ;
  assign n776 = ~n774 & n775 ;
  assign n777 = n459 & n776 ;
  assign n778 = n459 | n776 ;
  assign n779 = ~n777 & n778 ;
  assign n780 = n458 & n463 ;
  assign n781 = n457 | n780 ;
  assign n782 = n466 & n773 ;
  assign n783 = n781 | n782 ;
  assign n784 = n472 | n783 ;
  assign n785 = n472 & n783 ;
  assign n786 = n784 & ~n785 ;
  assign n787 = n465 & n773 ;
  assign n788 = n465 | n773 ;
  assign n789 = ~n787 & n788 ;
  assign n790 = n556 & n581 ;
  assign n791 = ~n565 & n790 ;
  assign n792 = n620 & n791 ;
  assign n793 = n610 & n792 ;
  assign n794 = n600 & n793 ;
  assign n795 = ~n789 & n794 ;
  assign n796 = ~n786 & n795 ;
  assign n797 = ~n779 & n796 ;
  assign n798 = G158 | n579 ;
  assign n799 = G158 & ~n561 ;
  assign n800 = G159 & ~n799 ;
  assign n801 = n798 & n800 ;
  assign n802 = G158 | G159 ;
  assign n803 = G81 & ~n802 ;
  assign n804 = G158 & ~G159 ;
  assign n805 = G80 & n804 ;
  assign n806 = n803 | n805 ;
  assign n807 = n801 | n806 ;
  assign n808 = G64 & n807 ;
  assign n809 = G160 | n579 ;
  assign n810 = G160 & ~n561 ;
  assign n811 = G161 & ~n810 ;
  assign n812 = n809 & n811 ;
  assign n813 = G160 | G161 ;
  assign n814 = G81 & ~n813 ;
  assign n815 = G160 & ~G161 ;
  assign n816 = G80 & n815 ;
  assign n817 = n814 | n816 ;
  assign n818 = n812 | n817 ;
  assign n819 = G64 & n818 ;
  assign n820 = G173 | n650 ;
  assign n821 = G173 & ~n605 ;
  assign n822 = G172 & ~n821 ;
  assign n823 = n820 & n822 ;
  assign n824 = G16 & n586 ;
  assign n825 = G14 & ~n588 ;
  assign n826 = n824 | n825 ;
  assign n827 = n823 | n826 ;
  assign n828 = G173 | n663 ;
  assign n829 = G173 & ~n615 ;
  assign n830 = G172 & ~n829 ;
  assign n831 = n828 & n830 ;
  assign n832 = G6 & ~n588 ;
  assign n833 = G27 & n586 ;
  assign n834 = n832 | n833 ;
  assign n835 = n831 | n834 ;
  assign n836 = G173 | n675 ;
  assign n837 = G173 & ~n625 ;
  assign n838 = G172 & ~n837 ;
  assign n839 = n836 & n838 ;
  assign n840 = G26 & n586 ;
  assign n841 = G5 & ~n588 ;
  assign n842 = n840 | n841 ;
  assign n843 = n839 | n842 ;
  assign n844 = G173 | n683 ;
  assign n845 = G173 & ~n570 ;
  assign n846 = G172 & ~n845 ;
  assign n847 = n844 & n846 ;
  assign n848 = G24 & n586 ;
  assign n849 = G25 & ~n588 ;
  assign n850 = n848 | n849 ;
  assign n851 = n847 | n850 ;
  assign n852 = G174 | n650 ;
  assign n853 = G174 & ~n605 ;
  assign n854 = G175 & ~n853 ;
  assign n855 = n852 & n854 ;
  assign n856 = G14 & ~n632 ;
  assign n857 = G16 & n630 ;
  assign n858 = n856 | n857 ;
  assign n859 = n855 | n858 ;
  assign n860 = G174 | n663 ;
  assign n861 = G174 & ~n615 ;
  assign n862 = G175 & ~n861 ;
  assign n863 = n860 & n862 ;
  assign n864 = G27 & n630 ;
  assign n865 = G6 & ~n632 ;
  assign n866 = n864 | n865 ;
  assign n867 = n863 | n866 ;
  assign n868 = G174 | n675 ;
  assign n869 = G174 & ~n625 ;
  assign n870 = G175 & ~n869 ;
  assign n871 = n868 & n870 ;
  assign n872 = G5 & ~n632 ;
  assign n873 = G26 & n630 ;
  assign n874 = n872 | n873 ;
  assign n875 = n871 | n874 ;
  assign n876 = G174 | n683 ;
  assign n877 = G174 & ~n570 ;
  assign n878 = G175 & ~n877 ;
  assign n879 = n876 & n878 ;
  assign n880 = G24 & n630 ;
  assign n881 = G25 & ~n632 ;
  assign n882 = n880 | n881 ;
  assign n883 = n879 | n882 ;
  assign n884 = G158 | n650 ;
  assign n885 = G158 & ~n605 ;
  assign n886 = G159 & ~n885 ;
  assign n887 = n884 & n886 ;
  assign n888 = G76 & ~n802 ;
  assign n889 = G86 & n804 ;
  assign n890 = n888 | n889 ;
  assign n891 = n887 | n890 ;
  assign n892 = G64 & n891 ;
  assign n893 = G158 | n683 ;
  assign n894 = G158 & ~n570 ;
  assign n895 = G159 & ~n894 ;
  assign n896 = n893 & n895 ;
  assign n897 = G72 & ~n802 ;
  assign n898 = G82 & n804 ;
  assign n899 = n897 | n898 ;
  assign n900 = n896 | n899 ;
  assign n901 = G64 & n900 ;
  assign n902 = G158 | n675 ;
  assign n903 = G158 & ~n625 ;
  assign n904 = G159 & ~n903 ;
  assign n905 = n902 & n904 ;
  assign n906 = G70 & ~n802 ;
  assign n907 = G71 & n804 ;
  assign n908 = n906 | n907 ;
  assign n909 = n905 | n908 ;
  assign n910 = G64 & n909 ;
  assign n911 = G158 | n663 ;
  assign n912 = G158 & ~n615 ;
  assign n913 = G159 & ~n912 ;
  assign n914 = n911 & n913 ;
  assign n915 = G68 & ~n802 ;
  assign n916 = G69 & n804 ;
  assign n917 = n915 | n916 ;
  assign n918 = n914 | n917 ;
  assign n919 = G64 & n918 ;
  assign n920 = G160 | n650 ;
  assign n921 = G160 & ~n605 ;
  assign n922 = G161 & ~n921 ;
  assign n923 = n920 & n922 ;
  assign n924 = G76 & ~n813 ;
  assign n925 = G86 & n815 ;
  assign n926 = n924 | n925 ;
  assign n927 = n923 | n926 ;
  assign n928 = G64 & n927 ;
  assign n929 = G160 | n683 ;
  assign n930 = G160 & ~n570 ;
  assign n931 = G161 & ~n930 ;
  assign n932 = n929 & n931 ;
  assign n933 = G72 & ~n813 ;
  assign n934 = G82 & n815 ;
  assign n935 = n933 | n934 ;
  assign n936 = n932 | n935 ;
  assign n937 = G64 & n936 ;
  assign n938 = G160 | n675 ;
  assign n939 = G160 & ~n625 ;
  assign n940 = G161 & ~n939 ;
  assign n941 = n938 & n940 ;
  assign n942 = G70 & ~n813 ;
  assign n943 = G71 & n815 ;
  assign n944 = n942 | n943 ;
  assign n945 = n941 | n944 ;
  assign n946 = G64 & n945 ;
  assign n947 = G160 | n663 ;
  assign n948 = G160 & ~n615 ;
  assign n949 = G161 & ~n948 ;
  assign n950 = n947 & n949 ;
  assign n951 = G68 & ~n813 ;
  assign n952 = G69 & n815 ;
  assign n953 = n951 | n952 ;
  assign n954 = n950 | n953 ;
  assign n955 = G64 & n954 ;
  assign n956 = G170 & n581 ;
  assign n957 = ~G61 & n469 ;
  assign n958 = G61 & ~n469 ;
  assign n959 = n957 | n958 ;
  assign n960 = G170 | n959 ;
  assign n961 = ~n956 & n960 ;
  assign n962 = G171 & ~n961 ;
  assign n963 = G178 & G62 ;
  assign n964 = G170 & ~G54 ;
  assign n965 = G170 | n246 ;
  assign n966 = ~n964 & n965 ;
  assign n967 = G171 | n966 ;
  assign n968 = ~n963 & n967 ;
  assign n969 = ~n962 & n968 ;
  assign n970 = n581 & n959 ;
  assign n971 = n581 | n959 ;
  assign n972 = n970 | ~n971 ;
  assign n973 = G54 & n552 ;
  assign n974 = ~G176 & n581 ;
  assign n975 = G176 & ~n246 ;
  assign n976 = G177 & ~n975 ;
  assign n977 = ~n974 & n976 ;
  assign n978 = ~n973 & ~n977 ;
  assign n979 = G52 & n552 ;
  assign n980 = G176 | n786 ;
  assign n981 = G176 & ~n249 ;
  assign n982 = G177 & ~n981 ;
  assign n983 = n980 & n982 ;
  assign n984 = ~n979 & ~n983 ;
  assign n985 = G47 & n552 ;
  assign n986 = G176 | n779 ;
  assign n987 = G176 & n224 ;
  assign n988 = G177 & ~n987 ;
  assign n989 = n986 & n988 ;
  assign n990 = ~n985 & ~n989 ;
  assign n991 = G43 & n552 ;
  assign n992 = G176 | n789 ;
  assign n993 = G176 & n233 ;
  assign n994 = G177 & ~n993 ;
  assign n995 = n992 & n994 ;
  assign n996 = ~n991 & ~n995 ;
  assign n997 = G155 & G99 ;
  assign n998 = n184 & n997 ;
  assign n999 = n179 & n998 ;
  assign n1000 = ~n506 & n999 ;
  assign n1001 = ~n533 & n1000 ;
  assign n1002 = ~n713 & n1001 ;
  assign n1003 = ~n743 & n1002 ;
  assign n1004 = G46 & n552 ;
  assign n1005 = ~G176 & n749 ;
  assign n1006 = G176 & n346 ;
  assign n1007 = G177 & ~n1006 ;
  assign n1008 = ~n1005 & n1007 ;
  assign n1009 = ~n1004 & ~n1008 ;
  assign n1010 = G45 & n552 ;
  assign n1011 = ~G176 & n763 ;
  assign n1012 = G176 & n298 ;
  assign n1013 = G177 & ~n1012 ;
  assign n1014 = ~n1011 & n1013 ;
  assign n1015 = ~n1010 & ~n1014 ;
  assign n1016 = G20 & n552 ;
  assign n1017 = G176 | n769 ;
  assign n1018 = G176 & n307 ;
  assign n1019 = G177 & ~n1018 ;
  assign n1020 = n1017 & n1019 ;
  assign n1021 = ~n1016 & ~n1020 ;
  assign n1022 = G44 & n552 ;
  assign n1023 = G176 | n752 ;
  assign n1024 = G176 & n289 ;
  assign n1025 = G177 & ~n1024 ;
  assign n1026 = n1023 & n1025 ;
  assign n1027 = ~n1022 & ~n1026 ;
  assign n1028 = G174 | n1009 ;
  assign n1029 = G174 & ~n978 ;
  assign n1030 = G175 & ~n1029 ;
  assign n1031 = n1028 & n1030 ;
  assign n1032 = G41 & ~n632 ;
  assign n1033 = G42 & n630 ;
  assign n1034 = n1032 | n1033 ;
  assign n1035 = n1031 | n1034 ;
  assign n1036 = G173 | n1009 ;
  assign n1037 = G173 & ~n978 ;
  assign n1038 = G172 & ~n1037 ;
  assign n1039 = n1036 & n1038 ;
  assign n1040 = G41 & ~n588 ;
  assign n1041 = G42 & n586 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = n1039 | n1042 ;
  assign n1044 = G173 & ~n984 ;
  assign n1045 = G173 | n1015 ;
  assign n1046 = G172 & n1045 ;
  assign n1047 = ~n1044 & n1046 ;
  assign n1048 = G17 & n586 ;
  assign n1049 = G18 & ~n588 ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = n1047 | n1050 ;
  assign n1052 = G173 & ~n990 ;
  assign n1053 = G173 | n1021 ;
  assign n1054 = G172 & n1053 ;
  assign n1055 = ~n1052 & n1054 ;
  assign n1056 = G39 & n586 ;
  assign n1057 = G40 & ~n588 ;
  assign n1058 = n1056 | n1057 ;
  assign n1059 = n1055 | n1058 ;
  assign n1060 = G173 & ~n996 ;
  assign n1061 = G173 | n1027 ;
  assign n1062 = G172 & n1061 ;
  assign n1063 = ~n1060 & n1062 ;
  assign n1064 = G36 & n586 ;
  assign n1065 = G15 & ~n588 ;
  assign n1066 = n1064 | n1065 ;
  assign n1067 = n1063 | n1066 ;
  assign n1068 = G174 | n1015 ;
  assign n1069 = G174 & ~n984 ;
  assign n1070 = G175 & ~n1069 ;
  assign n1071 = n1068 & n1070 ;
  assign n1072 = G17 & n630 ;
  assign n1073 = G18 & ~n632 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = n1071 | n1074 ;
  assign n1076 = G174 | n1021 ;
  assign n1077 = G174 & ~n990 ;
  assign n1078 = G175 & ~n1077 ;
  assign n1079 = n1076 & n1078 ;
  assign n1080 = G39 & n630 ;
  assign n1081 = G40 & ~n632 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = n1079 | n1082 ;
  assign n1084 = G174 | n1027 ;
  assign n1085 = G174 & ~n996 ;
  assign n1086 = G175 & ~n1085 ;
  assign n1087 = n1084 & n1086 ;
  assign n1088 = G36 & n630 ;
  assign n1089 = G15 & ~n632 ;
  assign n1090 = n1088 | n1089 ;
  assign n1091 = n1087 | n1090 ;
  assign n1092 = G158 & ~n996 ;
  assign n1093 = G158 | n1027 ;
  assign n1094 = G159 & n1093 ;
  assign n1095 = ~n1092 & n1094 ;
  assign n1096 = G77 & ~n802 ;
  assign n1097 = G87 & n804 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = n1095 | n1098 ;
  assign n1100 = G64 & n1099 ;
  assign n1101 = G158 & ~n990 ;
  assign n1102 = G158 | n1021 ;
  assign n1103 = G159 & n1102 ;
  assign n1104 = ~n1101 & n1103 ;
  assign n1105 = G75 & ~n802 ;
  assign n1106 = G85 & n804 ;
  assign n1107 = n1105 | n1106 ;
  assign n1108 = n1104 | n1107 ;
  assign n1109 = G64 & n1108 ;
  assign n1110 = G158 & ~n984 ;
  assign n1111 = G158 | n1015 ;
  assign n1112 = G159 & n1111 ;
  assign n1113 = ~n1110 & n1112 ;
  assign n1114 = G84 & n804 ;
  assign n1115 = G74 & ~n802 ;
  assign n1116 = n1114 | n1115 ;
  assign n1117 = n1113 | n1116 ;
  assign n1118 = G64 & n1117 ;
  assign n1119 = G158 | n1009 ;
  assign n1120 = G158 & ~n978 ;
  assign n1121 = G159 & ~n1120 ;
  assign n1122 = n1119 & n1121 ;
  assign n1123 = G73 & ~n802 ;
  assign n1124 = G83 & n804 ;
  assign n1125 = n1123 | n1124 ;
  assign n1126 = n1122 | n1125 ;
  assign n1127 = G64 & n1126 ;
  assign n1128 = G160 | n1027 ;
  assign n1129 = G160 & ~n996 ;
  assign n1130 = G161 & ~n1129 ;
  assign n1131 = n1128 & n1130 ;
  assign n1132 = G77 & ~n813 ;
  assign n1133 = G87 & n815 ;
  assign n1134 = n1132 | n1133 ;
  assign n1135 = n1131 | n1134 ;
  assign n1136 = G64 & n1135 ;
  assign n1137 = G160 | n1021 ;
  assign n1138 = G160 & ~n990 ;
  assign n1139 = G161 & ~n1138 ;
  assign n1140 = n1137 & n1139 ;
  assign n1141 = G85 & n815 ;
  assign n1142 = G75 & ~n813 ;
  assign n1143 = n1141 | n1142 ;
  assign n1144 = n1140 | n1143 ;
  assign n1145 = G64 & n1144 ;
  assign n1146 = G160 & ~n984 ;
  assign n1147 = G160 | n1015 ;
  assign n1148 = G161 & n1147 ;
  assign n1149 = ~n1146 & n1148 ;
  assign n1150 = G74 & ~n813 ;
  assign n1151 = G84 & n815 ;
  assign n1152 = n1150 | n1151 ;
  assign n1153 = n1149 | n1152 ;
  assign n1154 = G64 & n1153 ;
  assign n1155 = G160 | n1009 ;
  assign n1156 = G160 & ~n978 ;
  assign n1157 = G161 & ~n1156 ;
  assign n1158 = n1155 & n1157 ;
  assign n1159 = G73 & ~n813 ;
  assign n1160 = G83 & n815 ;
  assign n1161 = n1159 | n1160 ;
  assign n1162 = n1158 | n1161 ;
  assign n1163 = G64 & n1162 ;
  assign n1164 = ~G145 & n456 ;
  assign n1165 = n463 & ~n1164 ;
  assign n1166 = G145 & ~n464 ;
  assign n1167 = n1164 | n1166 ;
  assign n1168 = n456 & ~n465 ;
  assign n1169 = n1167 & ~n1168 ;
  assign n1170 = n1165 | n1169 ;
  assign n1171 = n686 & n1170 ;
  assign n1172 = n686 | n1170 ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1174 = n773 & ~n1173 ;
  assign n1175 = ~n457 & n463 ;
  assign n1176 = n458 & ~n1175 ;
  assign n1177 = ~n464 & n469 ;
  assign n1178 = n464 & ~n469 ;
  assign n1179 = n1177 | n1178 ;
  assign n1180 = n1176 & n1179 ;
  assign n1181 = n1176 | n1179 ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1183 = n773 | n1182 ;
  assign n1184 = ~n1174 & n1183 ;
  assign n1185 = n433 & ~n607 ;
  assign n1186 = ~n434 & n607 ;
  assign n1187 = n1185 | n1186 ;
  assign n1188 = G162 & n442 ;
  assign n1189 = n439 & n1188 ;
  assign n1190 = G162 | n439 ;
  assign n1191 = n444 & n1190 ;
  assign n1192 = ~n1189 & n1191 ;
  assign n1193 = ~n435 & n479 ;
  assign n1194 = n435 & ~n479 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = n1192 & n1195 ;
  assign n1197 = n1192 | n1195 ;
  assign n1198 = ~n1196 & n1197 ;
  assign n1199 = ~n451 & n1198 ;
  assign n1200 = n451 & ~n1198 ;
  assign n1201 = n1199 | n1200 ;
  assign n1202 = n1187 & ~n1201 ;
  assign n1203 = ~n1187 & n1201 ;
  assign n1204 = n1202 | n1203 ;
  assign n1205 = n1184 | n1204 ;
  assign n1206 = n1184 & n1204 ;
  assign n1207 = G176 | n1206 ;
  assign n1208 = n1205 & ~n1207 ;
  assign n1209 = ~G148 & G98 ;
  assign n1210 = ~G100 & G148 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = ~n253 & n1211 ;
  assign n1213 = n253 & ~n1211 ;
  assign n1214 = n1212 | n1213 ;
  assign n1215 = G100 | G121 ;
  assign n1216 = ~G101 & G121 ;
  assign n1217 = n1215 & ~n1216 ;
  assign n1218 = G147 & ~n1217 ;
  assign n1219 = G102 & G121 ;
  assign n1220 = ~G121 & G98 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = ~G147 & n1221 ;
  assign n1223 = n1218 | n1222 ;
  assign n1224 = n1214 | n1223 ;
  assign n1225 = n1214 & n1223 ;
  assign n1226 = n1224 & ~n1225 ;
  assign n1227 = G100 | G128 ;
  assign n1228 = ~G101 & G128 ;
  assign n1229 = n1227 & ~n1228 ;
  assign n1230 = G150 & ~n1229 ;
  assign n1231 = G102 & G128 ;
  assign n1232 = ~G128 & G98 ;
  assign n1233 = n1231 | n1232 ;
  assign n1234 = ~G150 & n1233 ;
  assign n1235 = n1230 | n1234 ;
  assign n1236 = G100 | G126 ;
  assign n1237 = ~G101 & G126 ;
  assign n1238 = n1236 & ~n1237 ;
  assign n1239 = G149 & ~n1238 ;
  assign n1240 = G102 & G126 ;
  assign n1241 = ~G126 & G98 ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = ~G149 & n1242 ;
  assign n1244 = n1239 | n1243 ;
  assign n1245 = n1235 | n1244 ;
  assign n1246 = n1235 & n1244 ;
  assign n1247 = n1245 & ~n1246 ;
  assign n1248 = n1226 | n1247 ;
  assign n1249 = n1226 & n1247 ;
  assign n1250 = n1248 & ~n1249 ;
  assign n1251 = n224 | n233 ;
  assign n1252 = ~n234 & n1251 ;
  assign n1253 = ~n246 & n249 ;
  assign n1254 = n250 | n1253 ;
  assign n1255 = n1252 | n1254 ;
  assign n1256 = n1252 & n1254 ;
  assign n1257 = n1255 & ~n1256 ;
  assign n1258 = n1250 | n1257 ;
  assign n1259 = n1250 & n1257 ;
  assign n1260 = G176 & ~n1259 ;
  assign n1261 = n1258 & n1260 ;
  assign n1262 = G177 & ~n1261 ;
  assign n1263 = ~n1208 & n1262 ;
  assign n1264 = ~G51 & n552 ;
  assign n1265 = ~n1263 & ~n1264 ;
  assign n1266 = n381 & n386 ;
  assign n1267 = n381 | n387 ;
  assign n1268 = ~n388 & n1267 ;
  assign n1269 = n379 | n386 ;
  assign n1270 = ~n534 & n1269 ;
  assign n1271 = n1268 | n1270 ;
  assign n1272 = ~n1266 & n1271 ;
  assign n1273 = n537 & ~n1272 ;
  assign n1274 = ~n537 & n1272 ;
  assign n1275 = n1273 | n1274 ;
  assign n1276 = n643 | n1275 ;
  assign n1277 = n643 & n1275 ;
  assign n1278 = G157 | n1277 ;
  assign n1279 = n1276 & ~n1278 ;
  assign n1280 = n380 & n385 ;
  assign n1281 = n380 | n386 ;
  assign n1282 = ~n1280 & n1281 ;
  assign n1283 = n653 & ~n1282 ;
  assign n1284 = ~n653 & n1282 ;
  assign n1285 = n1283 | n1284 ;
  assign n1286 = n375 | n1268 ;
  assign n1287 = n375 & n1268 ;
  assign n1288 = n1286 & ~n1287 ;
  assign n1289 = n402 | n640 ;
  assign n1290 = n1288 & ~n1289 ;
  assign n1291 = ~n1288 & n1289 ;
  assign n1292 = n1290 | n1291 ;
  assign n1293 = n1285 & n1292 ;
  assign n1294 = n1285 | n1292 ;
  assign n1295 = G157 & n1294 ;
  assign n1296 = ~n1293 & n1295 ;
  assign n1297 = n1279 | n1296 ;
  assign n1298 = n428 | n545 ;
  assign n1299 = ~n413 & n1298 ;
  assign n1300 = n414 & ~n1299 ;
  assign n1301 = n409 | n421 ;
  assign n1302 = n409 & n421 ;
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = n425 | n1298 ;
  assign n1305 = ~n544 & n1304 ;
  assign n1306 = n1303 & n1305 ;
  assign n1307 = n1303 | n1305 ;
  assign n1308 = ~n1306 & n1307 ;
  assign n1309 = n1300 & n1308 ;
  assign n1310 = n1300 | n1308 ;
  assign n1311 = ~n1309 & n1310 ;
  assign n1312 = n542 & n1311 ;
  assign n1313 = n413 | n545 ;
  assign n1314 = ~n546 & n1313 ;
  assign n1315 = ~n415 & n426 ;
  assign n1316 = n415 & ~n426 ;
  assign n1317 = n1315 | n1316 ;
  assign n1318 = n1303 & ~n1317 ;
  assign n1319 = ~n1303 & n1317 ;
  assign n1320 = n1318 | n1319 ;
  assign n1321 = n1314 | n1320 ;
  assign n1322 = n1314 & n1320 ;
  assign n1323 = n542 | n1322 ;
  assign n1324 = n1321 & ~n1323 ;
  assign n1325 = G157 | n1324 ;
  assign n1326 = n1312 | n1325 ;
  assign n1327 = n403 | n542 ;
  assign n1328 = n1311 & n1327 ;
  assign n1329 = ~n403 & n1324 ;
  assign n1330 = G157 & ~n1329 ;
  assign n1331 = ~n1328 & n1330 ;
  assign n1332 = n1326 & ~n1331 ;
  assign n1333 = n394 | n400 ;
  assign n1334 = ~n401 & n1333 ;
  assign n1335 = n1332 & ~n1334 ;
  assign n1336 = ~n1332 & n1334 ;
  assign n1337 = n1335 | n1336 ;
  assign n1338 = ~n1297 & n1337 ;
  assign n1339 = n1297 & ~n1337 ;
  assign n1340 = G176 | n1339 ;
  assign n1341 = n1338 | n1340 ;
  assign n1342 = G100 | G90 ;
  assign n1343 = ~G101 & G90 ;
  assign n1344 = n1342 & ~n1343 ;
  assign n1345 = G143 & ~n1344 ;
  assign n1346 = G102 & G90 ;
  assign n1347 = ~G90 & G98 ;
  assign n1348 = n1346 | n1347 ;
  assign n1349 = ~G143 & n1348 ;
  assign n1350 = n1345 | n1349 ;
  assign n1351 = G100 | G92 ;
  assign n1352 = ~G101 & G92 ;
  assign n1353 = n1351 & ~n1352 ;
  assign n1354 = G144 & ~n1353 ;
  assign n1355 = G102 & G92 ;
  assign n1356 = ~G92 & G98 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = ~G144 & n1357 ;
  assign n1359 = n1354 | n1358 ;
  assign n1360 = n1350 & ~n1359 ;
  assign n1361 = ~n1350 & n1359 ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = G100 | G94 ;
  assign n1364 = ~G101 & G94 ;
  assign n1365 = n1363 & ~n1364 ;
  assign n1366 = G140 & ~n1365 ;
  assign n1367 = G102 & G94 ;
  assign n1368 = ~G94 & G98 ;
  assign n1369 = n1367 | n1368 ;
  assign n1370 = ~G140 & n1369 ;
  assign n1371 = n1366 | n1370 ;
  assign n1372 = n346 & n1371 ;
  assign n1373 = n346 | n1371 ;
  assign n1374 = ~n1372 & n1373 ;
  assign n1375 = ~n1362 & n1374 ;
  assign n1376 = n1362 & ~n1374 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = G100 | G107 ;
  assign n1379 = ~G101 & G107 ;
  assign n1380 = n1378 & ~n1379 ;
  assign n1381 = G139 & ~n1380 ;
  assign n1382 = G102 & G107 ;
  assign n1383 = ~G107 & G98 ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = ~G139 & n1384 ;
  assign n1386 = n1381 | n1385 ;
  assign n1387 = G100 | G105 ;
  assign n1388 = ~G101 & G105 ;
  assign n1389 = n1387 & ~n1388 ;
  assign n1390 = G138 & ~n1389 ;
  assign n1391 = G102 & G105 ;
  assign n1392 = ~G105 & G98 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = ~G138 & n1393 ;
  assign n1395 = n1390 | n1394 ;
  assign n1396 = n1386 & n1395 ;
  assign n1397 = n1386 | n1395 ;
  assign n1398 = ~n1396 & n1397 ;
  assign n1399 = G100 | G96 ;
  assign n1400 = ~G101 & G96 ;
  assign n1401 = n1399 & ~n1400 ;
  assign n1402 = G141 & ~n1401 ;
  assign n1403 = G102 & G96 ;
  assign n1404 = ~G96 & G98 ;
  assign n1405 = n1403 | n1404 ;
  assign n1406 = ~G141 & n1405 ;
  assign n1407 = n1402 | n1406 ;
  assign n1408 = G100 | G109 ;
  assign n1409 = ~G101 & G109 ;
  assign n1410 = n1408 & ~n1409 ;
  assign n1411 = G135 & ~n1410 ;
  assign n1412 = G102 & G109 ;
  assign n1413 = ~G109 & G98 ;
  assign n1414 = n1412 | n1413 ;
  assign n1415 = ~G135 & n1414 ;
  assign n1416 = n1411 | n1415 ;
  assign n1417 = G100 | G103 ;
  assign n1418 = ~G101 & G103 ;
  assign n1419 = n1417 & ~n1418 ;
  assign n1420 = G137 & ~n1419 ;
  assign n1421 = G102 & G103 ;
  assign n1422 = ~G103 & G98 ;
  assign n1423 = n1421 | n1422 ;
  assign n1424 = ~G137 & n1423 ;
  assign n1425 = n1420 | n1424 ;
  assign n1426 = n1416 & n1425 ;
  assign n1427 = n1416 | n1425 ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = n1407 & ~n1428 ;
  assign n1430 = ~n1407 & n1428 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = ~n1398 & n1431 ;
  assign n1433 = n1398 & ~n1431 ;
  assign n1434 = n1432 | n1433 ;
  assign n1435 = ~n1377 & n1434 ;
  assign n1436 = n1377 & ~n1434 ;
  assign n1437 = G176 & ~n1436 ;
  assign n1438 = ~n1435 & n1437 ;
  assign n1439 = G177 & ~n1438 ;
  assign n1440 = n1341 & n1439 ;
  assign n1441 = ~G49 & n552 ;
  assign n1442 = ~n1440 & ~n1441 ;
  assign n1443 = ~G177 & G38 ;
  assign n1444 = n1440 | n1443 ;
  assign n1445 = G173 | n1444 ;
  assign n1446 = ~G177 & G37 ;
  assign n1447 = n1263 | n1446 ;
  assign n1448 = G173 & ~n1447 ;
  assign n1449 = G172 & ~n1448 ;
  assign n1450 = n1445 & n1449 ;
  assign n1451 = G23 & ~n588 ;
  assign n1452 = G4 & n586 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = n1450 | n1453 ;
  assign n1455 = G174 | n1444 ;
  assign n1456 = G174 & ~n1447 ;
  assign n1457 = G175 & ~n1456 ;
  assign n1458 = n1455 & n1457 ;
  assign n1459 = G23 & ~n632 ;
  assign n1460 = G4 & n630 ;
  assign n1461 = n1459 | n1460 ;
  assign n1462 = n1458 | n1461 ;
  assign n1463 = G158 | n1444 ;
  assign n1464 = G158 & ~n1447 ;
  assign n1465 = G159 & ~n1464 ;
  assign n1466 = n1463 & n1465 ;
  assign n1467 = G79 & ~n802 ;
  assign n1468 = G78 & n804 ;
  assign n1469 = n1467 | n1468 ;
  assign n1470 = n1466 | n1469 ;
  assign n1471 = ~G64 | ~n1470 ;
  assign n1472 = G160 | n1444 ;
  assign n1473 = G160 & ~n1447 ;
  assign n1474 = G161 & ~n1473 ;
  assign n1475 = n1472 & n1474 ;
  assign n1476 = G79 & ~n813 ;
  assign n1477 = G78 & n815 ;
  assign n1478 = n1476 | n1477 ;
  assign n1479 = n1475 | n1478 ;
  assign n1480 = ~G64 | ~n1479 ;
  assign G5193 = ~G66 ;
  assign G5194 = ~G113 ;
  assign G5195 = ~G165 ;
  assign G5196 = ~G151 ;
  assign G5197 = ~G127 ;
  assign G5198 = ~G131 ;
  assign G5199 = n179 ;
  assign G5200 = ~G152 ;
  assign G5201 = ~G151 ;
  assign G5202 = ~G151 ;
  assign G5203 = ~G125 ;
  assign G5204 = ~G129 ;
  assign G5205 = n180 ;
  assign G5206 = ~G99 ;
  assign G5207 = ~G153 ;
  assign G5208 = ~G156 ;
  assign G5209 = ~G155 ;
  assign G5210 = n181 ;
  assign G5211 = n182 ;
  assign G5212 = n183 ;
  assign G5213 = n184 ;
  assign G5214 = G64 ;
  assign G5215 = G66 ;
  assign G5216 = G1 ;
  assign G5217 = G152 ;
  assign G5218 = G114 ;
  assign G5219 = G152 ;
  assign G5220 = n186 ;
  assign G5221 = n185 ;
  assign G5222 = ~G1 ;
  assign G5223 = ~G1 ;
  assign G5224 = ~G1 ;
  assign G5225 = ~G1 ;
  assign G5226 = ~G114 ;
  assign G5227 = ~G114 ;
  assign G5228 = n190 ;
  assign G5229 = n194 ;
  assign G5230 = n194 ;
  assign G5231 = n195 ;
  assign G5232 = n200 ;
  assign G5233 = n205 ;
  assign G5234 = n210 ;
  assign G5235 = n215 ;
  assign G5236 = n280 ;
  assign G5237 = n369 ;
  assign G5238 = n431 ;
  assign G5239 = n482 ;
  assign G5240 = n482 ;
  assign G5241 = n431 ;
  assign G5242 = n506 ;
  assign G5243 = n533 ;
  assign G5244 = n550 ;
  assign G5245 = n551 ;
  assign G5246 = n550 ;
  assign G5247 = n551 ;
  assign G5248 = n561 ;
  assign G5249 = n570 ;
  assign G5250 = n579 ;
  assign G5251 = n581 ;
  assign G5252 = n591 ;
  assign G5253 = n605 ;
  assign G5254 = n615 ;
  assign G5255 = n625 ;
  assign G5256 = n635 ;
  assign G5257 = n650 ;
  assign G5258 = n663 ;
  assign G5259 = n675 ;
  assign G5260 = n683 ;
  assign G5261 = n713 ;
  assign G5262 = n743 ;
  assign G5263 = n771 ;
  assign G5264 = n797 ;
  assign G5265 = n808 ;
  assign G5266 = n819 ;
  assign G5267 = n827 ;
  assign G5268 = n835 ;
  assign G5269 = n843 ;
  assign G5270 = n851 ;
  assign G5271 = n859 ;
  assign G5272 = n867 ;
  assign G5273 = n875 ;
  assign G5274 = n883 ;
  assign G5275 = n892 ;
  assign G5276 = n901 ;
  assign G5277 = n910 ;
  assign G5278 = n919 ;
  assign G5279 = n928 ;
  assign G5280 = n937 ;
  assign G5281 = n946 ;
  assign G5282 = n955 ;
  assign G5283 = n969 ;
  assign G5284 = n972 ;
  assign G5285 = n978 ;
  assign G5286 = n984 ;
  assign G5287 = n990 ;
  assign G5288 = n996 ;
  assign G5289 = n1003 ;
  assign G5290 = n1009 ;
  assign G5291 = n1015 ;
  assign G5292 = n1021 ;
  assign G5293 = n1027 ;
  assign G5294 = n1035 ;
  assign G5295 = n1043 ;
  assign G5296 = n1051 ;
  assign G5297 = n1059 ;
  assign G5298 = n1067 ;
  assign G5299 = n1075 ;
  assign G5300 = n1083 ;
  assign G5301 = n1091 ;
  assign G5302 = n1100 ;
  assign G5303 = n1109 ;
  assign G5304 = n1118 ;
  assign G5305 = n1127 ;
  assign G5306 = n1136 ;
  assign G5307 = n1145 ;
  assign G5308 = n1154 ;
  assign G5309 = n1163 ;
  assign G5310 = n1265 ;
  assign G5311 = n1442 ;
  assign G5312 = n1454 ;
  assign G5313 = n1462 ;
  assign G5314 = n1471 ;
  assign G5315 = n1480 ;
endmodule