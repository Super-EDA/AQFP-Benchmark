module multiplier_8 (b_4_,a_1_,a_2_,b_1_,b_7_,a_6_,a_4_,b_2_,a_7_,a_5_,b_5_,b_3_,b_6_,b_0_,a_3_,a_0_,s_1_,s_8_,s_3_,s_5_,s_9_,s_2_,s_11_,s_15_,s_4_,s_10_,s_14_,s_7_,s_13_,s_12_,s_6_,s_0_);
  input b_4_,a_1_,a_2_,b_1_,b_7_,a_6_,a_4_,b_2_,a_7_,a_5_,b_5_,b_3_,b_6_,b_0_,a_3_,a_0_;
  output s_1_,s_8_,s_3_,s_5_,s_9_,s_2_,s_11_,s_15_,s_4_,s_10_,s_14_,s_7_,s_13_,s_12_,s_6_,s_0_;
  wire _w_2573,_w_2571,_w_2569,_w_2568,_w_2567,_w_2566,_w_2564,_w_2563,_w_2561,_w_2565,_w_2559,_w_2558,_w_2555,_w_2554,_w_2553,_w_2551,_w_2550,_w_2549,_w_2546,_w_2541,_w_2538,_w_2536,_w_2535,_w_2534,_w_2532,_w_2531,_w_2529,_w_2527,_w_2524,_w_2523,_w_2522,_w_2520,_w_2518,_w_2517,_w_2515,_w_2514,_w_2513,_w_2512,_w_2505,_w_2504,_w_2503,_w_2501,_w_2499,_w_2497,_w_2496,_w_2492,_w_2491,_w_2490,_w_2486,_w_2485,_w_2483,_w_2482,_w_2481,_w_2478,_w_2572,_w_2477,_w_2474,_w_2472,_w_2471,_w_2470,_w_2469,_w_2468,_w_2467,_w_2465,_w_2464,_w_2463,_w_2507,_w_2462,_w_2461,_w_2459,_w_2458,_w_2455,_w_2454,_w_2453,_w_2452,_w_2451,_w_2450,_w_2449,_w_2446,_w_2445,_w_2443,_w_2442,_w_2440,_w_2439,_w_2438,_w_2437,_w_2436,_w_2435,_w_2434,_w_2433,_w_2432,_w_2431,_w_2428,_w_2425,_w_2424,_w_2423,_w_2422,_w_2419,_w_2418,_w_2417,_w_2416,_w_2414,_w_2412,_w_2409,_w_2407,_w_2406,_w_2405,_w_2404,_w_2403,_w_2402,_w_2401,_w_2400,_w_2398,_w_2397,_w_2395,_w_2394,_w_2390,_w_2389,_w_2388,_w_2387,_w_2391,_w_2386,_w_2385,_w_2384,_w_2383,_w_2382,_w_2381,_w_2380,_w_2379,_w_2375,_w_2374,_w_2373,_w_2488,_w_2372,_w_2368,_w_2367,_w_2366,_w_2365,_w_2364,_w_2363,_w_2362,_w_2361,_w_2358,_w_2357,n326_1,n367_0,n168_0,n126_1,n126_0,_w_1970,n100_1,_w_1675,n122_0,n121_1,n218_0,_w_1623,_w_1385,n154_1,n175_0,n154_0,n122_1,n401_1,n115_0,_w_1744,_w_2326,n35_0,n295_0,a_7__11,_w_1694,a_7__5,a_7__3,_w_1632,b_0__9,b_0__8,n137,_w_1728,b_0__7,n225_1,_w_1937,n130_0,n310_1,n41_0,n390_1,n390_0,n305,n153_3,a_7__1,_w_2078,n153_0,n28_0,n25_1,_w_1468,b_3__3,n438,_w_1670,n164_0,n418_0,_w_1624,n109_0,_w_2539,n268_1,_w_2480,_w_1729,_w_1773,_w_2290,n24_0,n186_1,_w_2498,n186_0,n184_0,n255_1,n260_1,n255_0,_w_1659,_w_2530,n205_1,n375_1,n32_0,n197_1,_w_1940,n435,n284_3,n131_1,n284_0,b_1__8,n99_0,b_1__7,_w_1565,b_3__10,n253_1,b_1__6,b_0__3,b_1__4,_w_1414,n36_0,n350,n19_2,n56_1,n289_0,_w_1607,a_3__10,_w_2322,_w_1870,_w_2371,_w_1920,a_3__1,_w_1858,b_5__11,b_5__6,_w_1967,b_5__5,_w_1861,b_5__0,n214_0,_w_1780,_w_2218,a_5__10,a_5__7,_w_2248,a_5__2,_w_2429,_w_1484,_w_2203,a_6__9,n363_1,n378,a_6__8,n78_0,n211,a_6__7,_w_2202,a_6__6,n419,_w_1403,_w_1815,n62_2,_w_1994,n157_1,n242_0,_w_1849,n404_1,n404_0,_w_1821,b_7__11,_w_2159,n405_0,b_7__10,b_7__7,n394,a_3__4,_w_2162,_w_2548,n175_1,b_7__5,_w_1647,b_7__4,_w_2064,b_7__2,_w_1709,a_1__1,_w_2148,n43,n408_0,n54,_w_1382,b_4__11,_w_2151,b_4__10,n385,n321_1,b_4__7,b_4__4,b_4__3,_w_2344,n391_1,n261_1,a_5__5,n437_0,n287,_w_1449,n76_1,n139,n76_0,_w_1749,b_6__6,_w_1775,b_6__0,_w_2275,n133_1,n424_1,a_4__10,a_4__8,n178_1,n174_1,b_2__9,n385_1,n291,b_2__1,_w_2067,b_2__0,_w_2024,n73_0,a_5__8,n23,n142_0,a_2__10,_w_1518,a_2__8,a_2__7,n258_1,n367,a_2__6,a_2__3,n74,a_2__2,_w_1786,_w_1911,n214_1,_w_2164,n63_0,_w_1877,_w_1953,a_0__7,a_0__6,_w_2489,_w_1660,n74_0,_w_1996,a_0__2,n71,_w_2360,n45_0,n418_1,n95_0,n46_1,_w_2135,n69_1,n69_0,n168_1,_w_2276,n391_0,b_1__9,n55_2,n182_0,n416_1,a_4__1,a_7__9,n89,n190,n19_0,n40_0,n50_1,n103,n331_1,n331_0,_w_1363,n227_0,n242_1,_w_1717,_w_1929,n173_0,b_6__7,n285_0,b_6__3,_w_1730,_w_1928,n61_1,_w_1519,_w_1453,a_6__13,_w_1777,n61_0,_w_2460,_w_2298,n145_0,_w_1464,b_1__0,n230,_w_1523,n64_0,n172_1,n384_1,n85_0,n172_0,n26_0,n79_0,n205,n156_0,_w_1595,n227_1,n293_0,n130_1,_w_1381,_w_1547,n111_1,_w_1290,n92_1,n157,n62_6,n309_1,n92_0,n167_0,n188_1,n23_1,b_1__2,n411_0,n23_0,n44_1,_w_2188,b_1__3,a_4__7,n286_1,n190_0,_w_1423,n436_1,n410_1,_w_2004,_w_1763,_w_1433,n90_1,n44,_w_2071,n198_1,n93_1,n150_0,n156_1,b_0__4,n93_0,n364_1,b_0__6,n18_0,n56,_w_2201,n119_0,_w_1842,_w_2149,n305_1,_w_1956,n95_1,n208_0,_w_1452,n400_0,n200,_w_2186,n103_1,_w_1631,n398_1,n398_0,n65_1,n65,_w_1907,n199_1,_w_1604,n105_1,n123,n55_0,n105_0,n39_0,n134,n165_1,n110_1,n411,n197_0,_w_1418,n244_0,_w_1356,n133_0,n203_1,_w_1394,n378_0,n246_1,n332_1,_w_1446,_w_2312,_w_1748,n246_0,n248_0,n251_2,_w_1865,n403_1,_w_2495,n182_1,n403_0,n254_2,n433_0,b_5__8,n215_3,_w_2359,n254_1,_w_2519,_w_2070,n63_1,_w_1878,n254_0,_w_1401,n251_0,n259_1,n140_1,_w_1625,n259_0,_w_2457,a_0__5,_w_1746,_w_1978,n268_0,a_3__9,n272_1,b_7__6,n332,n272_0,_w_1320,n383_0,n274_0,b_6__1,_w_2020,n344_1,_w_2212,n79_1,_w_1493,n370_0,_w_1761,n344_0,n276_0,n436_0,n279_1,n209_0,n136_0,n279_0,b_4__6,n83_0,_w_2244,n324_3,_w_2557,n213_1,n324_2,n324_0,n77,n57,n287_0,n201,_w_2370,n294_0,_w_1573,n371_0,n372_1,n34_1,n307_1,_w_1795,n372_0,n408_1,n117,n298_1,n298_0,a_7__13,n300_1,n290_0,n34_0,n341_0,n269_0,n304_0,n422_0,b_3__11,n45,n260_0,n316_1,n401,n358_1,n423_0,n358_0,_w_2281,n39_1,n274,_w_1549,n317_1,_w_2346,n102_1,_w_2157,n319_1,n301_0,n416_0,_w_2421,n322_1,_w_1375,_w_1808,n322_0,_w_2376,b_4__5,n228,_w_2487,_w_1577,a_3__7,n342,a_6__10,n235,_w_1822,n347_1,_w_1361,_w_2181,_w_2313,n58_1,n219,n204_0,n174,n55_1,n213,a_7__4,_w_2196,n88,_w_2194,n353,n67_0,n209,_w_2117,n203,n432,_w_1725,n236,n364_0,n373,a_5__12,_w_1704,_w_2107,_w_2198,n229,a_6__2,n189,n64_1,_w_1944,_w_2065,_w_1892,n307,_w_1461,n180,n155,n179,n368,_w_1457,_w_2494,n171,_w_1983,n354,_w_1313,n166,n67_1,n289_1,n62,n25_0,n336_0,n396,n184,_w_1741,n429_0,n38_0,_w_1917,n257_0,n136_1,n280_0,n384,n202,_w_1508,n148,_w_2332,b_6__4,n49_0,n168_3,n53_1,n134_0,n159,n75_1,b_0__0,n300_0,_w_1671,n415,_w_1553,_w_2091,n141,n104,n142,n140,b_7__9,n52_0,n273_1,_w_1788,n142_1,_w_2289,n240,_w_2560,_w_1328,_w_2430,n84,n144_0,_w_2229,n288,n291_0,_w_2101,a_6__12,n430,_w_1790,n168,n216,n118,n135,n168_2,n175,n431,n37_1,n209_1,_w_1830,n130,_w_2042,n256,n127,_w_2441,n451,n17,_w_1654,_w_2134,_w_2350,n352,_w_1962,n149,_w_1359,n381_0,n70,_w_2230,b_3__0,_w_2223,a_3__2,n375_0,n121,n170,n261_0,n178,n154,n32_1,b_0__5,n360_0,a_3__8,_w_1578,n115,n78_1,n66,n314,_w_1421,_w_2204,n348_0,n138_0,_w_2476,_w_1350,a_4__2,n167_1,n119_1,n360_1,_w_2106,n82,_w_2155,n173,n59,n38,n68,_w_2377,a_7__12,n302_0,n404_2,_w_2183,n433_1,n363,_w_2178,n42,n436,n366,_w_1527,_w_1560,_w_2021,n390,n65_0,n170_1,n152,n317_0,n333,n212_1,n28,n24,n345,n392,a_5__11,n19,n392_0,n153_1,_w_1349,_w_2163,n225_0,n164_1,_w_1836,_w_1417,_w_1475,_w_2139,_w_1894,n214,n185,n443,_w_1326,b_1__5,n416,_w_1323,a_0__8,n138,n165_0,n286_0,n102,n376_1,n110_0,_w_2271,_w_2411,n150,n124,n197,b_5__2,n119,_w_2264,_w_1845,n422_1,a_5__6,n389_1,_w_1934,n223,n234_1,_w_2079,_w_2574,n284,n295,n217,n198,n439_1,n86_0,_w_1551,n60,n125,b_1__11,_w_1955,b_5__4,_w_1476,n337,n318_1,n324,n362,_w_2174,n386,n128_0,n35_1,_w_2392,_w_1927,_w_2552,_w_1693,n91,_w_2511,_w_1932,n143,_w_2351,n346,n369,_w_1481,n404,b_4__8,n40_1,_w_2274,n335_0,n294_1,n424_0,_w_1843,n280_1,n22_1,n405,n270_1,n397_1,_w_1465,_w_1628,b_2__2,_w_1335,_w_1314,n277,n438_0,_w_1422,_w_1667,n247,n252,a_5__9,n29_0,n22_0,_w_2168,n221,n206,n321_0,n348_1,n425,n167,b_3__7,n83,n52,_w_1436,n18,a_2__5,_w_1677,n237_1,_w_2034,n282_1,n308_0,a_5__3,_w_2547,_w_2369,n308,n69,n447,a_1__4,n367_1,_w_1517,_w_1764,_w_1991,n312,_w_1703,n40,_w_1691,_w_2023,n222,n68_0,_w_2190,n110,n50,n53,n227,n114_0,b_0__11,n375,n218_1,n290,_w_1918,_w_2228,n37,n44_0,_w_1972,_w_1666,n153_2,a_2__4,n27,n297_0,n132,_w_2126,n210,_w_1525,_w_2325,n102_0,n434_0,b_6__12,n176,a_3__3,n430_0,n50_0,n259,n144,_w_1834,n271,n218,_w_1747,n294,n331,b_6__5,_w_1367,n356_1,_w_2537,_w_1360,n304_1,n74_1,_w_2525,_w_1473,n46,n61,n449,n193,n435_1,n99_1,n147,n361,n64,_w_2266,n275,n425_0,n91_1,n357,n338_1,n305_0,n213_0,_w_1524,n41,_w_1448,_w_1301,n270,n273_0,_w_1672,_w_2160,n75,n58,n84_1,a_6__11,_w_1512,n111,n52_1,a_2__9,_w_2288,n172,a_0__11,n131,_w_1566,n59_0,n26,n103_0,b_2__5,n224_1,n173_1,_w_1824,n195,n297_1,_w_2249,n341_1,_w_2221,n269_1,_w_1743,n96,n414_1,_w_2039,n22,n79,n323_1,_w_2396,_w_1724,n156,n293,n309,n29,_w_1420,_w_1496,n161,n90_0,n391,n351_1,n445,n87,b_5__9,n240_0,a_0__1,a_6__5,n144_1,n106,n113,_w_1896,n31_1,n286,n285_1,n93,_w_2150,n95,n398,n301_1,b_3__4,a_4__6,n34,n400,n208_1,n97,_w_1306,n254,_w_2169,n345_0,_w_2543,_w_1793,n38_1,n284_1,_w_2540,n210_1,n250_0,_w_1636,n324_1,n101,n62_5,_w_1998,b_7__0,n192,n378_1,b_3__9,b_5__3,n376_0,n152_1,n163,n47_1,n122,n131_0,_w_2209,n68_1,n187,n377,n257_1,_w_1658,_w_1814,n347,n427,_w_1805,n243,_w_2123,n245,a_6__4,n370,_w_1462,n246,a_0__0,_w_2570,n300,n73_1,a_4__3,n287_1,n409_1,n224_0,b_1__1,n145_1,_w_1891,_w_1315,_w_2122,n249,n128,n321,n250,_w_1905,a_5__1,_w_1982,_w_1329,_w_1699,b_2__3,n403,_w_1586,_w_2211,_w_1450,n405_1,_w_1988,n257,n258,a_3__6,n420_0,_w_1856,n266,_w_1714,n420_1,n269,n397_0,n55,n273,_w_1341,_w_1325,n418,n407,_w_1477,n282,n182,n279,n129_0,n389_2,n280,n392_1,_w_2475,n281,n268,n283,n128_1,n309_0,n244,n285,n292,_w_2057,n255_2,_w_1366,_w_1947,n296,_w_1635,_w_1922,a_4__5,n372,a_2__0,n177_0,_w_1309,_w_1540,n278,_w_2329,n408,_w_2262,n389_3,n382,_w_2257,n297,_w_1487,_w_2047,a_4__9,_w_1721,n371,n109,n414,n298,n31,n240_2,_w_1357,b_6__8,n410,_w_1738,n303,_w_1888,n270_0,_w_1984,n423,n301,n117_0,n341,_w_2242,n199,n170_0,n306,n188,_w_2011,_w_1816,_w_2279,n25,_w_2246,n310,n387_0,_w_2225,n271_1,n356_0,n276_1,_w_1424,n311,a_5__0,n123_0,n109_1,_w_1416,a_7__2,n194_1,n51,n316,_w_2219,n358,_w_2081,b_3__6,_w_2104,_w_2053,_w_2493,_w_2285,n319,b_7__3,n260,_w_1942,_w_2185,n29_1,n307_0,n208,b_6__2,n226_0,n325,n253_0,n327,n152_0,n53_0,n244_1,_w_2214,_w_1903,n329,_w_2444,n186,_w_1931,n330,n334,_w_1985,n111_0,n36_1,n335,n425_1,n434_1,n325_0,_w_1338,n409_0,n336,b_0__1,_w_2076,n274_1,a_7__7,n45_1,n237_0,n437_1,n67,n338,n212,a_7__8,n420,n339,_w_2345,n121_0,_w_2033,n343,n355_0,_w_2132,n47_0,_w_2448,n422,n54_1,n238_1,n92,n248,n356,_w_2310,n46_0,n177,n282_0,_w_1426,_w_2251,n424,n207,n359,n434,_w_2255,b_4__0,n230_1,b_0__2,n360,b_0__10,n181,n85,n344,n364,n30_1,n231,n85_1,_w_2227,n393,n100,_w_2506,n81_0,n351,n99,n35,n376,n78,n264,n379,n97_0,n255,n277_1,_w_1990,n237,n114,n149_0,n381,_w_2210,n383,_w_1706,n318,_w_1506,n387,n389,_w_1646,n395,a_6__1,n368_0,_w_2051,_w_1690,n423_1,n406,n123_1,n379_1,_w_1579,_w_2037,n149_1,_w_1739,n28_1,b_7__1,n412,n304,n216_0,_w_2521,n421,a_0__10,b_6__9,n380,_w_2075,_w_1813,_w_2327,_w_2413,n43_0,n184_1,_w_2069,_w_1776,n90,n428,n330_1,n192_1,_w_1298,_w_1429,_w_1661,n409,n429,_w_2233,n441,_w_1495,n234,n56_0,_w_2187,n439,n339_1,n435_0,n277_0,n226,_w_2293,_w_2341,_w_2083,_w_1869,n453,_w_2156,n439_0,n438_1,n26_1,n129,n429_1,a_4__4,n410_0,n204,n248_1,n406_0,n49_1,n302,_w_1723,_w_2348,n406_1,n73,n427_1,n319_0,n401_0,n18_1,n37_0,n146,n339_0,n191,n98,n242,_w_2263,n399,n116,_w_1638,_w_1832,_w_2408,n387_1,n232,n379_0,n112_1,b_6__10,_w_2056,_w_2356,n151,n366_1,n164,_w_1316,n340,n329_0,_w_2231,a_7__0,n258_0,a_1__6,_w_2318,n357_0,_w_2192,n402,b_4__2,n107,n355_1,n345_1,_w_1472,n165,_w_1889,a_5__4,n345_2,n33,_w_2311,n183,n345_3,_w_1289,n389_0,n224,_w_2355,n338_0,n366_0,n337_0,n357_1,n337_1,_w_1354,b_5__1,b_3__5,n336_1,n58_0,n335_1,a_7__6,n332_0,n325_1,_w_2427,_w_1804,_w_2019,n204_1,n204_2,_w_2545,_w_2314,n204_3,n48,n138_1,n158_1,n84_0,n240_1,n207_0,n251,n146_1,a_0__3,n143_0,_w_1684,n143_1,n419_0,_w_2116,n419_1,_w_1897,n350_1,_w_2330,_w_1548,n148_0,_w_1412,_w_1437,_w_1732,_w_1754,n148_1,n151_0,_w_2426,n151_1,n157_0,n430_1,n198_0,_w_2035,n396_0,n193_0,n160_0,n179_1,n326_0,n62_1,_w_1317,n62_3,n62_4,n162_0,n162_1,_w_1943,_w_1539,n163_0,n163_1,b_5__7,n194_0,n166_1,_w_2509,n158,_w_1854,n98_0,_w_2287,n98_1,_w_1374,n177_1,_w_1651,_w_2410,n178_0,_w_1958,n368_1,n181_0,n323_0,_w_1756,n181_1,n256_0,n256_1,n188_0,n17_0,_w_1791,n190_1,n191_0,n310_0,n191_1,n241,a_1__0,_w_1431,_w_2297,a_1__2,a_1__3,a_1__5,b_3__1,a_1__8,_w_1959,_w_2533,a_1__9,n232_0,a_1__10,n133,n193_1,a_1__11,n196_0,n196_1,_w_1307,_w_2141,n192_0,n231_0,n231_1,n203_0,n203_2,n353_0,_w_2393,n353_1,n19_1,n174_0,_w_2189,_w_1372,n215_0,n371_1,n215_1,n215_2,n108,_w_1819,n216_1,_w_2043,n220_1,n295_1,_w_1801,_w_2048,n222_0,n220_0,n226_1,n134_1,_w_1796,_w_2113,n239_0,n239_1,n228_0,_w_1965,n228_1,n230_0,n427_0,n84_2,n233,n241_0,n107_0,n76,n232_1,_w_1531,n235_0,n235_1,n342_0,n328,n342_1,n238_0,n431_0,n431_1,n146_0,_w_1545,n241_1,n241_2,_w_1292,_w_1293,_w_1294,_w_1689,n75_0,_w_1295,_w_1296,_w_1297,_w_1299,a_6__3,_w_1302,n162,_w_1303,_w_2045,_w_1308,n397,_w_1310,n302_1,_w_1311,_w_1312,n234_0,_w_1318,_w_1319,_w_1321,_w_1322,_w_2112,_w_1324,_w_2158,_w_1327,n308_1,_w_1330,_w_1332,_w_2152,_w_1333,_w_1344,_w_2349,_w_1598,_w_2294,_w_1334,_w_1336,_w_2526,_w_1807,_w_2059,_w_2321,n220,_w_1339,_w_1430,_w_1340,_w_1342,_w_2010,_w_1343,_w_2473,n86,_w_1345,_w_1346,_w_1347,_w_1736,_w_2108,n222_1,_w_1348,n203_3,_w_1351,_w_2466,_w_1352,_w_1734,a_7__10,_w_1384,_w_1355,_w_1358,_w_2001,n124_0,_w_1362,_w_1950,a_1__7,_w_1364,_w_1368,n370_1,_w_1369,_w_1370,_w_1454,_w_1705,_w_1371,_w_1373,_w_1376,_w_1678,_w_1377,_w_1378,n43_1,_w_2027,_w_1380,_w_1564,_w_1383,_w_1386,_w_1974,_w_2291,_w_1387,_w_1488,_w_2193,_w_1388,n72,_w_1640,_w_1389,a_3__5,_w_1390,_w_1391,_w_1515,_w_1995,_w_1392,_w_1395,_w_1396,_w_2213,_w_2528,n112_0,_w_1398,n41_1,_w_1399,_w_2173,_w_2029,_w_1400,_w_1402,_w_2292,_w_1405,_w_1406,_w_1407,_w_1409,n47,_w_1410,_w_1411,n17_1,_w_1413,_w_1415,_w_1419,_w_1656,_w_1587,_w_1425,_w_1427,_w_1428,n32,_w_2352,_w_1432,b_2__6,_w_1434,_w_1435,_w_2147,n256_2,_w_1961,_w_1438,_w_1648,_w_1439,_w_1305,_w_1440,_w_2061,_w_2077,_w_2510,_w_1337,_w_1441,_w_1442,n239,_w_1443,_w_1855,_w_1444,_w_1447,_w_1451,b_6__11,_w_1455,n383_1,_w_1458,_w_1459,_w_1463,_w_1466,_w_1600,_w_1469,_w_1470,_w_1471,_w_1474,_w_1478,_w_1288,_w_1479,_w_1809,_w_2399,_w_1480,n413,_w_1483,_w_2195,_w_1485,_w_1486,n381_1,_w_1806,_w_1489,_w_2175,n120,_w_1491,_w_1494,n115_1,_w_1497,_w_1499,_w_1500,_w_1692,n238,_w_1501,_w_2508,_w_1502,b_2__7,_w_1503,_w_2236,_w_1504,_w_1507,n351_0,_w_1509,n30_0,_w_1767,_w_1901,_w_1510,_w_1300,_w_1511,n81,_w_1513,_w_2516,_w_1516,_w_1498,_w_1520,_w_1522,_w_1831,_w_1526,_w_1683,_w_1528,_w_1544,_w_1534,n24_1,_w_1535,_w_1408,_w_1536,_w_1555,_w_1538,_w_1541,a_0__9,_w_1542,_w_2170,_w_2378,_w_2315,_w_1546,_w_1550,_w_1552,_w_1556,_w_1557,_w_2502,n363_0,_w_1558,_w_1559,n160,_w_2058,n365,_w_1561,_w_2184,_w_1562,_w_1563,_w_1645,n126,_w_1567,_w_1568,_w_1570,_w_1571,_w_1572,_w_1575,_w_2098,_w_1576,_w_1837,_w_1582,_w_1583,n316_0,_w_2085,_w_1584,_w_1833,n129_1,_w_1585,_w_2062,_w_2129,_w_1588,_w_1589,_w_1590,n414_0,_w_1592,_w_1593,_w_1597,_w_1599,_w_2420,_w_1601,_w_1769,_w_1603,_w_1608,_w_1866,_w_1609,_w_2333,_w_1610,n194,_w_1627,_w_1612,b_5__10,_w_1997,n150_1,_w_1613,n196,_w_1482,_w_1614,_w_1617,_w_1618,_w_1619,_w_1620,_w_1621,n322,_w_1626,_w_1629,_w_1630,n49,_w_2082,_w_1633,_w_1811,_w_1713,_w_1634,_w_2177,_w_1637,_w_1639,_w_2038,_w_1641,_w_1642,n59_1,_w_1602,_w_1643,_w_1331,_w_1652,_w_1653,_w_1365,_w_1655,n86_1,_w_2335,_w_1662,_w_2447,_w_2084,_w_1663,n124_1,n299,_w_1664,_w_1657,_w_1665,n207_1,_w_2012,_w_2028,_w_1668,_w_2252,_w_1673,_w_1674,_w_1676,_w_1679,_w_1680,_w_1681,n261,_w_1682,_w_1685,_w_1353,_w_1686,n361_1,_w_1687,_w_1688,_w_1695,_w_2562,_w_1696,n169,n63,_w_1514,_w_1697,_w_1966,_w_1698,_w_1700,_w_1701,_w_2479,n81_1,n293_1,_w_1702,_w_2127,n114_1,_w_2179,n318_0,b_3__8,_w_1707,_w_2136,_w_2180,_w_1708,_w_1543,n317,_w_1710,_w_1711,_w_1712,_w_1521,_w_1812,n290_1,_w_2093,n158_0,_w_1715,_w_1716,n100_0,n268_2,_w_1718,_w_1720,_w_1722,_w_1726,n205_0,_w_1938,b_3__2,_w_1727,_w_2354,_w_1731,n116_1,n160_1,_w_1733,n284_2,_w_1893,n54_0,_w_1735,_w_2277,_w_1737,_w_1740,_w_1742,_w_1533,_w_1745,_w_1963,_w_1751,_w_1753,n112,_w_2003,_w_1755,_w_2484,n276,_w_1876,_w_1757,n253,_w_1758,_w_1759,_w_1760,_w_1762,_w_1765,_w_1766,_w_1770,_w_1771,_w_1404,_w_1772,_w_1774,_w_1778,_w_1779,_w_2336,_w_1467,_w_1781,n347_0,_w_1581,_w_2206,_w_1782,_w_1669,_w_1783,n355,_w_2238,_w_1445,_w_1784,n426,_w_1873,_w_2054,_w_1785,a_2__1,_w_1787,_w_1789,_w_1792,n433,n199_0,_w_1794,_w_1797,_w_1799,n62_0,_w_1798,_w_1800,b_4__9,_w_1802,_w_1803,_w_1835,_w_1810,_w_1817,n373_1,_w_1818,n400_1,_w_1820,_w_1823,_w_1825,n330_0,_w_2283,n212_0,_w_1529,_w_1826,_w_1827,_w_1828,b_1__10,n94,_w_1829,_w_1887,_w_1838,_w_1839,_w_1304,_w_1840,a_4__0,n107_1,_w_1379,_w_1841,n373_0,_w_1844,_w_2415,_w_1846,a_3__0,_w_1574,_w_1848,n215,_w_2055,_w_1850,n291_1,n153,_w_1851,n166_0,_w_1852,_w_1857,_w_1862,_w_2068,_w_1622,_w_1863,n36,_w_1914,_w_2118,_w_1649,_w_1864,n83_1,_w_1867,_w_2142,_w_1871,_w_1872,_w_1874,_w_1875,n350_0,_w_1879,n262,_w_1393,_w_1880,_w_1881,n329_1,_w_1883,_w_1969,_w_2060,_w_1884,_w_1847,_w_1885,b_2__4,_w_1859,_w_1886,_w_1895,_w_1898,_w_2200,_w_1899,_w_1902,_w_1904,_w_1882,_w_1906,n250_1,_w_1752,_w_2089,_w_2216,_w_1908,_w_1909,n349,_w_1860,_w_1912,n411_1,_w_1913,_w_1915,_w_2544,_w_1919,_w_1921,_w_1923,_w_1924,_w_1925,_w_1926,_w_1933,_w_2456,_w_1935,_w_2247,_w_1750,_w_1936,_w_1900,_w_1939,_w_1971,n97_1,_w_1941,_w_1945,_w_2205,_w_1946,_w_1615,_w_1948,_w_2286,_w_1949,_w_2046,_w_1952,_w_1954,_w_1957,n251_1,_w_1960,_w_1964,n116_0,_w_2340,n136,_w_1968,_w_1973,_w_1616,_w_1975,_w_1977,_w_1979,_w_1980,n20,_w_2278,_w_2119,_w_1981,_w_1986,_w_2542,_w_1987,_w_1456,_w_1989,_w_2102,_w_1992,_w_1606,_w_1768,_w_1993,n385_0,_w_2222,_w_1999,_w_2000,_w_2002,_w_2005,n348,n179_0,_w_2006,_w_2007,n272,_w_2008,_w_2009,n271_0,_w_2013,n105,_w_2014,_w_1569,_w_2015,_w_2018,_w_2025,_w_2026,n225,_w_2030,_w_1490,_w_2031,_w_2032,a_6__0,_w_1951,_w_2036,_w_2040,b_2__8,_w_2041,_w_1611,_w_2044,_w_2049,_w_2050,_w_2063,_w_1930,_w_2066,_w_1650,_w_2072,_w_2017,_w_2087,_w_2073,_w_2261,_w_1976,_w_2074,_w_2080,n396_1,_w_2239,_w_2306,_w_2086,_w_2088,n417,_w_2090,b_2__10,_w_2092,_w_2094,_w_2153,_w_2095,_w_2096,n320,_w_2097,_w_2099,_w_2309,_w_2100,_w_1868,_w_2103,_w_2105,_w_2109,n325_2,_w_2110,_w_1605,_w_2111,_w_1890,_w_2114,n80,_w_2115,b_4__1,_w_2120,_w_2121,_w_2124,_w_2125,_w_2128,n210_0,_w_2130,n437,_w_2347,_w_2131,n384_0,_w_2133,_w_1397,_w_2052,_w_2253,_w_2137,_w_2140,_w_1594,_w_2143,_w_2144,_w_2145,n140_0,_w_1580,_w_2146,n117_1,_w_1460,_w_2154,_w_2022,_w_2161,_w_2165,_w_2500,n374,_w_2166,_w_2167,n39,_w_2171,_w_2172,_w_2176,_w_2182,n145,_w_2191,_w_2197,b_7__8,_w_2199,n31_0,_w_2207,_w_2304,_w_2208,_w_2215,_w_1719,_w_2217,n91_0,_w_2016,_w_2220,_w_1596,_w_2224,_w_2226,_w_2342,_w_1554,_w_2232,_w_2234,_w_2235,_w_2237,_w_2240,_w_2241,_w_2243,n323,_w_2245,_w_2250,_w_2254,_w_2256,_w_2258,_w_2259,_w_2260,_w_2265,_w_1853,_w_2267,_w_2268,n289,_w_2269,_w_1291,_w_1532,_w_2270,_w_2272,_w_1910,_w_2273,_w_2280,n326,_w_2282,_w_2284,_w_2295,_w_1916,_w_2296,_w_1644,_w_2299,_w_2300,_w_1591,_w_2301,_w_2302,_w_2303,n30,_w_2305,a_0__4,_w_2307,n361_0,_w_2308,_w_2316,_w_1492,_w_2317,_w_2319,_w_2320,_w_2323,_w_2324,_w_1537,_w_2328,_w_2331,_w_2334,_w_2556,_w_2337,_w_2338,_w_2138,_w_1505,_w_2339,_w_2343,_w_1530,_w_2353;

  bfr _b_2115(.a(_w_2570),.q(_w_2571));
  bfr _b_2113(.a(_w_2568),.q(_w_2569));
  bfr _b_2112(.a(_w_2567),.q(_w_2568));
  bfr _b_2111(.a(a_0_),.q(_w_2567));
  bfr _b_2110(.a(a_3_),.q(_w_2565));
  bfr _b_2109(.a(_w_2564),.q(_w_2553));
  bfr _b_2108(.a(_w_2563),.q(_w_2564));
  bfr _b_2107(.a(_w_2562),.q(_w_2563));
  bfr _b_2106(.a(_w_2561),.q(_w_2562));
  bfr _b_2101(.a(_w_2556),.q(_w_2557));
  bfr _b_2100(.a(_w_2555),.q(_w_2556));
  bfr _b_2099(.a(_w_2554),.q(_w_2555));
  bfr _b_2097(.a(_w_2552),.q(_w_2549));
  bfr _b_2093(.a(_w_2548),.q(_w_2541));
  bfr _b_2091(.a(_w_2546),.q(_w_2547));
  bfr _b_2090(.a(_w_2545),.q(_w_2546));
  bfr _b_2089(.a(_w_2544),.q(_w_2545));
  bfr _b_2088(.a(_w_2543),.q(_w_2544));
  bfr _b_2085(.a(a_5_),.q(_w_2540));
  bfr _b_2084(.a(_w_2539),.q(_w_2536));
  bfr _b_2083(.a(_w_2538),.q(_w_2539));
  bfr _b_2082(.a(_w_2537),.q(_w_2538));
  bfr _b_2080(.a(a_4_),.q(_w_2535));
  bfr _b_2076(.a(_w_2531),.q(_w_2532));
  bfr _b_2075(.a(_w_2530),.q(_w_2531));
  bfr _b_2074(.a(_w_2529),.q(_w_2530));
  bfr _b_2071(.a(_w_2526),.q(_w_2527));
  bfr _b_2068(.a(_w_2523),.q(_w_2524));
  bfr _b_2065(.a(b_7_),.q(_w_2521));
  bfr _b_2061(.a(_w_2516),.q(_w_2517));
  bfr _b_2060(.a(_w_2515),.q(_w_2516));
  bfr _b_2059(.a(a_1_),.q(_w_2515));
  bfr _b_2057(.a(_w_2512),.q(_w_2513));
  bfr _b_2055(.a(b_4_),.q(_w_2511));
  bfr _b_2052(.a(_w_2507),.q(_w_2508));
  bfr _b_2050(.a(_w_2505),.q(_w_2506));
  bfr _b_2049(.a(_w_2504),.q(n274_1));
  bfr _b_2047(.a(_w_2502),.q(_w_2503));
  bfr _b_2045(.a(_w_2500),.q(n195));
  bfr _b_2043(.a(_w_2498),.q(_w_2499));
  bfr _b_2042(.a(_w_2497),.q(_w_2498));
  bfr _b_2041(.a(_w_2496),.q(_w_2497));
  bfr _b_2039(.a(_w_2494),.q(n318_1));
  bfr _b_2034(.a(_w_2489),.q(n167));
  bfr _b_2030(.a(_w_2485),.q(_w_2486));
  bfr _b_2072(.a(_w_2527),.q(_w_2528));
  bfr _b_2029(.a(_w_2484),.q(_w_2485));
  bfr _b_2026(.a(_w_2481),.q(a_7__12));
  bfr _b_2024(.a(_w_2479),.q(n451));
  bfr _b_2020(.a(_w_2475),.q(_w_2476));
  bfr _b_2019(.a(_w_2474),.q(n373));
  bfr _b_2018(.a(_w_2473),.q(_w_2474));
  bfr _b_2027(.a(_w_2482),.q(n453));
  bfr _b_2016(.a(_w_2471),.q(_w_2472));
  bfr _b_2014(.a(_w_2469),.q(_w_2470));
  bfr _b_2013(.a(_w_2468),.q(_w_2469));
  bfr _b_2011(.a(_w_2466),.q(_w_2467));
  bfr _b_2007(.a(_w_2462),.q(s_7_));
  bfr _b_2005(.a(_w_2460),.q(_w_2461));
  bfr _b_2004(.a(_w_2459),.q(_w_2460));
  bfr _b_2002(.a(_w_2457),.q(_w_2458));
  bfr _b_2001(.a(_w_2456),.q(_w_2457));
  bfr _b_2000(.a(_w_2455),.q(_w_2456));
  bfr _b_1998(.a(_w_2453),.q(_w_2454));
  bfr _b_1997(.a(_w_2452),.q(_w_2453));
  bfr _b_1996(.a(_w_2451),.q(_w_2452));
  bfr _b_2058(.a(_w_2513),.q(_w_2510));
  bfr _b_1994(.a(_w_2449),.q(_w_2450));
  bfr _b_1993(.a(_w_2448),.q(_w_2449));
  bfr _b_1992(.a(_w_2447),.q(_w_2448));
  bfr _b_1991(.a(_w_2446),.q(_w_2447));
  bfr _b_1990(.a(_w_2445),.q(_w_2446));
  bfr _b_1987(.a(_w_2442),.q(_w_2443));
  bfr _b_1986(.a(_w_2441),.q(_w_2442));
  bfr _b_1985(.a(_w_2440),.q(_w_2441));
  bfr _b_1984(.a(_w_2439),.q(_w_2440));
  bfr _b_1983(.a(_w_2438),.q(_w_2439));
  bfr _b_1982(.a(_w_2437),.q(_w_2438));
  bfr _b_1981(.a(_w_2436),.q(_w_2437));
  bfr _b_1979(.a(_w_2434),.q(_w_2435));
  bfr _b_1977(.a(_w_2432),.q(_w_2433));
  bfr _b_2035(.a(_w_2490),.q(n417));
  bfr _b_1975(.a(_w_2430),.q(_w_2431));
  bfr _b_1974(.a(_w_2429),.q(_w_2430));
  bfr _b_1972(.a(_w_2427),.q(_w_2428));
  bfr _b_1971(.a(_w_2426),.q(_w_2427));
  bfr _b_1970(.a(_w_2425),.q(_w_2426));
  bfr _b_1968(.a(_w_2423),.q(_w_2424));
  bfr _b_1964(.a(_w_2419),.q(_w_2420));
  bfr _b_2102(.a(_w_2557),.q(_w_2558));
  bfr _b_1958(.a(_w_2413),.q(_w_2414));
  bfr _b_1957(.a(_w_2412),.q(_w_2413));
  bfr _b_1952(.a(_w_2407),.q(n424));
  bfr _b_1951(.a(_w_2406),.q(_w_2407));
  bfr _b_1950(.a(_w_2405),.q(_w_2406));
  bfr _b_1949(.a(_w_2404),.q(_w_2405));
  bfr _b_1948(.a(_w_2403),.q(_w_2404));
  bfr _b_1946(.a(_w_2401),.q(_w_2402));
  bfr _b_1944(.a(_w_2399),.q(_w_2400));
  bfr _b_1943(.a(_w_2398),.q(_w_2399));
  bfr _b_1937(.a(_w_2392),.q(_w_2393));
  bfr _b_1934(.a(_w_2389),.q(_w_2390));
  bfr _b_1933(.a(_w_2388),.q(_w_2389));
  bfr _b_1929(.a(_w_2384),.q(n420));
  bfr _b_1927(.a(_w_2382),.q(_w_2383));
  bfr _b_1926(.a(_w_2381),.q(_w_2382));
  bfr _b_1925(.a(_w_2380),.q(_w_2381));
  bfr _b_1924(.a(_w_2379),.q(_w_2380));
  bfr _b_1923(.a(_w_2378),.q(_w_2379));
  bfr _b_1922(.a(_w_2377),.q(n416));
  bfr _b_1919(.a(_w_2374),.q(_w_2375));
  bfr _b_1914(.a(_w_2369),.q(_w_2370));
  bfr _b_1913(.a(_w_2368),.q(_w_2369));
  bfr _b_1912(.a(_w_2367),.q(_w_2368));
  bfr _b_1910(.a(_w_2365),.q(_w_2366));
  bfr _b_1907(.a(_w_2362),.q(_w_2363));
  bfr _b_1906(.a(_w_2361),.q(_w_2362));
  bfr _b_2009(.a(_w_2464),.q(_w_2465));
  bfr _b_1905(.a(_w_2360),.q(_w_2361));
  bfr _b_1969(.a(_w_2424),.q(s_10_));
  bfr _b_1904(.a(_w_2359),.q(_w_2360));
  bfr _b_1903(.a(_w_2358),.q(_w_2359));
  bfr _b_1898(.a(_w_2353),.q(n414));
  bfr _b_1895(.a(_w_2350),.q(_w_2351));
  bfr _b_1893(.a(_w_2348),.q(_w_2349));
  bfr _b_1892(.a(_w_2347),.q(_w_2348));
  bfr _b_1891(.a(_w_2346),.q(_w_2347));
  bfr _b_1887(.a(_w_2342),.q(_w_2343));
  bfr _b_1881(.a(_w_2336),.q(_w_2337));
  bfr _b_1879(.a(_w_2334),.q(_w_2335));
  bfr _b_1878(.a(_w_2333),.q(_w_2334));
  bfr _b_1876(.a(_w_2331),.q(_w_2332));
  bfr _b_1869(.a(_w_2324),.q(n33));
  bfr _b_1868(.a(_w_2323),.q(n392));
  bfr _b_1867(.a(_w_2322),.q(_w_2323));
  bfr _b_1866(.a(_w_2321),.q(_w_2322));
  bfr _b_1863(.a(_w_2318),.q(_w_2319));
  bfr _b_1861(.a(_w_2316),.q(_w_2317));
  bfr _b_1859(.a(_w_2314),.q(_w_2315));
  bfr _b_2056(.a(_w_2511),.q(_w_2512));
  bfr _b_1858(.a(_w_2313),.q(_w_2314));
  bfr _b_1857(.a(_w_2312),.q(_w_2313));
  bfr _b_1855(.a(_w_2310),.q(_w_2311));
  bfr _b_1854(.a(_w_2309),.q(_w_2310));
  bfr _b_1852(.a(_w_2307),.q(n406));
  bfr _b_2048(.a(_w_2503),.q(_w_2504));
  bfr _b_1850(.a(_w_2305),.q(_w_2306));
  bfr _b_1847(.a(_w_2302),.q(_w_2303));
  bfr _b_1846(.a(_w_2301),.q(n377));
  bfr _b_1844(.a(_w_2299),.q(_w_2300));
  bfr _b_1843(.a(_w_2298),.q(_w_2299));
  bfr _b_1842(.a(_w_2297),.q(_w_2298));
  bfr _b_1836(.a(_w_2291),.q(_w_2292));
  bfr _b_1833(.a(_w_2288),.q(_w_2289));
  bfr _b_1832(.a(_w_2287),.q(n372));
  bfr _b_1831(.a(_w_2286),.q(_w_2287));
  bfr _b_1829(.a(_w_2284),.q(b_6__5));
  bfr _b_1827(.a(_w_2282),.q(_w_2283));
  bfr _b_1825(.a(_w_2280),.q(_w_2281));
  bfr _b_1824(.a(_w_2279),.q(_w_2280));
  bfr _b_1823(.a(_w_2278),.q(_w_2279));
  bfr _b_1821(.a(_w_2276),.q(_w_2277));
  bfr _b_1819(.a(_w_2274),.q(_w_2275));
  bfr _b_1814(.a(_w_2269),.q(_w_2270));
  bfr _b_1813(.a(_w_2268),.q(_w_2269));
  bfr _b_1812(.a(_w_2267),.q(_w_2268));
  bfr _b_1808(.a(_w_2263),.q(_w_2264));
  bfr _b_1976(.a(_w_2431),.q(_w_2432));
  bfr _b_1807(.a(_w_2262),.q(_w_2263));
  bfr _b_1884(.a(_w_2339),.q(_w_2340));
  bfr _b_1805(.a(_w_2260),.q(_w_2261));
  bfr _b_1804(.a(_w_2259),.q(_w_2260));
  bfr _b_1799(.a(_w_2254),.q(_w_2255));
  bfr _b_1794(.a(_w_2249),.q(_w_2250));
  bfr _b_1849(.a(_w_2304),.q(_w_2305));
  bfr _b_1793(.a(_w_2248),.q(_w_2249));
  bfr _b_1789(.a(_w_2244),.q(n359));
  bfr _b_1989(.a(_w_2444),.q(_w_2445));
  bfr _b_1788(.a(_w_2243),.q(a_6__13));
  bfr _b_1787(.a(_w_2242),.q(_w_2243));
  bfr _b_1786(.a(_w_2241),.q(_w_2242));
  bfr _b_1781(.a(_w_2236),.q(n352));
  bfr _b_1777(.a(_w_2232),.q(_w_2233));
  bfr _b_1774(.a(_w_2229),.q(_w_2230));
  bfr _b_1770(.a(_w_2225),.q(_w_2226));
  bfr _b_1768(.a(_w_2223),.q(n443));
  bfr _b_1767(.a(_w_2222),.q(n343));
  bfr _b_1763(.a(_w_2218),.q(_w_2219));
  bfr _b_1759(.a(_w_2214),.q(_w_2215));
  bfr _b_1920(.a(_w_2375),.q(_w_2376));
  bfr _b_1757(.a(_w_2212),.q(_w_2213));
  bfr _b_1755(.a(_w_2210),.q(s_4_));
  bfr _b_1752(.a(_w_2207),.q(_w_2208));
  bfr _b_1963(.a(_w_2418),.q(_w_2419));
  bfr _b_1750(.a(_w_2205),.q(_w_2206));
  bfr _b_1749(.a(_w_2204),.q(_w_2205));
  bfr _b_1748(.a(_w_2203),.q(_w_2204));
  bfr _b_1747(.a(_w_2202),.q(_w_2203));
  bfr _b_1745(.a(_w_2200),.q(_w_2201));
  bfr _b_1742(.a(_w_2197),.q(_w_2198));
  bfr _b_1839(.a(_w_2294),.q(_w_2295));
  bfr _b_1741(.a(_w_2196),.q(_w_2197));
  bfr _b_1740(.a(_w_2195),.q(_w_2196));
  bfr _b_1739(.a(_w_2194),.q(_w_2195));
  bfr _b_1736(.a(_w_2191),.q(_w_2192));
  bfr _b_1735(.a(_w_2190),.q(_w_2191));
  bfr _b_1732(.a(_w_2187),.q(_w_2188));
  bfr _b_1730(.a(_w_2185),.q(_w_2186));
  bfr _b_1725(.a(_w_2180),.q(_w_2181));
  bfr _b_1723(.a(_w_2178),.q(_w_2179));
  bfr _b_1722(.a(_w_2177),.q(_w_2178));
  bfr _b_1720(.a(_w_2175),.q(n328));
  bfr _b_1717(.a(_w_2172),.q(_w_2173));
  bfr _b_1714(.a(_w_2169),.q(_w_2170));
  bfr _b_1713(.a(_w_2168),.q(_w_2169));
  bfr _b_1712(.a(_w_2167),.q(_w_2168));
  bfr _b_1710(.a(_w_2165),.q(_w_2166));
  bfr _b_1709(.a(_w_2164),.q(n433));
  bfr _b_1738(.a(_w_2193),.q(_w_2194));
  bfr _b_1708(.a(_w_2163),.q(_w_2164));
  bfr _b_1705(.a(_w_2160),.q(_w_2161));
  bfr _b_1704(.a(_w_2159),.q(_w_2160));
  bfr _b_1703(.a(_w_2158),.q(_w_2159));
  bfr _b_1702(.a(_w_2157),.q(_w_2158));
  bfr _b_1701(.a(_w_2156),.q(_w_2157));
  bfr _b_1699(.a(_w_2154),.q(_w_2155));
  bfr _b_2053(.a(_w_2508),.q(n367_1));
  bfr _b_1696(.a(_w_2151),.q(_w_2152));
  bfr _b_1692(.a(_w_2147),.q(n323));
  bfr _b_2119(.a(_w_2574),.q(_w_2566));
  bfr _b_1691(.a(_w_2146),.q(_w_2147));
  bfr _b_1689(.a(_w_2144),.q(_w_2145));
  bfr _b_1688(.a(_w_2143),.q(_w_2144));
  bfr _b_1687(.a(_w_2142),.q(_w_2143));
  bfr _b_1686(.a(_w_2141),.q(_w_2142));
  bfr _b_1684(.a(_w_2139),.q(_w_2140));
  bfr _b_1681(.a(_w_2136),.q(n302_1));
  bfr _b_1680(.a(_w_2135),.q(_w_2136));
  bfr _b_1679(.a(_w_2134),.q(_w_2135));
  bfr _b_1677(.a(_w_2132),.q(n37));
  bfr _b_1988(.a(_w_2443),.q(_w_2444));
  bfr _b_1672(.a(_w_2127),.q(n319));
  bfr _b_1671(.a(_w_2126),.q(n398_1));
  bfr _b_2104(.a(_w_2559),.q(_w_2560));
  bfr _b_1874(.a(_w_2329),.q(_w_2330));
  bfr _b_1670(.a(_w_2125),.q(_w_2126));
  bfr _b_2094(.a(b_3_),.q(_w_2550));
  bfr _b_1666(.a(_w_2121),.q(_w_2122));
  bfr _b_1664(.a(_w_2119),.q(_w_2120));
  bfr _b_1658(.a(_w_2113),.q(_w_2114));
  bfr _b_1657(.a(_w_2112),.q(_w_2113));
  bfr _b_1938(.a(_w_2393),.q(_w_2394));
  bfr _b_1656(.a(_w_2111),.q(_w_2112));
  bfr _b_1651(.a(_w_2106),.q(_w_2107));
  bfr _b_1649(.a(_w_2104),.q(_w_2105));
  bfr _b_1648(.a(_w_2103),.q(_w_2104));
  bfr _b_1646(.a(_w_2101),.q(n127));
  bfr _b_1645(.a(_w_2100),.q(n362));
  bfr _b_1641(.a(_w_2096),.q(_w_2097));
  bfr _b_1640(.a(_w_2095),.q(n309));
  bfr _b_1638(.a(_w_2093),.q(_w_2094));
  bfr _b_1900(.a(_w_2355),.q(_w_2356));
  bfr _b_1728(.a(_w_2183),.q(_w_2184));
  bfr _b_1634(.a(_w_2089),.q(_w_2090));
  bfr _b_1632(.a(_w_2087),.q(n219));
  bfr _b_1631(.a(_w_2086),.q(n168_1));
  bfr _b_1630(.a(_w_2085),.q(_w_2086));
  bfr _b_1629(.a(_w_2084),.q(_w_2085));
  bfr _b_1628(.a(_w_2083),.q(_w_2084));
  bfr _b_1637(.a(_w_2092),.q(_w_2093));
  bfr _b_1627(.a(_w_2082),.q(_w_2083));
  bfr _b_1625(.a(_w_2080),.q(_w_2081));
  bfr _b_1624(.a(_w_2079),.q(_w_2080));
  bfr _b_1623(.a(_w_2078),.q(_w_2079));
  bfr _b_1621(.a(_w_2076),.q(n299));
  bfr _b_1620(.a(_w_2075),.q(s_2_));
  bfr _b_1618(.a(_w_2073),.q(_w_2074));
  bfr _b_1616(.a(_w_2071),.q(_w_2072));
  bfr _b_1614(.a(_w_2069),.q(_w_2070));
  bfr _b_1611(.a(_w_2066),.q(_w_2067));
  bfr _b_1610(.a(_w_2065),.q(_w_2066));
  bfr _b_1609(.a(_w_2064),.q(_w_2065));
  bfr _b_1894(.a(_w_2349),.q(_w_2350));
  bfr _b_1607(.a(_w_2062),.q(_w_2063));
  bfr _b_1603(.a(_w_2058),.q(_w_2059));
  bfr _b_1597(.a(_w_2052),.q(_w_2053));
  bfr _b_1595(.a(_w_2050),.q(_w_2051));
  bfr _b_1594(.a(_w_2049),.q(_w_2050));
  bfr _b_1593(.a(_w_2048),.q(_w_2049));
  bfr _b_1853(.a(_w_2308),.q(_w_2309));
  bfr _b_1591(.a(_w_2046),.q(_w_2047));
  bfr _b_1590(.a(_w_2045),.q(_w_2046));
  bfr _b_1588(.a(_w_2043),.q(_w_2044));
  bfr _b_1773(.a(_w_2228),.q(_w_2229));
  bfr _b_1587(.a(_w_2042),.q(_w_2043));
  bfr _b_1586(.a(_w_2041),.q(_w_2042));
  bfr _b_1584(.a(_w_2039),.q(_w_2040));
  bfr _b_1583(.a(_w_2038),.q(_w_2039));
  bfr _b_1582(.a(_w_2037),.q(_w_2038));
  bfr _b_1580(.a(_w_2035),.q(n389_1));
  bfr _b_1579(.a(_w_2034),.q(_w_2035));
  bfr _b_1578(.a(_w_2033),.q(n292));
  bfr _b_1577(.a(_w_2032),.q(n290));
  bfr _b_1575(.a(_w_2030),.q(_w_2031));
  bfr _b_1574(.a(_w_2029),.q(_w_2030));
  bfr _b_1573(.a(_w_2028),.q(_w_2029));
  bfr _b_1569(.a(_w_2024),.q(n25_1));
  bfr _b_1568(.a(_w_2023),.q(_w_2024));
  bfr _b_1567(.a(_w_2022),.q(_w_2023));
  bfr _b_1566(.a(_w_2021),.q(_w_2022));
  bfr _b_1565(.a(_w_2020),.q(n308));
  bfr _b_1562(.a(_w_2017),.q(_w_2018));
  bfr _b_2066(.a(_w_2521),.q(_w_2522));
  bfr _b_1561(.a(_w_2016),.q(_w_2017));
  bfr _b_1652(.a(_w_2107),.q(_w_2108));
  bfr _b_1560(.a(_w_2015),.q(_w_2016));
  bfr _b_1559(.a(_w_2014),.q(_w_2015));
  bfr _b_1556(.a(_w_2011),.q(n151_1));
  bfr _b_1555(.a(_w_2010),.q(_w_2011));
  bfr _b_1962(.a(_w_2417),.q(_w_2418));
  bfr _b_1945(.a(_w_2400),.q(_w_2401));
  bfr _b_1605(.a(_w_2060),.q(_w_2061));
  bfr _b_1554(.a(_w_2009),.q(_w_2010));
  bfr _b_1917(.a(_w_2372),.q(_w_2373));
  bfr _b_1841(.a(_w_2296),.q(_w_2297));
  bfr _b_1553(.a(_w_2008),.q(_w_2009));
  bfr _b_2028(.a(_w_2483),.q(n42));
  bfr _b_1871(.a(_w_2326),.q(n413));
  bfr _b_1551(.a(_w_2006),.q(n19));
  bfr _b_1550(.a(_w_2005),.q(_w_2006));
  bfr _b_1547(.a(_w_2002),.q(_w_2003));
  bfr _b_1546(.a(_w_2001),.q(_w_2002));
  bfr _b_1545(.a(_w_2000),.q(_w_2001));
  bfr _b_1633(.a(_w_2088),.q(_w_2089));
  bfr _b_1544(.a(_w_1999),.q(n132));
  bfr _b_1540(.a(_w_1995),.q(s_11_));
  bfr _b_1604(.a(_w_2059),.q(_w_2060));
  bfr _b_1539(.a(_w_1994),.q(_w_1995));
  bfr _b_1690(.a(_w_2145),.q(_w_2146));
  bfr _b_1537(.a(_w_1992),.q(_w_1993));
  bfr _b_1536(.a(_w_1991),.q(_w_1992));
  bfr _b_1535(.a(_w_1990),.q(_w_1991));
  bfr _b_1534(.a(_w_1989),.q(_w_1990));
  bfr _b_1533(.a(_w_1988),.q(_w_1989));
  bfr _b_1541(.a(_w_1996),.q(n187));
  bfr _b_1528(.a(_w_1983),.q(n296));
  bfr _b_1526(.a(_w_1981),.q(_w_1982));
  bfr _b_1524(.a(_w_1979),.q(a_1__2));
  bfr _b_1523(.a(_w_1978),.q(_w_1979));
  bfr _b_1522(.a(_w_1977),.q(_w_1978));
  bfr _b_1521(.a(_w_1976),.q(n445));
  bfr _b_1520(.a(_w_1975),.q(n118));
  bfr _b_1519(.a(_w_1974),.q(n234));
  bfr _b_1516(.a(_w_1971),.q(_w_1972));
  bfr _b_2086(.a(b_5_),.q(_w_2542));
  bfr _b_1513(.a(_w_1968),.q(_w_1969));
  bfr _b_1511(.a(_w_1966),.q(n106));
  bfr _b_1956(.a(_w_2411),.q(_w_2412));
  bfr _b_1510(.a(_w_1965),.q(n282_1));
  bfr _b_2032(.a(_w_2487),.q(n351_1));
  bfr _b_1782(.a(_w_2237),.q(n354));
  bfr _b_1507(.a(_w_1962),.q(n32));
  bfr _b_1506(.a(_w_1961),.q(_w_1962));
  bfr _b_1504(.a(_w_1959),.q(_w_1960));
  bfr _b_1503(.a(_w_1958),.q(_w_1959));
  bfr _b_1502(.a(_w_1957),.q(_w_1958));
  bfr _b_1883(.a(_w_2338),.q(_w_2339));
  bfr _b_1499(.a(_w_1954),.q(_w_1955));
  bfr _b_1497(.a(_w_1952),.q(n199_1));
  bfr _b_1496(.a(_w_1951),.q(_w_1952));
  bfr _b_1493(.a(_w_1948),.q(a_7__3));
  bfr _b_1491(.a(_w_1946),.q(n80));
  bfr _b_1911(.a(_w_2366),.q(_w_2367));
  bfr _b_1483(.a(_w_1938),.q(_w_1939));
  bfr _b_1480(.a(_w_1935),.q(_w_1936));
  bfr _b_1479(.a(_w_1934),.q(_w_1935));
  bfr _b_1475(.a(_w_1930),.q(_w_1931));
  bfr _b_1474(.a(_w_1929),.q(_w_1930));
  bfr _b_1472(.a(_w_1927),.q(_w_1928));
  bfr _b_1470(.a(_w_1925),.q(n270));
  bfr _b_1468(.a(_w_1923),.q(_w_1924));
  bfr _b_1467(.a(_w_1922),.q(_w_1923));
  bfr _b_1734(.a(_w_2189),.q(_w_2190));
  bfr _b_1466(.a(_w_1921),.q(_w_1922));
  bfr _b_1465(.a(_w_1920),.q(_w_1921));
  bfr _b_1826(.a(_w_2281),.q(_w_2282));
  bfr _b_1463(.a(_w_1918),.q(_w_1919));
  bfr _b_1462(.a(_w_1917),.q(n373_1));
  bfr _b_1459(.a(_w_1914),.q(_w_1915));
  bfr _b_1458(.a(_w_1913),.q(n242_1));
  bfr _b_1456(.a(_w_1911),.q(_w_1912));
  bfr _b_1455(.a(_w_1910),.q(_w_1911));
  bfr _b_1886(.a(_w_2341),.q(_w_2342));
  bfr _b_1454(.a(_w_1909),.q(a_2__8));
  bfr _b_1756(.a(_w_2211),.q(_w_2212));
  bfr _b_1453(.a(_w_1908),.q(_w_1909));
  bfr _b_1450(.a(_w_1905),.q(n139));
  bfr _b_1449(.a(_w_1904),.q(n161));
  bfr _b_1676(.a(_w_2131),.q(n320));
  bfr _b_1448(.a(_w_1903),.q(a_1__9));
  bfr _b_1446(.a(_w_1901),.q(_w_1902));
  bfr _b_1442(.a(_w_1897),.q(n339_1));
  bfr _b_1461(.a(_w_1916),.q(_w_1917));
  bfr _b_1441(.a(_w_1896),.q(_w_1897));
  bfr _b_1440(.a(_w_1895),.q(_w_1896));
  bfr _b_1585(.a(_w_2040),.q(_w_2041));
  bfr _b_1431(.a(_w_1886),.q(n113));
  bfr _b_1430(.a(_w_1885),.q(n249));
  bfr _b_1429(.a(_w_1884),.q(n266));
  bfr _b_1427(.a(_w_1882),.q(_w_1883));
  bfr _b_1548(.a(_w_2003),.q(_w_2004));
  bfr _b_1424(.a(_w_1879),.q(_w_1880));
  bfr _b_1422(.a(_w_1877),.q(_w_1878));
  bfr _b_1419(.a(_w_1874),.q(_w_1875));
  bfr _b_1418(.a(_w_1873),.q(_w_1874));
  bfr _b_1417(.a(_w_1872),.q(_w_1873));
  bfr _b_1571(.a(_w_2026),.q(n236));
  bfr _b_1412(.a(_w_1867),.q(_w_1868));
  bfr _b_1410(.a(_w_1865),.q(_w_1866));
  bfr _b_1408(.a(_w_1863),.q(_w_1864));
  bfr _b_1407(.a(_w_1862),.q(_w_1863));
  bfr _b_1406(.a(_w_1861),.q(_w_1862));
  bfr _b_1795(.a(_w_2250),.q(_w_2251));
  bfr _b_1405(.a(_w_1860),.q(_w_1861));
  bfr _b_1635(.a(_w_2090),.q(_w_2091));
  bfr _b_1404(.a(_w_1859),.q(_w_1860));
  bfr _b_1403(.a(_w_1858),.q(_w_1859));
  bfr _b_1402(.a(_w_1857),.q(_w_1858));
  bfr _b_1674(.a(_w_2129),.q(_w_2130));
  bfr _b_1530(.a(_w_1985),.q(_w_1986));
  bfr _b_1401(.a(_w_1856),.q(_w_1857));
  bfr _b_1864(.a(_w_2319),.q(_w_2320));
  bfr _b_1399(.a(_w_1854),.q(_w_1855));
  bfr _b_1865(.a(_w_2320),.q(_w_2321));
  bfr _b_1398(.a(_w_1853),.q(_w_1854));
  bfr _b_1396(.a(_w_1851),.q(_w_1852));
  bfr _b_1391(.a(_w_1846),.q(_w_1847));
  bfr _b_1700(.a(_w_2155),.q(_w_2156));
  bfr _b_1388(.a(_w_1843),.q(_w_1844));
  bfr _b_1387(.a(_w_1842),.q(_w_1843));
  bfr _b_1477(.a(_w_1932),.q(n425_1));
  bfr _b_1385(.a(_w_1840),.q(_w_1841));
  bfr _b_1384(.a(_w_1839),.q(_w_1840));
  bfr _b_1381(.a(_w_1836),.q(_w_1837));
  bfr _b_1378(.a(_w_1833),.q(_w_1834));
  bfr _b_1377(.a(_w_1832),.q(_w_1833));
  bfr _b_1413(.a(_w_1868),.q(_w_1869));
  bfr _b_1375(.a(_w_1830),.q(n108));
  bfr _b_1374(.a(_w_1829),.q(n222));
  bfr _b_1371(.a(_w_1826),.q(_w_1827));
  bfr _b_1707(.a(_w_2162),.q(_w_2163));
  bfr _b_1369(.a(_w_1824),.q(_w_1825));
  bfr _b_1368(.a(_w_1823),.q(n63));
  bfr _b_2070(.a(_w_2525),.q(_w_2526));
  bfr _b_1367(.a(_w_1822),.q(n284_1));
  bfr _b_1365(.a(_w_1820),.q(_w_1821));
  bfr _b_1364(.a(_w_1819),.q(n22));
  bfr _b_1834(.a(_w_2289),.q(_w_2290));
  bfr _b_1359(.a(_w_1814),.q(n376));
  bfr _b_1358(.a(_w_1813),.q(_w_1814));
  bfr _b_1357(.a(_w_1812),.q(_w_1813));
  bfr _b_1356(.a(_w_1811),.q(_w_1812));
  bfr _b_1660(.a(_w_2115),.q(_w_2116));
  bfr _b_1355(.a(_w_1810),.q(_w_1811));
  bfr _b_1354(.a(_w_1809),.q(_w_1810));
  bfr _b_1351(.a(_w_1806),.q(_w_1807));
  bfr _b_1350(.a(_w_1805),.q(_w_1806));
  bfr _b_1349(.a(_w_1804),.q(_w_1805));
  bfr _b_1348(.a(_w_1803),.q(n405_1));
  bfr _b_1347(.a(_w_1802),.q(_w_1803));
  bfr _b_2021(.a(_w_2476),.q(_w_2477));
  bfr _b_1460(.a(_w_1915),.q(_w_1916));
  bfr _b_1345(.a(_w_1800),.q(_w_1801));
  bfr _b_1451(.a(_w_1906),.q(n77));
  bfr _b_1393(.a(_w_1848),.q(_w_1849));
  bfr _b_1343(.a(_w_1798),.q(n432));
  bfr _b_1626(.a(_w_2081),.q(_w_2082));
  bfr _b_1341(.a(_w_1796),.q(_w_1797));
  bfr _b_1337(.a(_w_1792),.q(n51));
  bfr _b_1336(.a(_w_1791),.q(n136));
  bfr _b_1335(.a(_w_1790),.q(_w_1791));
  bfr _b_1334(.a(_w_1789),.q(_w_1790));
  bfr _b_1488(.a(_w_1943),.q(_w_1944));
  bfr _b_1333(.a(_w_1788),.q(_w_1789));
  bfr _b_1329(.a(_w_1784),.q(n210_1));
  bfr _b_1328(.a(_w_1783),.q(_w_1784));
  bfr _b_1810(.a(_w_2265),.q(_w_2266));
  bfr _b_1669(.a(_w_2124),.q(_w_2125));
  bfr _b_1332(.a(_w_1787),.q(n141));
  bfr _b_1322(.a(_w_1777),.q(_w_1778));
  bfr _b_1321(.a(_w_1776),.q(_w_1777));
  bfr _b_1899(.a(_w_2354),.q(n415));
  bfr _b_1320(.a(_w_1775),.q(_w_1776));
  bfr _b_1525(.a(_w_1980),.q(n125));
  bfr _b_1319(.a(_w_1774),.q(_w_1775));
  bfr _b_1897(.a(_w_2352),.q(_w_2353));
  bfr _b_1314(.a(_w_1769),.q(_w_1770));
  bfr _b_2006(.a(_w_2461),.q(_w_2462));
  bfr _b_1312(.a(_w_1767),.q(_w_1768));
  bfr _b_1397(.a(_w_1852),.q(_w_1853));
  bfr _b_1311(.a(_w_1766),.q(_w_1767));
  bfr _b_1890(.a(_w_2345),.q(_w_2346));
  bfr _b_1307(.a(_w_1762),.q(_w_1763));
  bfr _b_1306(.a(_w_1761),.q(_w_1762));
  bfr _b_1305(.a(_w_1760),.q(_w_1761));
  bfr _b_1304(.a(_w_1759),.q(_w_1760));
  bfr _b_1303(.a(_w_1758),.q(_w_1759));
  bfr _b_1302(.a(_w_1757),.q(_w_1758));
  bfr _b_1301(.a(_w_1756),.q(_w_1757));
  bfr _b_2116(.a(_w_2571),.q(_w_2572));
  bfr _b_1300(.a(_w_1755),.q(_w_1756));
  bfr _b_1818(.a(_w_2273),.q(_w_2274));
  bfr _b_1298(.a(_w_1753),.q(_w_1754));
  bfr _b_1297(.a(_w_1752),.q(_w_1753));
  bfr _b_1295(.a(_w_1750),.q(_w_1751));
  bfr _b_1294(.a(_w_1749),.q(_w_1750));
  bfr _b_1292(.a(_w_1747),.q(_w_1748));
  bfr _b_1654(.a(_w_2109),.q(_w_2110));
  bfr _b_1291(.a(_w_1746),.q(_w_1747));
  bfr _b_1290(.a(_w_1745),.q(_w_1746));
  bfr _b_1289(.a(_w_1744),.q(_w_1745));
  bfr _b_1514(.a(_w_1969),.q(_w_1970));
  bfr _b_1287(.a(_w_1742),.q(_w_1743));
  bfr _b_1966(.a(_w_2421),.q(_w_2422));
  bfr _b_1286(.a(_w_1741),.q(_w_1742));
  bfr _b_1283(.a(_w_1738),.q(a_4__2));
  bfr _b_1282(.a(_w_1737),.q(_w_1738));
  bfr _b_1279(.a(_w_1734),.q(_w_1735));
  bfr _b_1276(.a(_w_1731),.q(a_6__3));
  bfr _b_1274(.a(_w_1729),.q(_w_1730));
  bfr _b_1278(.a(_w_1733),.q(n393));
  bfr _b_1272(.a(_w_1727),.q(_w_1728));
  bfr _b_1683(.a(_w_2138),.q(_w_2139));
  bfr _b_1268(.a(_w_1723),.q(_w_1724));
  bfr _b_1277(.a(_w_1732),.q(_w_1733));
  bfr _b_1267(.a(_w_1722),.q(s_3_));
  bfr _b_1978(.a(_w_2433),.q(_w_2434));
  bfr _b_1264(.a(_w_1719),.q(_w_1720));
  bfr _b_1258(.a(_w_1713),.q(_w_1714));
  bfr _b_1256(.a(_w_1711),.q(_w_1712));
  bfr _b_1255(.a(_w_1710),.q(_w_1711));
  bfr _b_1251(.a(_w_1706),.q(_w_1707));
  bfr _b_1250(.a(_w_1705),.q(_w_1706));
  bfr _b_1249(.a(_w_1704),.q(_w_1705));
  bfr _b_1901(.a(_w_2356),.q(_w_2357));
  bfr _b_1248(.a(_w_1703),.q(_w_1704));
  bfr _b_1771(.a(_w_2226),.q(b_1__7));
  bfr _b_1372(.a(_w_1827),.q(n179));
  bfr _b_1246(.a(_w_1701),.q(_w_1702));
  bfr _b_1242(.a(_w_1697),.q(_w_1698));
  bfr _b_1241(.a(_w_1696),.q(_w_1697));
  bfr _b_1239(.a(_w_1694),.q(_w_1695));
  bfr _b_1494(.a(_w_1949),.q(_w_1950));
  bfr _b_1238(.a(_w_1693),.q(_w_1694));
  bfr _b_1324(.a(_w_1779),.q(_w_1780));
  bfr _b_1235(.a(_w_1690),.q(_w_1691));
  bfr _b_1234(.a(_w_1689),.q(_w_1690));
  bfr _b_1233(.a(_w_1688),.q(_w_1689));
  bfr _b_1361(.a(_w_1816),.q(n308_1));
  bfr _b_1232(.a(_w_1687),.q(_w_1688));
  bfr _b_1608(.a(_w_2063),.q(_w_2064));
  bfr _b_1231(.a(_w_1686),.q(_w_1687));
  bfr _b_1230(.a(_w_1685),.q(n428));
  bfr _b_1229(.a(_w_1684),.q(n306));
  bfr _b_1228(.a(_w_1683),.q(a_4__10));
  bfr _b_1227(.a(_w_1682),.q(_w_1683));
  bfr _b_1225(.a(_w_1680),.q(_w_1681));
  bfr _b_1224(.a(_w_1679),.q(n169));
  bfr _b_1222(.a(_w_1677),.q(_w_1678));
  bfr _b_1221(.a(_w_1676),.q(n426));
  bfr _b_1806(.a(_w_2261),.q(_w_2262));
  bfr _b_1598(.a(_w_2053),.q(_w_2054));
  bfr _b_1270(.a(_w_1725),.q(n153_3));
  bfr _b_1263(.a(_w_1718),.q(_w_1719));
  bfr _b_1220(.a(_w_1675),.q(n252));
  bfr _b_1219(.a(_w_1674),.q(n180));
  bfr _b_1443(.a(_w_1898),.q(n183));
  bfr _b_1216(.a(_w_1671),.q(_w_1672));
  bfr _b_1942(.a(_w_2397),.q(_w_2398));
  bfr _b_1213(.a(_w_1668),.q(n185));
  bfr _b_1265(.a(_w_1720),.q(_w_1721));
  bfr _b_1212(.a(_w_1667),.q(n189));
  bfr _b_1211(.a(_w_1666),.q(n202));
  bfr _b_1207(.a(_w_1662),.q(_w_1663));
  bfr _b_1206(.a(_w_1661),.q(_w_1662));
  bfr _b_1205(.a(_w_1660),.q(n82));
  bfr _b_1482(.a(_w_1937),.q(n176));
  bfr _b_1203(.a(_w_1658),.q(n253));
  bfr _b_1615(.a(_w_2070),.q(_w_2071));
  bfr _b_1200(.a(_w_1655),.q(n211));
  bfr _b_1549(.a(_w_2004),.q(_w_2005));
  bfr _b_1199(.a(_w_1654),.q(n382));
  bfr _b_1198(.a(_w_1653),.q(n217));
  bfr _b_1196(.a(_w_1651),.q(n229));
  bfr _b_1194(.a(_w_1649),.q(n224));
  bfr _b_1916(.a(_w_2371),.q(_w_2372));
  bfr _b_1775(.a(_w_2230),.q(_w_2231));
  bfr _b_1193(.a(_w_1648),.q(_w_1649));
  bfr _b_1995(.a(_w_2450),.q(_w_2451));
  bfr _b_1192(.a(_w_1647),.q(_w_1648));
  bfr _b_1191(.a(_w_1646),.q(_w_1647));
  bfr _b_1190(.a(_w_1645),.q(_w_1646));
  bfr _b_1931(.a(_w_2386),.q(n429));
  bfr _b_1189(.a(_w_1644),.q(_w_1645));
  bfr _b_1790(.a(_w_2245),.q(n365));
  bfr _b_1188(.a(_w_1643),.q(_w_1644));
  bfr _b_1187(.a(_w_1642),.q(_w_1643));
  bfr _b_1389(.a(_w_1844),.q(_w_1845));
  bfr _b_1183(.a(_w_1638),.q(n20));
  bfr _b_1180(.a(_w_1635),.q(_w_1636));
  bfr _b_1798(.a(_w_2253),.q(_w_2254));
  bfr _b_1179(.a(_w_1634),.q(_w_1635));
  bfr _b_1177(.a(_w_1632),.q(_w_1633));
  bfr _b_1176(.a(_w_1631),.q(_w_1632));
  bfr _b_1175(.a(_w_1630),.q(n247));
  bfr _b_1174(.a(_w_1629),.q(n449));
  bfr _b_1173(.a(_w_1628),.q(s_6_));
  bfr _b_1171(.a(_w_1626),.q(_w_1627));
  bfr _b_1169(.a(_w_1624),.q(_w_1625));
  bfr _b_1168(.a(_w_1623),.q(_w_1624));
  bfr _b_1167(.a(_w_1622),.q(_w_1623));
  bfr _b_1421(.a(_w_1876),.q(_w_1877));
  bfr _b_1164(.a(_w_1619),.q(_w_1620));
  bfr _b_1163(.a(_w_1618),.q(_w_1619));
  bfr _b_1716(.a(_w_2171),.q(_w_2172));
  bfr _b_1162(.a(_w_1617),.q(_w_1618));
  bfr _b_1159(.a(_w_1614),.q(_w_1615));
  bfr _b_1158(.a(_w_1613),.q(_w_1614));
  bfr _b_1156(.a(_w_1611),.q(_w_1612));
  bfr _b_1154(.a(_w_1609),.q(_w_1610));
  bfr _b_1153(.a(_w_1608),.q(_w_1609));
  bfr _b_1150(.a(_w_1605),.q(_w_1606));
  bfr _b_1148(.a(_w_1603),.q(_w_1604));
  bfr _b_1147(.a(_w_1602),.q(_w_1603));
  bfr _b_1146(.a(_w_1601),.q(_w_1602));
  bfr _b_1144(.a(_w_1599),.q(_w_1600));
  bfr _b_2064(.a(a_2_),.q(_w_2519));
  bfr _b_1142(.a(_w_1597),.q(n233));
  bfr _b_1141(.a(_w_1596),.q(n243));
  bfr _b_1140(.a(_w_1595),.q(n262));
  bfr _b_1138(.a(_w_1593),.q(_w_1594));
  bfr _b_1137(.a(_w_1592),.q(_w_1593));
  bfr _b_1136(.a(_w_1591),.q(_w_1592));
  bfr _b_2067(.a(_w_2522),.q(_w_2523));
  bfr _b_1133(.a(_w_1588),.q(_w_1589));
  bfr _b_1132(.a(_w_1587),.q(_w_1588));
  bfr _b_1293(.a(_w_1748),.q(_w_1749));
  bfr _b_1131(.a(_w_1586),.q(_w_1587));
  bfr _b_1129(.a(_w_1584),.q(_w_1585));
  bfr _b_1128(.a(_w_1583),.q(_w_1584));
  bfr _b_1127(.a(_w_1582),.q(_w_1583));
  bfr _b_1126(.a(_w_1581),.q(_w_1582));
  bfr _b_1125(.a(_w_1580),.q(_w_1581));
  bfr _b_1124(.a(_w_1579),.q(_w_1580));
  bfr _b_1160(.a(_w_1615),.q(_w_1616));
  bfr _b_1122(.a(_w_1577),.q(_w_1578));
  bfr _b_1121(.a(_w_1576),.q(_w_1577));
  bfr _b_1120(.a(_w_1575),.q(_w_1576));
  bfr _b_1119(.a(_w_1574),.q(_w_1575));
  bfr _b_1118(.a(_w_1573),.q(_w_1574));
  bfr _b_1776(.a(_w_2231),.q(_w_2232));
  bfr _b_1116(.a(_w_1571),.q(n386));
  bfr _b_1114(.a(_w_1569),.q(n60));
  bfr _b_1113(.a(_w_1568),.q(s_5_));
  bfr _b_1111(.a(_w_1566),.q(_w_1567));
  bfr _b_1110(.a(_w_1565),.q(_w_1566));
  bfr _b_1109(.a(_w_1564),.q(_w_1565));
  spl2 g34_s_0(.a(n34),.q0(n34_0),.q1(n34_1));
  bfr _b_1261(.a(_w_1716),.q(_w_1717));
  bfr _b_872(.a(_w_1327),.q(_w_1328));
  spl2 g400_s_0(.a(n400),.q0(n400_0),.q1(n400_1));
  and_bb g281(.a(a_5__7),.b(b_4__8),.q(n281));
  and_bb g40(.a(a_4__3),.b(b_3__2),.q(n40));
  bfr _b_1428(.a(_w_1883),.q(s_0_));
  bfr _b_1376(.a(_w_1831),.q(n407));
  bfr _b_1039(.a(_w_1494),.q(n227_1));
  spl2 g110_s_0(.a(n110),.q0(n110_0),.q1(n110_1));
  bfr _b_1967(.a(_w_2422),.q(_w_2423));
  spl2 g248_s_0(.a(n248),.q0(n248_0),.q1(n248_1));
  and_bi g34(.a(n33),.b(n31_0),.q(n34));
  spl2 g115_s_0(.a(n115),.q0(n115_0),.q1(n115_1));
  and_bi g97(.a(n96),.b(n93_0),.q(n97));
  spl3L g268_s_0(.a(n268),.q0(n268_0),.q1(n268_1),.q2(n268_2));
  bfr _b_2036(.a(_w_2491),.q(_w_2492));
  spl2 g367_s_0(.a(n367),.q0(n367_0),.q1(_w_2505));
  spl2 g273_s_0(.a(n273),.q0(n273_0),.q1(n273_1));
  and_bi g237(.a(n236),.b(n235_0),.q(n237));
  spl2 g279_s_0(.a(n279),.q0(n279_0),.q1(n279_1));
  spl2 g285_s_0(.a(n285),.q0(n285_0),.q1(_w_2496));
  spl2 g345_s_1(.a(n345_1),.q0(n345_2),.q1(n345_3));
  bfr _b_924(.a(_w_1379),.q(b_3__0));
  spl2 g294_s_0(.a(n294),.q0(n294_0),.q1(n294_1));
  spl2 g371_s_0(.a(n371),.q0(n371_0),.q1(n371_1));
  spl2 g372_s_0(.a(n372),.q0(n372_0),.q1(n372_1));
  bfr _b_1762(.a(_w_2217),.q(n329));
  or_bb g135(.a(n133_1),.b(n36_1),.q(_w_2495));
  bfr _b_1161(.a(_w_1616),.q(_w_1617));
  spl2 g408_s_0(.a(n408),.q0(n408_0),.q1(n408_1));
  bfr _b_1339(.a(_w_1794),.q(_w_1795));
  and_bi g58(.a(n57),.b(n56_0),.q(n58));
  bfr _b_908(.a(_w_1363),.q(_w_1364));
  bfr _b_1098(.a(_w_1553),.q(_w_1554));
  bfr _b_2038(.a(_w_2493),.q(_w_2494));
  bfr _b_1373(.a(_w_1828),.q(_w_1829));
  spl2 g423_s_0(.a(n423),.q0(n423_0),.q1(n423_1));
  spl2 g274_s_0(.a(n274),.q0(n274_0),.q1(_w_2501));
  and_bb g291(.a(n289_0),.b(n290_0),.q(n291));
  bfr _b_1313(.a(_w_1768),.q(_w_1769));
  and_bb g241(.a(n222_0),.b(n240_0),.q(n241));
  bfr _b_1471(.a(_w_1926),.q(_w_1927));
  spl2 g422_s_0(.a(n422),.q0(n422_0),.q1(n422_1));
  bfr _b_990(.a(_w_1445),.q(_w_1446));
  and_bi g248(.a(n247),.b(n240_1),.q(n248));
  spl2 g45_s_0(.a(n45),.q0(n45_0),.q1(n45_1));
  bfr _b_1721(.a(_w_2176),.q(_w_2177));
  spl3L g254_s_0(.a(n254),.q0(n254_0),.q1(n254_1),.q2(n254_2));
  spl2 g182_s_0(.a(n182),.q0(n182_0),.q1(n182_1));
  or_bb g167(.a(n156_1),.b(n158_1),.q(_w_2488));
  bfr _b_1045(.a(_w_1500),.q(_w_1501));
  spl2 g336_s_0(.a(n336),.q0(n336_0),.q1(n336_1));
  spl2 g337_s_0(.a(n337),.q0(n337_0),.q1(n337_1));
  spl2 g323_s_0(.a(n323),.q0(n323_0),.q1(n323_1));
  spl2 g351_s_0(.a(n351),.q0(n351_0),.q1(_w_2484));
  bfr _b_1338(.a(_w_1793),.q(b_1__5));
  spl2 g260_s_0(.a(n260),.q0(n260_0),.q1(n260_1));
  spl2 g406_s_0(.a(n406),.q0(n406_0),.q1(n406_1));
  bfr _b_1344(.a(_w_1799),.q(n57));
  and_bb g317(.a(a_4__9),.b(b_6__4),.q(n317));
  spl2 g411_s_0(.a(n411),.q0(n411_0),.q1(n411_1));
  bfr _b_1751(.a(_w_2206),.q(_w_2207));
  bfr _b_1170(.a(_w_1625),.q(_w_1626));
  or_bb g42(.a(n39_1),.b(n40_1),.q(_w_2483));
  spl2 g244_s_0(.a(n244),.q0(n244_0),.q1(n244_1));
  spl3L g256_s_0(.a(n256),.q0(n256_0),.q1(n256_1),.q2(n256_2));
  bfr _b_1500(.a(_w_1955),.q(_w_1956));
  spl2 g277_s_0(.a(n277),.q0(n277_0),.q1(n277_1));
  or_bb g453(.a(n244_1),.b(n256_2),.q(_w_2482));
  spl2 a_7__s_6(.a(a_7__11),.q0(_w_2480),.q1(a_7__13));
  bfr _b_905(.a(_w_1360),.q(n31_1));
  bfr _b_1433(.a(_w_1888),.q(_w_1889));
  spl2 g385_s_0(.a(n385),.q0(n385_0),.q1(n385_1));
  and_bi g446(.a(n445),.b(n439_1),.q(s_14_));
  bfr _b_1259(.a(_w_1714),.q(_w_1715));
  and_bi g444(.a(n443),.b(n384_1),.q(_w_2409));
  and_bb g240(.a(n224_0),.b(n239_0),.q(n240));
  spl2 g318_s_0(.a(n318),.q0(n318_0),.q1(_w_2491));
  or_bb g440(.a(n412),.b(n439_0),.q(s_15_));
  bfr _b_1327(.a(_w_1782),.q(_w_1783));
  bfr _b_1280(.a(_w_1735),.q(n396));
  or_bb g438(.a(n425_1),.b(n437_0),.q(n438));
  and_bb g302(.a(n300_0),.b(n301_0),.q(n302));
  spl2 a_1__s_4(.a(a_1__9),.q0(a_1__10),.q1(a_1__11));
  or_bb g430(.a(n358_1),.b(n361_1),.q(n430));
  and_bi g427(.a(n426),.b(n425_0),.q(n427));
  and_bb g26(.a(a_1__3),.b(b_5__2),.q(n26));
  spl2 g23_s_0(.a(n23),.q0(n23_0),.q1(n23_1));
  and_bb g425(.a(n416_0),.b(n424_0),.q(n425));
  bfr _b_1908(.a(_w_2363),.q(_w_2364));
  spl2 g366_s_0(.a(n366),.q0(n366_0),.q1(n366_1));
  bfr _b_1706(.a(_w_2161),.q(_w_2162));
  or_bb g424(.a(n419_1),.b(n423_0),.q(_w_2387));
  and_bi g429(.a(n428),.b(n423_1),.q(_w_2386));
  bfr _b_1665(.a(_w_2120),.q(_w_2121));
  bfr _b_1068(.a(_w_1523),.q(_w_1524));
  bfr _b_1733(.a(_w_2188),.q(_w_2189));
  or_bb g147(.a(n143_1),.b(n144_1),.q(_w_2408));
  or_bb g421(.a(n345_3),.b(n418_1),.q(_w_2385));
  or_bb g420(.a(n339_1),.b(n342_1),.q(_w_2378));
  and_bi g418(.a(n417),.b(n404_1),.q(n418));
  spl2 g18_s_0(.a(n18),.q0(n18_0),.q1(n18_1));
  spl2 a_7__s_2(.a(a_7__3),.q0(a_7__4),.q1(a_7__5));
  bfr _b_1636(.a(_w_2091),.q(_w_2092));
  bfr _b_1415(.a(_w_1870),.q(_w_1871));
  bfr _b_942(.a(_w_1397),.q(_w_1398));
  or_bb g415(.a(n406_1),.b(n408_1),.q(_w_2354));
  bfr _b_1724(.a(_w_2179),.q(_w_2180));
  and_bi g414(.a(n413),.b(n411_0),.q(_w_2327));
  or_bb g413(.a(n392_1),.b(n410_1),.q(_w_2326));
  and_bb g85(.a(n62_1),.b(n84_0),.q(n85));
  bfr _b_1928(.a(_w_2383),.q(_w_2384));
  and_bb g261(.a(n182_0),.b(n260_0),.q(n261));
  and_bb g411(.a(n392_0),.b(n410_0),.q(n411));
  and_bi g403(.a(n402),.b(n401_0),.q(n403));
  bfr _b_1240(.a(_w_1695),.q(_w_1696));
  and_bb g398(.a(b_6__11),.b(n325_1),.q(n398));
  and_bb g397(.a(a_5__12),.b(b_7__8),.q(_w_2325));
  bfr _b_1490(.a(_w_1945),.q(n250));
  and_bb g394(.a(a_6__13),.b(b_7__11),.q(n394));
  and_bi g366(.a(n365),.b(n356_1),.q(n366));
  or_bb g33(.a(n22_1),.b(n30_1),.q(_w_2324));
  and_bb g390(.a(a_7__12),.b(b_7__10),.q(n390));
  bfr _b_1973(.a(_w_2428),.q(_w_2429));
  and_bb g152(.a(a_0__0),.b(b_5__5),.q(n152));
  and_bb g387(.a(n375_0),.b(n385_0),.q(n387));
  bfr _b_1961(.a(_w_2416),.q(_w_2417));
  spl2 g198_s_0(.a(n198),.q0(n198_0),.q1(n198_1));
  bfr _b_1260(.a(_w_1715),.q(_w_1716));
  or_bb g406(.a(n398_1),.b(n401_1),.q(_w_2302));
  bfr _b_1596(.a(_w_2051),.q(_w_2052));
  or_bb g377(.a(n368_1),.b(n370_1),.q(_w_2301));
  or_bb g374(.a(n363_1),.b(n372_1),.q(_w_2288));
  bfr _b_914(.a(_w_1369),.q(_w_1370));
  and_bb g371(.a(n368_0),.b(n370_0),.q(n371));
  bfr _b_1613(.a(_w_2068),.q(_w_2069));
  and_bi g61(.a(n60),.b(n59_0),.q(n61));
  and_bb g242(.a(n220_0),.b(n241_0),.q(n242));
  bfr _b_957(.a(_w_1412),.q(n56_1));
  bfr _b_1754(.a(_w_2209),.q(_w_2210));
  and_bi g370(.a(n369),.b(n367_0),.q(n370));
  bfr _b_1033(.a(_w_1488),.q(_w_1489));
  bfr _b_1394(.a(_w_1849),.q(_w_1850));
  spl2 g434_s_0(.a(n434),.q0(n434_0),.q1(n434_1));
  or_bb g368(.a(n274_1),.b(n277_1),.q(_w_2276));
  bfr _b_915(.a(_w_1370),.q(_w_1371));
  or_bb g412(.a(n391_1),.b(n411_1),.q(_w_2246));
  and_bb g367(.a(n364_0),.b(n366_0),.q(n367));
  bfr _b_1860(.a(_w_2315),.q(_w_2316));
  spl2 g191_s_0(.a(n191),.q0(n191_0),.q1(n191_1));
  bfr _b_1342(.a(_w_1797),.q(n93_1));
  or_bb g365(.a(n353_1),.b(n355_1),.q(_w_2245));
  bfr _b_1880(.a(_w_2335),.q(_w_2336));
  or_bb g364(.a(n295_1),.b(n298_1),.q(n364));
  and_bb g272(.a(a_3__9),.b(b_6__3),.q(n272));
  or_bb g359(.a(n347_1),.b(n357_1),.q(_w_2244));
  spl2 a_6__s_6(.a(a_6__11),.q0(a_6__12),.q1(_w_2241));
  or_bb g357(.a(n351_1),.b(n356_0),.q(_w_2238));
  bfr _b_1552(.a(_w_2007),.q(n137));
  bfr _b_981(.a(_w_1436),.q(_w_1437));
  bfr _b_1601(.a(_w_2056),.q(_w_2057));
  and_bi g355(.a(n354),.b(n322_0),.q(n355));
  and_bi g121(.a(n120),.b(n117_0),.q(n121));
  or_bb g354(.a(n319_1),.b(n321_1),.q(_w_2237));
  and_bb g326(.a(a_7__6),.b(b_4__10),.q(n326));
  or_bb g283(.a(n281),.b(n282_0),.q(n283));
  bfr _b_1761(.a(_w_2216),.q(_w_2217));
  bfr _b_1698(.a(_w_2153),.q(_w_2154));
  or_bb g36(.a(n31_1),.b(n35_1),.q(_w_2228));
  and_bi g350(.a(n349),.b(n336_1),.q(_w_2227));
  spl2 b_1__s_2(.a(b_1__5),.q0(b_1__6),.q1(_w_2224));
  bfr _b_940(.a(_w_1395),.q(_w_1396));
  bfr _b_1835(.a(_w_2290),.q(_w_2291));
  bfr _b_1024(.a(_w_1479),.q(_w_1480));
  or_bb g443(.a(n381_1),.b(n383_1),.q(_w_2223));
  and_bi g246(.a(n245),.b(n241_1),.q(n246));
  bfr _b_1659(.a(_w_2114),.q(_w_2115));
  or_bb g314(.a(n19_2),.b(n250_1),.q(_w_2509));
  spl2 g345_s_0(.a(n345),.q0(n345_0),.q1(n345_1));
  and_bb g342(.a(n330_0),.b(n341_0),.q(n342));
  and_bb g255(.a(n248_0),.b(n254_0),.q(n255));
  spl2 b_7__s_4(.a(b_7__9),.q0(b_7__10),.q1(b_7__11));
  bfr _b_2008(.a(_w_2463),.q(_w_2464));
  bfr _b_1425(.a(_w_1880),.q(_w_1881));
  and_bb g339(.a(n337_0),.b(n338_0),.q(n339));
  and_bb g338(.a(a_5__11),.b(b_6__7),.q(_w_2221));
  and_bb g336(.a(n332_0),.b(n335_0),.q(n336));
  bfr _b_1935(.a(_w_2390),.q(_w_2391));
  and_bi g335(.a(n334),.b(n331_0),.q(n335));
  bfr _b_1269(.a(_w_1724),.q(_w_1725));
  bfr _b_1087(.a(_w_1542),.q(_w_1543));
  bfr _b_1501(.a(_w_1956),.q(_w_1957));
  or_bb g334(.a(n284_2),.b(n333),.q(n334));
  bfr _b_1182(.a(_w_1637),.q(_w_1638));
  bfr _b_929(.a(_w_1384),.q(_w_1385));
  and_bb g333(.a(a_7__8),.b(b_3__11),.q(n333));
  bfr _b_1040(.a(_w_1495),.q(_w_1496));
  bfr _b_2078(.a(_w_2533),.q(_w_2534));
  bfr _b_2063(.a(_w_2518),.q(_w_2514));
  and_bb g332(.a(a_5__9),.b(b_5__8),.q(n332));
  and_bb g330(.a(a_4__10),.b(b_7__6),.q(_w_2218));
  bfr _b_1965(.a(_w_2420),.q(_w_2421));
  bfr _b_1210(.a(_w_1665),.q(n48));
  bfr _b_898(.a(_w_1353),.q(_w_1354));
  bfr _b_1512(.a(_w_1967),.q(_w_1968));
  and_bi g442(.a(n441),.b(n255_1),.q(_w_2176));
  or_bb g328(.a(n326_1),.b(n327),.q(_w_2174));
  bfr _b_2003(.a(_w_2458),.q(_w_2459));
  spl2 g324_s_0(.a(n324),.q0(n324_0),.q1(_w_2165));
  and_bb g23(.a(a_2__2),.b(b_4__2),.q(n23));
  spl2 g215_s_1(.a(n215_1),.q0(n215_2),.q1(n215_3));
  and_bi g433(.a(n432),.b(n431_0),.q(_w_2149));
  and_bb g405(.a(n396_0),.b(n404_0),.q(n405));
  or_bb g402(.a(n397_1),.b(n400_1),.q(_w_2148));
  and_bi g360(.a(n359),.b(n358_0),.q(n360));
  spl2 g335_s_0(.a(n335),.q0(n335_0),.q1(n335_1));
  bfr _b_1025(.a(_w_1480),.q(_w_1481));
  bfr _b_863(.a(_w_1318),.q(_w_1319));
  bfr _b_2117(.a(_w_2572),.q(_w_2573));
  and_bb g327(.a(a_6__10),.b(b_5__11),.q(n327));
  bfr _b_1092(.a(_w_1547),.q(_w_1548));
  spl2 g403_s_0(.a(n403),.q0(n403_0),.q1(n403_1));
  bfr _b_1076(.a(_w_1531),.q(a_3__2));
  and_bb g391(.a(n389_2),.b(n390_0),.q(n391));
  spl2 g355_s_0(.a(n355),.q0(n355_0),.q1(n355_1));
  and_bb g37(.a(a_1__10),.b(b_7__2),.q(_w_2132));
  bfr _b_1370(.a(_w_1825),.q(_w_1826));
  bfr _b_1323(.a(_w_1778),.q(_w_1779));
  bfr _b_1226(.a(_w_1681),.q(_w_1682));
  spl2 g173_s_0(.a(n173),.q0(n173_0),.q1(n173_1));
  bfr _b_1400(.a(_w_1855),.q(_w_1856));
  bfr _b_891(.a(_w_1346),.q(_w_1347));
  spl2 g250_s_0(.a(n250),.q0(n250_0),.q1(n250_1));
  bfr _b_1939(.a(_w_2394),.q(_w_2395));
  spl2 b_7__s_2(.a(b_7__5),.q0(b_7__6),.q1(b_7__7));
  or_bb g395(.a(n393),.b(n394),.q(_w_2129));
  or_bb g96(.a(n83_1),.b(n92_1),.q(_w_2128));
  spl2 g398_s_0(.a(n398),.q0(n398_0),.q1(_w_2123));
  and_bb g312(.a(n268_1),.b(n310_1),.q(n312));
  or_bb g27(.a(n23_1),.b(n24_1),.q(_w_2102));
  bfr _b_1281(.a(_w_1736),.q(_w_1737));
  or_bb g311(.a(n268_0),.b(n310_0),.q(n311));
  or_bb g127(.a(n107_1),.b(n123_1),.q(_w_2101));
  spl2 g326_s_0(.a(n326),.q0(n326_0),.q1(_w_2096));
  or_bb g380(.a(n268_2),.b(n308_1),.q(n380));
  and_bi g310(.a(n309_0),.b(n308_0),.q(n310));
  bfr _b_1123(.a(_w_1578),.q(_w_1579));
  and_bi g196(.a(n195),.b(n193_0),.q(n196));
  and_bi g78(.a(n77),.b(n76_0),.q(n78));
  or_bb g309(.a(n269_1),.b(n307_1),.q(_w_2088));
  spl2 b_0__s_4(.a(b_0__9),.q0(b_0__10),.q1(b_0__11));
  and_bi g307(.a(n306),.b(n305_0),.q(n307));
  bfr _b_1856(.a(_w_2311),.q(n193_1));
  bfr _b_1395(.a(_w_1850),.q(_w_1851));
  bfr _b_1151(.a(_w_1606),.q(_w_1607));
  bfr _b_1139(.a(_w_1594),.q(s_8_));
  or_bb g219(.a(n186_1),.b(n214_1),.q(_w_2087));
  spl2 g149_s_0(.a(n149),.q0(n149_0),.q1(n149_1));
  bfr _b_1063(.a(_w_1518),.q(_w_1519));
  bfr _b_1642(.a(_w_2097),.q(_w_2098));
  and_bb g305(.a(n270_0),.b(n304_0),.q(n305));
  spl2 g435_s_0(.a(n435),.q0(n435_0),.q1(n435_1));
  and_bi g383(.a(n382),.b(n379_0),.q(n383));
  spl2 g168_s_0(.a(n168),.q0(n168_0),.q1(_w_2078));
  spl2 g146_s_0(.a(n146),.q0(n146_0),.q1(n146_1));
  and_bi g300(.a(n299),.b(n298_0),.q(n300));
  or_bb g92(.a(n85_1),.b(n91_0),.q(n92));
  and_bb g379(.a(n376_0),.b(n378_0),.q(n379));
  or_bb g299(.a(n279_1),.b(n297_1),.q(_w_2076));
  and_bi g315(.a(n314),.b(n251_1),.q(_w_2037));
  and_bi g297(.a(n296),.b(n295_0),.q(n297));
  spl2 g272_s_0(.a(n272),.q0(n272_0),.q1(n272_1));
  or_bb g288(.a(n280_1),.b(n286_1),.q(_w_2036));
  bfr _b_2025(.a(_w_2480),.q(_w_2481));
  bfr _b_1083(.a(_w_1538),.q(_w_1539));
  bfr _b_1870(.a(_w_2325),.q(n397));
  bfr _b_1484(.a(_w_1939),.q(_w_1940));
  or_bb g294(.a(n76_1),.b(n79_1),.q(n294));
  bfr _b_1166(.a(_w_1621),.q(_w_1622));
  spl2 g389_s_0(.a(n389),.q0(n389_0),.q1(_w_2034));
  or_bb g292(.a(n289_1),.b(n290_1),.q(_w_2033));
  and_bi g289(.a(n288),.b(n287_0),.q(n289));
  bfr _b_874(.a(_w_1329),.q(_w_1330));
  bfr _b_1909(.a(_w_2364),.q(_w_2365));
  and_bb g358(.a(n347_0),.b(n357_0),.q(n358));
  bfr _b_2118(.a(_w_2573),.q(_w_2574));
  and_bb g287(.a(n280_0),.b(n286_0),.q(n287));
  or_bb g269(.a(n131_1),.b(n134_1),.q(n269));
  bfr _b_1955(.a(_w_2410),.q(_w_2411));
  bfr _b_1527(.a(_w_1982),.q(n168));
  bfr _b_1518(.a(_w_1973),.q(_w_1974));
  and_bb g282(.a(a_6__6),.b(b_3__6),.q(n282));
  bfr _b_1822(.a(_w_2277),.q(_w_2278));
  bfr _b_1186(.a(_w_1641),.q(a_7__9));
  spl2 g364_s_0(.a(n364),.q0(n364_0),.q1(n364_1));
  and_bb g280(.a(a_4__7),.b(b_5__6),.q(n280));
  bfr _b_1134(.a(_w_1589),.q(_w_1590));
  spl2 g317_s_0(.a(n317),.q0(n317_0),.q1(n317_1));
  bfr _b_1682(.a(_w_2137),.q(_w_2138));
  and_bb g308(.a(n269_0),.b(n307_0),.q(_w_2013));
  and_bb g274(.a(n272_0),.b(n273_0),.q(n274));
  and_bi g140(.a(n139),.b(n122_1),.q(n140));
  and_bi g138(.a(n137),.b(n129_1),.q(n138));
  and_bb g257(.a(n244_0),.b(n256_0),.q(n257));
  spl4L b_2__s_2(.a(b_2__1),.q0(b_2__5),.q1(b_2__6),.q2(b_2__7),.q3(_w_2012));
  and_bi g329(.a(n328),.b(n325_0),.q(_w_2211));
  and_bb g88(.a(a_6__2),.b(b_0__6),.q(n88));
  spl2 g54_s_0(.a(n54),.q0(n54_0),.q1(n54_1));
  spl2 g401_s_0(.a(n401),.q0(n401_0),.q1(n401_1));
  or_bb g137(.a(n126_1),.b(n128_1),.q(_w_2007));
  bfr _b_1145(.a(_w_1600),.q(_w_1601));
  spl2 g269_s_0(.a(n269),.q0(n269_0),.q1(n269_1));
  and_bb g151(.a(n142_0),.b(n150_0),.q(n151));
  bfr _b_1445(.a(_w_1900),.q(a_1__7));
  or_bb g436(.a(n431_1),.b(n435_0),.q(n436));
  bfr _b_1653(.a(_w_2108),.q(_w_2109));
  and_bi g148(.a(n147),.b(n145_0),.q(n148));
  and_bi g90(.a(n89),.b(n85_0),.q(n90));
  bfr _b_1873(.a(_w_2328),.q(_w_2329));
  bfr _b_1811(.a(_w_2266),.q(_w_2267));
  and_bi g95(.a(n94),.b(n45_1),.q(n95));
  bfr _b_1581(.a(_w_2036),.q(n288));
  bfr _b_859(.a(_w_1314),.q(n181_1));
  or_bb g132(.a(n105_1),.b(n130_1),.q(_w_1999));
  bfr _b_1380(.a(_w_1835),.q(_w_1836));
  spl2 a_6__s_5(.a(a_6__9),.q0(a_6__10),.q1(_w_1997));
  or_bb g130(.a(n124_1),.b(n129_0),.q(n130));
  bfr _b_967(.a(_w_1422),.q(_w_1423));
  and_bb g129(.a(n126_0),.b(n128_0),.q(n129));
  spl2 g287_s_0(.a(n287),.q0(n287_0),.q1(n287_1));
  and_bb g53(.a(a_3__7),.b(b_5__4),.q(n53));
  bfr _b_1117(.a(_w_1572),.q(_w_1573));
  or_bb g187(.a(n160_1),.b(n162_1),.q(_w_1996));
  bfr _b_1888(.a(_w_2343),.q(_w_2344));
  and_bi g388(.a(n386),.b(n387_0),.q(_w_1984));
  or_bb g296(.a(n293_1),.b(n294_1),.q(_w_1983));
  and_bb g168(.a(n166_0),.b(n167_0),.q(_w_1981));
  bfr _b_1617(.a(_w_2072),.q(_w_2073));
  and_bi g128(.a(n127),.b(n124_0),.q(n128));
  and_bb g193(.a(n191_0),.b(n192_0),.q(n193));
  bfr _b_926(.a(_w_1381),.q(_w_1382));
  bfr _b_1362(.a(_w_1817),.q(n325_2));
  bfr _b_1215(.a(_w_1670),.q(n346));
  and_bi g375(.a(n374),.b(n373_0),.q(n375));
  and_bb g194(.a(a_1__1),.b(b_2__7),.q(n194));
  bfr _b_2081(.a(b_2_),.q(_w_2537));
  or_bb g123(.a(n117_1),.b(n122_0),.q(n123));
  bfr _b_1143(.a(_w_1598),.q(_w_1599));
  and_bb g319(.a(a_3__10),.b(b_7__4),.q(_w_2127));
  spl2 g439_s_0(.a(n439),.q0(n439_0),.q1(n439_1));
  spl3L a_1__s_0(.a(_w_2514),.q0(a_1__0),.q1(a_1__1),.q2(_w_1977));
  bfr _b_1030(.a(_w_1485),.q(_w_1486));
  and_bb g325(.a(n284_3),.b(n324_0),.q(n325));
  and_bi g119(.a(n118),.b(n29_1),.q(n119));
  bfr _b_844(.a(_w_1299),.q(n216_1));
  bfr _b_1877(.a(_w_2332),.q(_w_2333));
  or_bb g445(.a(n414_1),.b(n438_1),.q(_w_1976));
  or_bb g118(.a(n26_1),.b(n28_1),.q(_w_1975));
  spl2 g97_s_0(.a(n97),.q0(n97_0),.q1(n97_1));
  bfr _b_842(.a(_w_1297),.q(_w_1298));
  bfr _b_1379(.a(_w_1834),.q(_w_1835));
  spl2 g397_s_0(.a(n397),.q0(n397_0),.q1(n397_1));
  bfr _b_1056(.a(_w_1511),.q(_w_1512));
  and_bi g234(.a(n233),.b(n197_1),.q(_w_1967));
  bfr _b_1715(.a(_w_2170),.q(_w_2171));
  and_bb g111(.a(n110_0),.b(n84_1),.q(n111));
  bfr _b_1673(.a(_w_2128),.q(n96));
  bfr _b_1420(.a(_w_1875),.q(_w_1876));
  spl3L a_1__s_1(.a(a_1__2),.q0(a_1__3),.q1(a_1__4),.q2(a_1__5));
  spl2 g282_s_0(.a(n282),.q0(n282_0),.q1(_w_1964));
  and_bi g105(.a(n104),.b(n103_0),.q(n105));
  or_bb g106(.a(n95_1),.b(n97_1),.q(_w_1966));
  and_bb g115(.a(n112_0),.b(n114_0),.q(n115));
  or_bb g434(.a(n373_1),.b(n387_1),.q(n434));
  bfr _b_1726(.a(_w_2181),.q(_w_2182));
  bfr _b_983(.a(_w_1438),.q(_w_1439));
  bfr _b_1760(.a(_w_2215),.q(_w_2216));
  bfr _b_1589(.a(_w_2044),.q(_w_2045));
  and_bi g160(.a(n159),.b(n158_0),.q(n160));
  and_bi g230(.a(n229),.b(n227_0),.q(n230));
  or_bb g369(.a(n364_1),.b(n366_1),.q(_w_1963));
  and_bb g32(.a(a_0__7),.b(b_7__0),.q(_w_1961));
  spl2 g62_s_2(.a(n62_4),.q0(n62_5),.q1(n62_6));
  bfr _b_1612(.a(_w_2067),.q(_w_2068));
  spl2 g316_s_0(.a(n316),.q0(n316_0),.q1(n316_1));
  bfr _b_1106(.a(_w_1561),.q(_w_1562));
  and_bb g254(.a(n251_0),.b(n253_0),.q(n254));
  and_bi g452(.a(n451),.b(n435_1),.q(_w_1953));
  bfr _b_1531(.a(_w_1986),.q(_w_1987));
  or_bb g125(.a(n32_1),.b(n34_1),.q(_w_1980));
  spl2 g297_s_0(.a(n297),.q0(n297_0),.q1(n297_1));
  spl2 g199_s_0(.a(n199),.q0(n199_0),.q1(_w_1949));
  spl2 a_7__s_1(.a(a_7__1),.q0(a_7__2),.q1(_w_1948));
  bfr _b_1042(.a(_w_1497),.q(_w_1498));
  bfr _b_1043(.a(_w_1498),.q(_w_1499));
  or_bb g441(.a(n248_1),.b(n254_2),.q(_w_1947));
  bfr _b_2015(.a(_w_2470),.q(_w_2471));
  bfr _b_1817(.a(_w_2272),.q(_w_2273));
  spl2 g298_s_0(.a(n298),.q0(n298_0),.q1(n298_1));
  or_bb g80(.a(n61_1),.b(n78_1),.q(_w_1946));
  and_bi g250(.a(n249),.b(n231_1),.q(_w_1938));
  or_bb g176(.a(n138_1),.b(n174_1),.q(_w_1937));
  bfr _b_1564(.a(_w_2019),.q(_w_2020));
  bfr _b_1414(.a(_w_1869),.q(_w_1870));
  and_bb g73(.a(a_7__2),.b(b_2__3),.q(n73));
  spl4L a_2__s_1(.a(a_2__1),.q0(a_2__2),.q1(a_2__3),.q2(a_2__4),.q3(_w_1934));
  spl3L g251_s_0(.a(n251),.q0(n251_0),.q1(n251_1),.q2(n251_2));
  and_bb g91(.a(n86_0),.b(n90_0),.q(n91));
  spl2 a_0__s_4(.a(a_0__9),.q0(a_0__10),.q1(a_0__11));
  and_bb g134(.a(n133_0),.b(n36_0),.q(n134));
  bfr _b_1845(.a(_w_2300),.q(n374));
  or_bb g89(.a(n87),.b(n88),.q(n89));
  bfr _b_1655(.a(_w_2110),.q(_w_2111));
  and_bi g83(.a(n82),.b(n68_1),.q(n83));
  spl2 g425_s_0(.a(n425),.q0(n425_0),.q1(_w_1929));
  and_bb g404(.a(n324_2),.b(n403_0),.q(n404));
  bfr _b_1784(.a(_w_2239),.q(_w_2240));
  and_bb g251(.a(n19_1),.b(n250_0),.q(n251));
  and_bb g112(.a(a_3__5),.b(b_2__5),.q(n112));
  or_bb g270(.a(n47_1),.b(n50_1),.q(_w_1918));
  bfr _b_1697(.a(_w_2152),.q(_w_2153));
  spl2 g373_s_0(.a(n373),.q0(n373_0),.q1(_w_1914));
  bfr _b_1165(.a(_w_1620),.q(_w_1621));
  and_bi g218(.a(n217),.b(n216_0),.q(n218));
  and_bb g318(.a(n316_0),.b(n317_0),.q(n318));
  bfr _b_880(.a(_w_1335),.q(_w_1336));
  bfr _b_1778(.a(_w_2233),.q(_w_2234));
  bfr _b_1130(.a(_w_1585),.q(_w_1586));
  bfr _b_890(.a(_w_1345),.q(_w_1346));
  bfr _b_2054(.a(_w_2509),.q(n314));
  and_bb g144(.a(a_3__0),.b(b_1__3),.q(n144));
  and_bi g126(.a(n125),.b(n35_0),.q(n126));
  bfr _b_1746(.a(_w_2201),.q(_w_2202));
  and_bi g448(.a(n447),.b(n259_1),.q(_w_2436));
  spl2 b_0__s_0(.a(b_0_),.q0(b_0__0),.q1(b_0__1));
  and_bb g45(.a(n43_0),.b(n44_0),.q(n45));
  bfr _b_1436(.a(_w_1891),.q(a_5__8));
  or_bb g385(.a(n379_1),.b(n384_0),.q(n385));
  bfr _b_875(.a(_w_1330),.q(n100_1));
  spl3L a_2__s_2(.a(a_2__5),.q0(a_2__6),.q1(a_2__7),.q2(_w_1907));
  spl2 g166_s_0(.a(n166),.q0(n166_0),.q1(n166_1));
  and_bb g437(.a(n427_0),.b(n436_0),.q(n437));
  bfr _b_951(.a(_w_1406),.q(_w_1407));
  or_bb g77(.a(n69_1),.b(n75_1),.q(_w_1906));
  spl2 g22_s_0(.a(n22),.q0(n22_0),.q1(n22_1));
  bfr _b_1149(.a(_w_1604),.q(_w_1605));
  bfr _b_1086(.a(_w_1541),.q(_w_1542));
  and_bb g25(.a(n23_0),.b(n24_0),.q(n25));
  bfr _b_2023(.a(_w_2478),.q(s_13_));
  and_bb g322(.a(n319_0),.b(n321_0),.q(n322));
  spl3L g55_s_0(.a(n55),.q0(n55_0),.q1(n55_1),.q2(n55_2));
  and_bb g39(.a(a_3__4),.b(b_4__3),.q(n39));
  spl2 g112_s_0(.a(n112),.q0(n112_0),.q1(n112_1));
  and_bi g321(.a(n320),.b(n318_0),.q(n321));
  or_bb g161(.a(n142_1),.b(n150_1),.q(_w_1904));
  and_bb g38(.a(a_2__9),.b(b_6__2),.q(n38));
  bfr _b_1195(.a(_w_1650),.q(n223));
  or_bb g316(.a(n285_1),.b(n287_1),.q(n316));
  or_bb g372(.a(n367_1),.b(n371_0),.q(_w_2285));
  bfr _b_922(.a(_w_1377),.q(_w_1378));
  and_bb g84(.a(a_5__0),.b(b_0__2),.q(n84));
  and_bb g100(.a(n81_0),.b(n99_0),.q(n100));
  spl2 a_1__s_2(.a(a_1__5),.q0(a_1__6),.q1(_w_1900));
  and_bb g76(.a(n69_0),.b(n75_0),.q(n76));
  or_bb g349(.a(n332_1),.b(n335_1),.q(_w_1899));
  bfr _b_1489(.a(_w_1944),.q(_w_1945));
  spl2 g310_s_0(.a(n310),.q0(n310_0),.q1(n310_1));
  and_bb g373(.a(n363_0),.b(n372_0),.q(_w_2463));
  or_bb g183(.a(n168_3),.b(n177_1),.q(_w_1898));
  bfr _b_2040(.a(_w_2495),.q(n135));
  spl2 g90_s_0(.a(n90),.q0(n90_0),.q1(n90_1));
  bfr _b_1809(.a(_w_2264),.q(_w_2265));
  bfr _b_1663(.a(_w_2118),.q(_w_2119));
  spl2 g430_s_0(.a(n430),.q0(n430_0),.q1(n430_1));
  bfr _b_1600(.a(_w_2055),.q(_w_2056));
  and_bb g31(.a(n22_0),.b(n30_0),.q(n31));
  spl2 g339_s_0(.a(n339),.q0(n339_0),.q1(_w_1894));
  spl2 g192_s_0(.a(n192),.q0(n192_0),.q1(n192_1));
  bfr _b_1529(.a(_w_1984),.q(_w_1985));
  spl2 g92_s_0(.a(n92),.q0(n92_0),.q1(n92_1));
  or_bb g340(.a(n337_1),.b(n338_1),.q(_w_1893));
  bfr _b_964(.a(_w_1419),.q(_w_1420));
  and_bb g143(.a(a_4__1),.b(b_0__3),.q(n143));
  and_bb g235(.a(n232_0),.b(n234_0),.q(n235));
  and_bb g149(.a(n146_0),.b(n148_0),.q(n149));
  spl2 a_6__s_2(.a(a_6__3),.q0(a_6__4),.q1(a_6__5));
  bfr _b_1959(.a(_w_2414),.q(_w_2415));
  bfr _b_1181(.a(_w_1636),.q(_w_1637));
  bfr _b_1103(.a(_w_1558),.q(_w_1559));
  bfr _b_1310(.a(_w_1765),.q(_w_1766));
  and_bb g93(.a(n83_0),.b(n92_0),.q(n93));
  and_bb g271(.a(a_2__10),.b(b_7__3),.q(_w_2077));
  spl2 g143_s_0(.a(n143),.q0(n143_0),.q1(n143_1));
  spl2 g381_s_0(.a(n381),.q0(n381_0),.q1(n381_1));
  and_bi g276(.a(n275),.b(n274_0),.q(n276));
  or_bb g104(.a(n102_1),.b(n52_1),.q(_w_1892));
  and_bb g41(.a(n39_0),.b(n40_0),.q(n41));
  bfr _b_1936(.a(_w_2391),.q(_w_2392));
  spl2 a_5__s_3(.a(a_5__6),.q0(a_5__7),.q1(_w_1888));
  spl2 g302_s_0(.a(n302),.q0(n302_0),.q1(_w_2133));
  spl2 g342_s_0(.a(n342),.q0(n342_0),.q1(n342_1));
  or_bb g171(.a(n140_1),.b(n164_1),.q(_w_1887));
  bfr _b_1592(.a(_w_2047),.q(_w_2048));
  or_bb g164(.a(n151_1),.b(n163_0),.q(n164));
  and_bb g79(.a(n61_0),.b(n78_0),.q(n79));
  or_bb g113(.a(n110_1),.b(n84_2),.q(_w_1886));
  and_bb g201(.a(a_0__3),.b(b_4__11),.q(n201));
  bfr _b_1498(.a(_w_1953),.q(_w_1954));
  or_bb g249(.a(n228_1),.b(n230_1),.q(_w_1885));
  bfr _b_1711(.a(_w_2166),.q(_w_2167));
  spl2 g257_s_0(.a(n257),.q0(n257_0),.q1(n257_1));
  bfr _b_1085(.a(_w_1540),.q(_w_1541));
  bfr _b_1352(.a(_w_1807),.q(_w_1808));
  and_bb g455(.a(a_0__11),.b(b_0__11),.q(_w_1832));
  bfr _b_2114(.a(_w_2569),.q(_w_2570));
  or_bb g337(.a(n331_1),.b(n336_0),.q(n337));
  and_bb g56(.a(n54_0),.b(n55_0),.q(n56));
  spl3L a_0__s_3(.a(a_0__6),.q0(a_0__7),.q1(a_0__8),.q2(a_0__9));
  spl2 g437_s_0(.a(n437),.q0(n437_0),.q1(n437_1));
  or_bb g407(.a(n396_1),.b(n404_2),.q(_w_1831));
  or_bb g108(.a(n86_1),.b(n90_1),.q(_w_1830));
  spl2 g301_s_0(.a(n301),.q0(n301_0),.q1(n301_1));
  and_bi g408(.a(n407),.b(n405_0),.q(n408));
  and_bi g222(.a(n221),.b(n213_1),.q(_w_1828));
  bfr _b_1622(.a(_w_2077),.q(n271));
  and_bi g220(.a(n219),.b(n215_0),.q(n220));
  and_bi g43(.a(n42),.b(n41_0),.q(n43));
  and_bi g182(.a(n180),.b(n181_0),.q(n182));
  bfr _b_1744(.a(_w_2199),.q(_w_2200));
  and_bb g63(.a(a_7__0),.b(b_0__0),.q(_w_1823));
  or_bb g150(.a(n145_1),.b(n149_0),.q(n150));
  spl2 g158_s_0(.a(n158),.q0(n158_0),.q1(n158_1));
  and_bb g158(.a(n152_0),.b(n157_0),.q(n158));
  spl2 g284_s_0(.a(n284),.q0(n284_0),.q1(_w_1820));
  spl2 g121_s_0(.a(n121),.q0(n121_0),.q1(n121_1));
  and_bb g431(.a(n429_0),.b(n430_0),.q(n431));
  and_bi g190(.a(n189),.b(n149_1),.q(n190));
  bfr _b_1386(.a(_w_1841),.q(_w_1842));
  bfr _b_1244(.a(_w_1699),.q(_w_1700));
  bfr _b_873(.a(_w_1328),.q(_w_1329));
  bfr _b_1152(.a(_w_1607),.q(_w_1608));
  and_bb g22(.a(a_1__8),.b(b_6__0),.q(_w_1819));
  bfr _b_1247(.a(_w_1702),.q(_w_1703));
  and_bb g356(.a(n353_0),.b(n355_0),.q(n356));
  and_bi g378(.a(n377),.b(n371_1),.q(_w_2425));
  spl3L g84_s_0(.a(n84),.q0(n84_0),.q1(n84_1),.q2(n84_2));
  bfr _b_944(.a(_w_1399),.q(_w_1400));
  bfr _b_970(.a(_w_1425),.q(_w_1426));
  or_bb g66(.a(n62_3),.b(n63_1),.q(n66));
  bfr _b_1457(.a(_w_1912),.q(_w_1913));
  and_bb g122(.a(n119_0),.b(n121_0),.q(n122));
  and_bb g86(.a(a_4__5),.b(b_2__4),.q(n86));
  bfr _b_1902(.a(_w_2357),.q(_w_2358));
  and_bb g50(.a(n37_0),.b(n49_0),.q(n50));
  spl2 g420_s_0(.a(n420),.q0(n420_0),.q1(n420_1));
  or_bb g236(.a(n232_1),.b(n234_1),.q(_w_2026));
  spl2 g324_s_1(.a(n324_1),.q0(n324_2),.q1(n324_3));
  or_bb g46(.a(n41_1),.b(n45_0),.q(n46));
  and_bb g110(.a(a_4__0),.b(b_1__2),.q(n110));
  bfr _b_1325(.a(_w_1780),.q(s_1_));
  spl2 g291_s_0(.a(n291),.q0(n291_0),.q1(n291_1));
  and_bb g47(.a(n38_0),.b(n46_0),.q(n47));
  bfr _b_1557(.a(_w_2012),.q(b_2__8));
  spl2 g308_s_0(.a(n308),.q0(n308_0),.q1(_w_1815));
  spl2 g389_s_1(.a(n389_1),.q0(n389_2),.q1(n389_3));
  bfr _b_2079(.a(_w_2534),.q(_w_2520));
  spl3L g19_s_0(.a(n19),.q0(n19_0),.q1(n19_1),.q2(n19_2));
  or_bb g376(.a(n302_1),.b(n305_1),.q(_w_1804));
  bfr _b_1838(.a(_w_2293),.q(_w_2294));
  bfr _b_1266(.a(_w_1721),.q(_w_1722));
  bfr _b_1172(.a(_w_1627),.q(_w_1628));
  and_bi g49(.a(n48),.b(n47_0),.q(n49));
  and_bb g345(.a(n329_0),.b(n344_0),.q(n345));
  spl2 g414_s_0(.a(n414),.q0(n414_0),.q1(n414_1));
  bfr _b_1765(.a(_w_2220),.q(n330));
  spl2 g405_s_0(.a(n405),.q0(n405_0),.q1(_w_1800));
  or_bb g57(.a(n54_1),.b(n55_2),.q(_w_1799));
  and_bi g162(.a(n161),.b(n151_0),.q(n162));
  spl2 g383_s_0(.a(n383),.q0(n383_0),.q1(n383_1));
  and_bi g142(.a(n141),.b(n115_1),.q(n142));
  spl2 g28_s_0(.a(n28),.q0(n28_0),.q1(n28_1));
  bfr _b_1214(.a(_w_1669),.q(n264));
  or_bb g432(.a(n429_1),.b(n430_1),.q(_w_1798));
  bfr _b_928(.a(_w_1383),.q(n165_1));
  and_bb g178(.a(n168_2),.b(n177_0),.q(n178));
  spl2 g93_s_0(.a(n93),.q0(n93_0),.q1(_w_1794));
  bfr _b_2033(.a(_w_2488),.q(_w_2489));
  bfr _b_1218(.a(_w_1673),.q(n101));
  and_bi g290(.a(n73_1),.b(n62_6),.q(_w_2027));
  and_bb g285(.a(n284_0),.b(n55_1),.q(n285));
  bfr _b_1662(.a(_w_2117),.q(_w_2118));
  or_bb g399(.a(n325_2),.b(n389_0),.q(n399));
  bfr _b_1253(.a(_w_1708),.q(_w_1709));
  and_bb g381(.a(n309_1),.b(n380),.q(n381));
  bfr _b_999(.a(_w_1454),.q(n391_1));
  and_bb g165(.a(n140_0),.b(n164_0),.q(n165));
  spl2 g356_s_0(.a(n356),.q0(n356_0),.q1(n356_1));
  bfr _b_1064(.a(_w_1519),.q(_w_1520));
  bfr _b_1082(.a(_w_1537),.q(_w_1538));
  spl2 g433_s_0(.a(n433),.q0(n433_0),.q1(n433_1));
  and_bi g75(.a(n72),.b(n74_0),.q(n75));
  and_bi g136(.a(n135),.b(n134_0),.q(_w_1788));
  and_bb g59(.a(n53_0),.b(n58_0),.q(n59));
  or_bb g141(.a(n112_1),.b(n114_1),.q(_w_1787));
  spl2 g122_s_0(.a(n122),.q0(n122_0),.q1(n122_1));
  or_bb g245(.a(n222_1),.b(n240_2),.q(_w_1786));
  bfr _b_1729(.a(_w_2184),.q(_w_2185));
  and_bb g145(.a(n143_0),.b(n144_0),.q(n145));
  spl2 g144_s_0(.a(n144),.q0(n144_0),.q1(n144_1));
  and_bb g62(.a(a_6__0),.b(b_1__0),.q(_w_1785));
  bfr _b_1695(.a(_w_2150),.q(_w_2151));
  bfr _b_1077(.a(_w_1532),.q(_w_1533));
  and_bb g389(.a(a_6__12),.b(b_6__9),.q(n389));
  bfr _b_1797(.a(_w_2252),.q(_w_2253));
  bfr _b_1643(.a(_w_2098),.q(_w_2099));
  bfr _b_1416(.a(_w_1871),.q(_w_1872));
  spl2 g210_s_0(.a(n210),.q0(n210_0),.q1(_w_1781));
  and_bb g64(.a(n62_0),.b(n63_0),.q(n64));
  bfr _b_1785(.a(_w_2240),.q(n357));
  bfr _b_1473(.a(_w_1928),.q(a_0__6));
  spl2 a_0__s_1(.a(a_0__2),.q0(a_0__3),.q1(a_0__4));
  and_bi g21(.a(n20),.b(n19_0),.q(_w_1740));
  bfr _b_1432(.a(_w_1887),.q(n171));
  and_bb g393(.a(a_7__13),.b(b_6__12),.q(_w_1732));
  bfr _b_1999(.a(_w_2454),.q(_w_2455));
  spl2 g105_s_0(.a(n105),.q0(n105_0),.q1(n105_1));
  and_bb g439(.a(n414_0),.b(n438_0),.q(n439));
  or_bb g99(.a(n93_1),.b(n98_0),.q(n99));
  spl2 a_6__s_1(.a(a_6__1),.q0(a_6__2),.q1(_w_1731));
  bfr _b_1727(.a(_w_2182),.q(_w_2183));
  spl2 g79_s_0(.a(n79),.q0(n79_0),.q1(n79_1));
  bfr _b_1052(.a(_w_1507),.q(_w_1508));
  or_bb g303(.a(n300_1),.b(n301_1),.q(_w_1818));
  spl2 g358_s_0(.a(n358),.q0(n358_0),.q1(_w_1727));
  and_bb g213(.a(n204_2),.b(n212_0),.q(n213));
  spl2 g293_s_0(.a(n293),.q0(n293_0),.q1(n293_1));
  and_bb g103(.a(n102_0),.b(n52_0),.q(n103));
  or_bb g72(.a(n70),.b(n71),.q(n72));
  bfr _b_1743(.a(_w_2198),.q(_w_2199));
  or_bb g275(.a(n272_1),.b(n273_1),.q(_w_1726));
  bfr _b_1299(.a(_w_1754),.q(_w_1755));
  bfr _b_1262(.a(_w_1717),.q(_w_1718));
  spl2 g153_s_1(.a(n153_1),.q0(n153_2),.q1(_w_1723));
  bfr _b_1543(.a(_w_1998),.q(a_6__11));
  and_bb g70(.a(a_7__4),.b(b_1__8),.q(n70));
  and_bb g146(.a(a_2__3),.b(b_2__6),.q(n146));
  and_bi g207(.a(n206),.b(n199_0),.q(n207));
  and_bi g265(.a(n264),.b(n254_1),.q(_w_1686));
  bfr _b_1201(.a(_w_1656),.q(n159));
  spl2 g348_s_0(.a(n348),.q0(n348_0),.q1(n348_1));
  bfr _b_836(.a(_w_1291),.q(n235_1));
  bfr _b_867(.a(_w_1322),.q(_w_1323));
  bfr _b_1023(.a(_w_1478),.q(_w_1479));
  bfr _b_1932(.a(_w_2387),.q(_w_2388));
  and_bb g154(.a(a_2__4),.b(b_3__4),.q(n154));
  and_bi g353(.a(n352),.b(n351_0),.q(n353));
  spl2 g232_s_0(.a(n232),.q0(n232_0),.q1(n232_1));
  bfr _b_1028(.a(_w_1483),.q(_w_1484));
  and_bb g200(.a(a_1__6),.b(b_3__10),.q(n200));
  or_bb g428(.a(n420_1),.b(n422_1),.q(_w_1685));
  bfr _b_1769(.a(_w_2224),.q(_w_2225));
  spl2 g126_s_0(.a(n126),.q0(n126_0),.q1(n126_1));
  and_bb g423(.a(n420_0),.b(n422_0),.q(n423));
  bfr _b_1606(.a(_w_2061),.q(_w_2062));
  bfr _b_1447(.a(_w_1902),.q(_w_1903));
  bfr _b_1073(.a(_w_1528),.q(n85_1));
  or_bb g155(.a(n153_2),.b(n154_1),.q(n155));
  spl3L g62_s_0(.a(n62),.q0(n62_0),.q1(n62_1),.q2(n62_2));
  and_bb g65(.a(a_5__5),.b(b_2__2),.q(n65));
  and_bb g163(.a(n160_0),.b(n162_0),.q(n163));
  bfr _b_1426(.a(_w_1881),.q(_w_1882));
  spl2 g387_s_0(.a(n387),.q0(n387_0),.q1(n387_1));
  or_bb g174(.a(n165_1),.b(n173_0),.q(n174));
  spl2 g53_s_0(.a(n53),.q0(n53_0),.q1(n53_1));
  bfr _b_1273(.a(_w_1728),.q(_w_1729));
  bfr _b_861(.a(_w_1316),.q(n62_4));
  spl2 g258_s_0(.a(n258),.q0(n258_0),.q1(n258_1));
  or_bb g209(.a(n199_1),.b(n208_0),.q(n209));
  bfr _b_1275(.a(_w_1730),.q(n358_1));
  spl2 g116_s_0(.a(n116),.q0(n116_0),.q1(n116_1));
  spl2 g438_s_0(.a(n438),.q0(n438_0),.q1(n438_1));
  bfr _b_2077(.a(_w_2532),.q(_w_2533));
  and_bb g435(.a(n433_0),.b(n434_0),.q(n435));
  or_bb g306(.a(n270_1),.b(n304_1),.q(_w_1684));
  bfr _b_1647(.a(_w_2102),.q(n27));
  bfr _b_1439(.a(_w_1894),.q(_w_1895));
  bfr _b_1363(.a(_w_1818),.q(n303));
  bfr _b_1288(.a(_w_1743),.q(_w_1744));
  bfr _b_1091(.a(_w_1546),.q(_w_1547));
  and_bi g102(.a(n101),.b(n100_0),.q(n102));
  spl2 a_4__s_3(.a(a_4__8),.q0(a_4__9),.q1(_w_1680));
  and_bi g114(.a(n113),.b(n111_0),.q(n114));
  spl2 g341_s_0(.a(n341),.q0(n341_0),.q1(n341_1));
  or_bb g169(.a(n166_1),.b(n167_1),.q(_w_1677));
  or_bb g198(.a(n193_1),.b(n197_0),.q(n198));
  and_bb g175(.a(n138_0),.b(n174_0),.q(n175));
  spl3L a_4__s_0(.a(_w_2535),.q0(a_4__0),.q1(a_4__1),.q2(_w_1736));
  and_bi g170(.a(n169),.b(n168_0),.q(n170));
  spl2 g329_s_0(.a(n329),.q0(n329_0),.q1(n329_1));
  spl2 g138_s_0(.a(n138),.q0(n138_0),.q1(n138_1));
  bfr _b_1000(.a(_w_1455),.q(_w_1456));
  or_bb g30(.a(n25_1),.b(n29_0),.q(n30));
  spl2 g416_s_0(.a(n416),.q0(n416_0),.q1(n416_1));
  spl2 g322_s_0(.a(n322),.q0(n322_0),.q1(n322_1));
  bfr _b_894(.a(_w_1349),.q(_w_1350));
  bfr _b_1980(.a(_w_2435),.q(n378));
  bfr _b_1340(.a(_w_1795),.q(_w_1796));
  and_bb g173(.a(n170_0),.b(n172_0),.q(n173));
  or_bb g426(.a(n416_1),.b(n424_1),.q(_w_1676));
  bfr _b_882(.a(_w_1337),.q(_w_1338));
  bfr _b_1257(.a(_w_1712),.q(_w_1713));
  or_bb g252(.a(n203_3),.b(n237_1),.q(_w_1675));
  or_bb g451(.a(n433_1),.b(n434_1),.q(_w_2479));
  bfr _b_899(.a(_w_1354),.q(_w_1355));
  or_bb g180(.a(n136_1),.b(n179_1),.q(_w_1674));
  or_bb g260(.a(n216_1),.b(n259_0),.q(n260));
  or_bb g101(.a(n81_1),.b(n99_1),.q(_w_1673));
  spl2 g330_s_0(.a(n330),.q0(n330_0),.q1(n330_1));
  and_bi g286(.a(n283),.b(n285_0),.q(n286));
  and_bb g131(.a(n105_0),.b(n130_0),.q(n131));
  bfr _b_1851(.a(_w_2306),.q(_w_2307));
  and_bb g216(.a(n184_0),.b(n215_2),.q(n216));
  and_bb g228(.a(a_0__5),.b(b_2__10),.q(_w_1671));
  bfr _b_1940(.a(_w_2395),.q(_w_2396));
  bfr _b_1157(.a(_w_1612),.q(_w_1613));
  spl2 g246_s_0(.a(n246),.q0(n246_0),.q1(n246_1));
  spl2 g103_s_0(.a(n103),.q0(n103_0),.q1(n103_1));
  bfr _b_996(.a(_w_1451),.q(_w_1452));
  bfr _b_1678(.a(_w_2133),.q(_w_2134));
  or_bb g346(.a(n329_1),.b(n344_1),.q(_w_1670));
  bfr _b_1517(.a(_w_1972),.q(_w_1973));
  or_bb g264(.a(n251_2),.b(n253_1),.q(_w_1669));
  bfr _b_1792(.a(_w_2247),.q(_w_2248));
  spl2 g153_s_0(.a(n153),.q0(n153_0),.q1(n153_1));
  or_bb g185(.a(n170_1),.b(n172_1),.q(_w_1668));
  and_bi g188(.a(n187),.b(n163_1),.q(n188));
  spl2 g188_s_0(.a(n188),.q0(n188_0),.q1(n188_1));
  and_bb g166(.a(a_0__8),.b(b_6__6),.q(n166));
  and_bb g409(.a(n406_0),.b(n408_0),.q(n409));
  or_bb g273(.a(n56_1),.b(n59_1),.q(n273));
  and_bi g157(.a(n155),.b(n156_0),.q(n157));
  spl3L g325_s_0(.a(n325),.q0(n325_0),.q1(n325_1),.q2(_w_1817));
  and_bb g331(.a(n282_1),.b(n326_0),.q(n331));
  or_bb g268(.a(n181_1),.b(n261_1),.q(n268));
  bfr _b_2103(.a(_w_2558),.q(_w_2559));
  bfr _b_2046(.a(_w_2501),.q(_w_2502));
  bfr _b_1737(.a(_w_2192),.q(_w_2193));
  and_bi g244(.a(n243),.b(n242_0),.q(n244));
  and_bb g199(.a(n190_0),.b(n198_0),.q(n199));
  and_bb g401(.a(n397_0),.b(n400_0),.q(n401));
  and_bi g392(.a(n390_1),.b(n389_3),.q(_w_2312));
  and_bb g117(.a(n109_0),.b(n116_0),.q(n117));
  bfr _b_912(.a(_w_1367),.q(_w_1368));
  bfr _b_1921(.a(_w_2376),.q(_w_2377));
  or_bb g202(.a(n200),.b(n201),.q(_w_1666));
  and_bb g226(.a(a_2__7),.b(b_0__8),.q(n226));
  bfr _b_2087(.a(_w_2542),.q(_w_2543));
  spl2 g162_s_0(.a(n162),.q0(n162_0),.q1(n162_1));
  spl2 g117_s_0(.a(n117),.q0(n117_0),.q1(_w_1661));
  and_bi g400(.a(n399),.b(n398_0),.q(n400));
  spl2 g157_s_0(.a(n157),.q0(n157_0),.q1(n157_1));
  and_bb g204(.a(n153_3),.b(n203_0),.q(n204));
  bfr _b_1204(.a(_w_1659),.q(n206));
  spl2 g376_s_0(.a(n376),.q0(n376_0),.q1(n376_1));
  bfr _b_1532(.a(_w_1987),.q(_w_1988));
  bfr _b_1464(.a(_w_1919),.q(_w_1920));
  bfr _b_1309(.a(_w_1764),.q(_w_1765));
  or_bb g82(.a(n65_1),.b(n67_1),.q(_w_1660));
  or_bb g301(.a(n100_1),.b(n103_1),.q(n301));
  bfr _b_943(.a(_w_1398),.q(_w_1399));
  bfr _b_1112(.a(_w_1567),.q(_w_1568));
  or_bb g206(.a(n190_1),.b(n198_1),.q(_w_1659));
  and_bb g35(.a(n32_0),.b(n34_0),.q(n35));
  and_bb g74(.a(n62_5),.b(n73_0),.q(n74));
  and_bb g210(.a(n188_0),.b(n209_0),.q(n210));
  bfr _b_1816(.a(_w_2271),.q(_w_2272));
  spl2 g276_s_0(.a(n276),.q0(n276_0),.q1(n276_1));
  and_bi g253(.a(n252),.b(n238_1),.q(_w_1657));
  spl2 g357_s_0(.a(n357),.q0(n357_0),.q1(n357_1));
  bfr _b_1317(.a(_w_1772),.q(_w_1773));
  spl2 g370_s_0(.a(n370),.q0(n370_0),.q1(n370_1));
  or_bb g211(.a(n188_1),.b(n209_1),.q(_w_1655));
  bfr _b_2069(.a(_w_2524),.q(_w_2525));
  or_bb g343(.a(n330_1),.b(n341_1),.q(_w_2222));
  spl2 g213_s_0(.a(n213),.q0(n213_0),.q1(n213_1));
  bfr _b_1236(.a(_w_1691),.q(_w_1692));
  and_bi g67(.a(n66),.b(n64_0),.q(n67));
  or_bb g214(.a(n210_1),.b(n213_0),.q(n214));
  bfr _b_1360(.a(_w_1815),.q(_w_1816));
  and_bb g384(.a(n381_0),.b(n383_0),.q(n384));
  bfr _b_858(.a(_w_1313),.q(_w_1314));
  and_bb g215(.a(n186_0),.b(n214_0),.q(n215));
  or_bb g217(.a(n184_1),.b(n215_3),.q(_w_1653));
  spl2 g259_s_0(.a(n259),.q0(n259_0),.q1(n259_1));
  or_bb g116(.a(n111_1),.b(n115_0),.q(n116));
  or_bb g221(.a(n204_3),.b(n212_1),.q(_w_1652));
  or_bb g229(.a(n225_1),.b(n226_1),.q(_w_1651));
  bfr _b_1779(.a(_w_2234),.q(_w_2235));
  or_bb g223(.a(n205_1),.b(n207_1),.q(_w_1650));
  bfr _b_1061(.a(_w_1516),.q(_w_1517));
  and_bi g224(.a(n223),.b(n208_1),.q(_w_1642));
  spl2 a_7__s_4(.a(a_7__7),.q0(a_7__8),.q1(_w_1640));
  or_bb g447(.a(n218_1),.b(n258_1),.q(_w_1639));
  bfr _b_1155(.a(_w_1610),.q(_w_1611));
  and_bb g192(.a(a_3__1),.b(b_0__4),.q(n192));
  bfr _b_1100(.a(_w_1555),.q(_w_1556));
  and_bb g227(.a(n225_0),.b(n226_0),.q(n227));
  or_bb g20(.a(n17_1),.b(n18_1),.q(_w_1631));
  or_bb g247(.a(n224_1),.b(n239_1),.q(_w_1630));
  or_bb g69(.a(n64_1),.b(n68_0),.q(n69));
  spl2 g338_s_0(.a(n338),.q0(n338_0),.q1(n338_1));
  and_bb g259(.a(n218_0),.b(n258_0),.q(n259));
  and_bi g344(.a(n343),.b(n342_0),.q(n344));
  spl2 g239_s_0(.a(n239),.q0(n239_0),.q1(n239_1));
  and_bb g238(.a(n203_2),.b(n237_0),.q(n238));
  spl2 g344_s_0(.a(n344),.q0(n344_0),.q1(n344_1));
  and_bi g212(.a(n211),.b(n210_0),.q(n212));
  spl2 g300_s_0(.a(n300),.q0(n300_0),.q1(n300_1));
  or_bb g449(.a(n427_1),.b(n436_1),.q(_w_1629));
  bfr _b_1067(.a(_w_1522),.q(_w_1523));
  or_bb g232(.a(n227_1),.b(n231_0),.q(n232));
  bfr _b_1115(.a(_w_1570),.q(a_5__6));
  spl2 g73_s_0(.a(n73),.q0(n73_0),.q1(n73_1));
  and_bi g454(.a(n453),.b(n257_1),.q(_w_1598));
  bfr _b_1801(.a(_w_2256),.q(_w_2257));
  or_bb g233(.a(n194_1),.b(n196_1),.q(_w_1597));
  and_bi g304(.a(n303),.b(n302_0),.q(n304));
  bfr _b_1018(.a(_w_1473),.q(_w_1474));
  or_bb g243(.a(n220_1),.b(n241_2),.q(_w_1596));
  bfr _b_1830(.a(_w_2285),.q(_w_2286));
  spl2 g179_s_0(.a(n179),.q0(n179_0),.q1(n179_1));
  and_bi g177(.a(n176),.b(n175_0),.q(n177));
  spl2 g424_s_0(.a(n424),.q0(n424_0),.q1(n424_1));
  or_bb g410(.a(n405_1),.b(n409_0),.q(n410));
  and_bb g419(.a(n345_2),.b(n418_0),.q(n419));
  or_bb g120(.a(n109_1),.b(n116_1),.q(_w_1739));
  or_bb g262(.a(n182_1),.b(n260_1),.q(_w_1595));
  bfr _b_1481(.a(_w_1936),.q(a_2__5));
  and_bi g263(.a(n262),.b(n261_0),.q(_w_1572));
  and_bi g341(.a(n340),.b(n339_0),.q(n341));
  bfr _b_1047(.a(_w_1502),.q(_w_1503));
  spl2 g409_s_0(.a(n409),.q0(n409_0),.q1(n409_1));
  or_bb g386(.a(n375_1),.b(n385_1),.q(_w_1571));
  bfr _b_1815(.a(_w_2270),.q(_w_2271));
  bfr _b_1217(.a(_w_1672),.q(n228));
  and_bb g361(.a(n323_0),.b(n360_0),.q(n361));
  spl2 b_4__s_0(.a(_w_2510),.q0(b_4__0),.q1(b_4__1));
  spl3L a_5__s_2(.a(a_5__3),.q0(a_5__4),.q1(a_5__5),.q2(_w_1570));
  spl2 g128_s_0(.a(n128),.q0(n128_0),.q1(n128_1));
  spl2 g78_s_0(.a(n78),.q0(n78_0),.q1(n78_1));
  spl2 g58_s_0(.a(n58),.q0(n58_0),.q1(n58_1));
  or_bb g60(.a(n53_1),.b(n58_1),.q(_w_1569));
  and_bi g267(.a(n266),.b(n256_1),.q(_w_1536));
  spl2 g379_s_0(.a(n379),.q0(n379_0),.q1(_w_1532));
  bfr _b_1515(.a(_w_1970),.q(_w_1971));
  spl3L a_3__s_0(.a(_w_2565),.q0(a_3__0),.q1(a_3__1),.q2(_w_1529));
  bfr _b_1508(.a(_w_1963),.q(n369));
  bfr _b_871(.a(_w_1326),.q(n215_1));
  spl2 b_1__s_0(.a(b_1_),.q0(b_1__0),.q1(b_1__1));
  and_bi g109(.a(n108),.b(n91_1),.q(n109));
  spl2 g95_s_0(.a(n95),.q0(n95_0),.q1(n95_1));
  bfr _b_1693(.a(_w_2148),.q(n402));
  and_bi g313(.a(n311),.b(n312),.q(_w_2103));
  and_bb g156(.a(n153_0),.b(n154_0),.q(n156));
  spl2 g410_s_0(.a(n410),.q0(n410_0),.q1(n410_1));
  and_bb g208(.a(n205_0),.b(n207_0),.q(n208));
  spl2 g286_s_0(.a(n286),.q0(n286_0),.q1(n286_1));
  bfr _b_1135(.a(_w_1590),.q(_w_1591));
  spl2 g86_s_0(.a(n86),.q0(n86_0),.q1(n86_1));
  bfr _b_1837(.a(_w_2292),.q(_w_2293));
  and_bb g24(.a(a_3__3),.b(b_3__0),.q(n24));
  spl2 g85_s_0(.a(n85),.q0(n85_0),.q1(_w_1525));
  bfr _b_2051(.a(_w_2506),.q(_w_2507));
  bfr _b_1840(.a(_w_2295),.q(_w_2296));
  bfr _b_850(.a(_w_1305),.q(_w_1306));
  or_bb g258(.a(n242_1),.b(n257_0),.q(n258));
  spl2 g81_s_0(.a(n81),.q0(n81_0),.q1(n81_1));
  bfr _b_1435(.a(_w_1890),.q(_w_1891));
  and_bi g133(.a(n132),.b(n131_0),.q(n133));
  spl2 g150_s_0(.a(n150),.q0(n150_0),.q1(n150_1));
  bfr _b_1057(.a(_w_1512),.q(_w_1513));
  bfr _b_1862(.a(_w_2317),.q(_w_2318));
  bfr _b_1070(.a(_w_1525),.q(_w_1526));
  spl2 g156_s_0(.a(n156),.q0(n156_0),.q1(_w_1518));
  spl2 g174_s_0(.a(n174),.q0(n174_0),.q1(n174_1));
  spl2 g305_s_0(.a(n305),.q0(n305_0),.q1(n305_1));
  spl2 g347_s_0(.a(n347),.q0(n347_0),.q1(n347_1));
  spl2 g102_s_0(.a(n102),.q0(n102_0),.q1(n102_1));
  bfr _b_1346(.a(_w_1801),.q(_w_1802));
  bfr _b_906(.a(_w_1361),.q(_w_1362));
  spl2 g26_s_0(.a(n26),.q0(n26_0),.q1(n26_1));
  spl2 g129_s_0(.a(n129),.q0(n129_0),.q1(n129_1));
  spl2 g75_s_0(.a(n75),.q0(n75_0),.q1(n75_1));
  bfr _b_1947(.a(_w_2402),.q(_w_2403));
  spl2 g238_s_0(.a(n238),.q0(n238_0),.q1(n238_1));
  bfr _b_2105(.a(_w_2560),.q(_w_2561));
  spl2 g172_s_0(.a(n172),.q0(n172_0),.q1(n172_1));
  spl2 g140_s_0(.a(n140),.q0(n140_0),.q1(n140_1));
  bfr _b_1178(.a(_w_1633),.q(_w_1634));
  spl2 g360_s_0(.a(n360),.q0(n360_0),.q1(n360_1));
  spl2 g111_s_0(.a(n111),.q0(n111_0),.q1(_w_1514));
  bfr _b_2095(.a(_w_2550),.q(_w_2551));
  spl2 g175_s_0(.a(n175),.q0(n175_0),.q1(_w_1510));
  spl2 g270_s_0(.a(n270),.q0(n270_0),.q1(n270_1));
  bfr _b_865(.a(_w_1320),.q(_w_1321));
  bfr _b_1576(.a(_w_2031),.q(_w_2032));
  bfr _b_1542(.a(_w_1997),.q(_w_1998));
  spl2 g64_s_0(.a(n64),.q0(n64_0),.q1(_w_1506));
  spl2 g361_s_0(.a(n361),.q0(n361_0),.q1(n361_1));
  spl2 g145_s_0(.a(n145),.q0(n145_0),.q1(_w_1502));
  spl2 g61_s_0(.a(n61),.q0(n61_0),.q1(n61_1));
  or_bb g320(.a(n316_1),.b(n317_1),.q(_w_2131));
  and_bb g18(.a(a_0__10),.b(b_1__11),.q(n18));
  spl2 g218_s_0(.a(n218),.q0(n218_0),.q1(n218_1));
  spl2 b_1__s_4(.a(b_1__9),.q0(b_1__10),.q1(_w_1495));
  bfr _b_1872(.a(_w_2327),.q(_w_2328));
  spl2 g37_s_0(.a(n37),.q0(n37_0),.q1(n37_1));
  bfr _b_1783(.a(_w_2238),.q(_w_2239));
  spl2 g375_s_0(.a(n375),.q0(n375_0),.q1(n375_1));
  bfr _b_1694(.a(_w_2149),.q(_w_2150));
  spl2 g204_s_1(.a(n204_1),.q0(n204_2),.q1(n204_3));
  bfr _b_930(.a(_w_1385),.q(_w_1386));
  spl2 g227_s_0(.a(n227),.q0(n227_0),.q1(_w_1491));
  and_bi g422(.a(n421),.b(n419_0),.q(n422));
  bfr _b_959(.a(_w_1414),.q(_w_1415));
  spl2 g331_s_0(.a(n331),.q0(n331_0),.q1(_w_1487));
  spl2 g50_s_0(.a(n50),.q0(n50_0),.q1(n50_1));
  bfr _b_1718(.a(_w_2173),.q(n324_1));
  bfr _b_1089(.a(_w_1544),.q(_w_1545));
  spl4L b_7__s_1(.a(b_7__1),.q0(b_7__2),.q1(b_7__3),.q2(b_7__4),.q3(b_7__5));
  or_bb g179(.a(n175_1),.b(n178_0),.q(_w_1824));
  spl2 g40_s_0(.a(n40),.q0(n40_0),.q1(n40_1));
  bfr _b_2044(.a(_w_2499),.q(n285_1));
  spl2 g67_s_0(.a(n67),.q0(n67_0),.q1(n67_1));
  bfr _b_1719(.a(_w_2174),.q(_w_2175));
  bfr _b_1570(.a(_w_2025),.q(n278));
  bfr _b_1060(.a(_w_1515),.q(_w_1516));
  and_bb g191(.a(a_2__0),.b(b_1__4),.q(n191));
  spl2 g47_s_0(.a(n47),.q0(n47_0),.q1(_w_1483));
  or_bb g352(.a(n348_1),.b(n350_1),.q(_w_2236));
  spl2 g69_s_0(.a(n69),.q0(n69_0),.q1(n69_1));
  bfr _b_1599(.a(_w_2054),.q(_w_2055));
  spl2 g46_s_0(.a(n46),.q0(n46_0),.q1(n46_1));
  bfr _b_1889(.a(_w_2344),.q(_w_2345));
  and_bb g197(.a(n194_0),.b(n196_0),.q(n197));
  spl2 g49_s_0(.a(n49),.q0(n49_0),.q1(n49_1));
  bfr _b_1820(.a(_w_2275),.q(n412));
  spl2 g196_s_0(.a(n196),.q0(n196_0),.q1(n196_1));
  spl2 g225_s_0(.a(n225),.q0(n225_0),.q1(n225_1));
  bfr _b_1915(.a(_w_2370),.q(_w_2371));
  spl2 g74_s_0(.a(n74),.q0(n74_0),.q1(_w_1475));
  spl2 g418_s_0(.a(n418),.q0(n418_0),.q1(n418_1));
  spl3L a_0__s_0(.a(_w_2566),.q0(a_0__0),.q1(a_0__1),.q2(a_0__2));
  spl2 a_2__s_0(.a(_w_2519),.q0(a_2__0),.q1(_w_1472));
  spl2 a_2__s_3(.a(a_2__8),.q0(a_2__9),.q1(_w_1469));
  spl2 g52_s_0(.a(n52),.q0(n52_0),.q1(n52_1));
  spl2 g83_s_0(.a(n83),.q0(n83_0),.q1(n83_1));
  spl2 b_2__s_0(.a(_w_2536),.q0(b_2__0),.q1(b_2__1));
  and_bb g54(.a(a_4__4),.b(b_4__4),.q(n54));
  spl2 b_3__s_4(.a(b_3__9),.q0(b_3__10),.q1(b_3__11));
  bfr _b_965(.a(_w_1420),.q(_w_1421));
  spl4L b_3__s_1(.a(b_3__1),.q0(b_3__2),.q1(b_3__3),.q2(b_3__4),.q3(b_3__5));
  spl3L b_2__s_1(.a(b_2__0),.q0(b_2__2),.q1(b_2__3),.q2(b_2__4));
  bfr _b_1021(.a(_w_1476),.q(_w_1477));
  spl2 b_6__s_3(.a(b_6__8),.q0(b_6__9),.q1(b_6__10));
  spl2 b_2__s_3(.a(b_2__8),.q0(b_2__9),.q1(_w_1465));
  spl4L a_4__s_1(.a(a_4__2),.q0(a_4__3),.q1(a_4__4),.q2(a_4__5),.q3(_w_1462));
  bfr _b_2092(.a(_w_2547),.q(_w_2548));
  bfr _b_1316(.a(_w_1771),.q(_w_1772));
  or_bb g195(.a(n191_1),.b(n192_1),.q(_w_2500));
  spl2 a_4__s_2(.a(a_4__6),.q0(a_4__7),.q1(_w_1459));
  spl2 g59_s_0(.a(n59),.q0(n59_0),.q1(n59_1));
  spl2 g290_s_0(.a(n290),.q0(n290_0),.q1(n290_1));
  bfr _b_984(.a(_w_1439),.q(b_4__11));
  spl2 g271_s_0(.a(n271),.q0(n271_0),.q1(n271_1));
  spl2 g133_s_0(.a(n133),.q0(n133_0),.q1(n133_1));
  spl2 g261_s_0(.a(n261),.q0(n261_0),.q1(n261_1));
  bfr _b_1004(.a(_w_1459),.q(_w_1460));
  spl2 b_6__s_0(.a(_w_2553),.q0(b_6__0),.q1(b_6__1));
  bfr _b_841(.a(_w_1296),.q(_w_1297));
  spl2 g253_s_0(.a(n253),.q0(n253_0),.q1(n253_1));
  spl2 b_6__s_4(.a(b_6__10),.q0(b_6__11),.q1(b_6__12));
  spl2 g427_s_0(.a(n427),.q0(n427_0),.q1(n427_1));
  bfr _b_1254(.a(_w_1709),.q(_w_1710));
  spl2 g76_s_0(.a(n76),.q0(n76_0),.q1(_w_1455));
  spl2 g391_s_0(.a(n391),.q0(n391_0),.q1(_w_1441));
  bfr _b_1079(.a(_w_1534),.q(_w_1535));
  spl2 b_4__s_1(.a(b_4__0),.q0(b_4__2),.q1(b_4__3));
  bfr _b_1764(.a(_w_2219),.q(_w_2220));
  bfr _b_1675(.a(_w_2130),.q(n395));
  spl4L b_1__s_1(.a(b_1__1),.q0(b_1__2),.q1(b_1__3),.q2(b_1__4),.q3(_w_1793));
  spl4L b_4__s_2(.a(b_4__1),.q0(b_4__4),.q1(b_4__5),.q2(b_4__6),.q3(_w_1440));
  bfr _b_958(.a(_w_1413),.q(_w_1414));
  spl2 b_4__s_3(.a(b_4__7),.q0(b_4__8),.q1(b_4__9));
  spl2 g119_s_0(.a(n119),.q0(n119_0),.q1(n119_1));
  spl2 b_4__s_4(.a(b_4__9),.q0(b_4__10),.q1(_w_1438));
  bfr _b_1444(.a(_w_1899),.q(n349));
  spl2 b_7__s_0(.a(_w_2520),.q0(b_7__0),.q1(b_7__1));
  bfr _b_980(.a(_w_1435),.q(a_6__9));
  spl2 b_7__s_3(.a(b_7__7),.q0(b_7__8),.q1(b_7__9));
  spl2 g214_s_0(.a(n214),.q0(n214_0),.q1(n214_1));
  spl3L g404_s_0(.a(n404),.q0(n404_0),.q1(n404_1),.q2(n404_2));
  bfr _b_2098(.a(b_6_),.q(_w_2554));
  and_bb g55(.a(a_5__4),.b(b_3__3),.q(n55));
  spl2 a_6__s_3(.a(a_6__5),.q0(a_6__6),.q1(a_6__7));
  spl2 a_6__s_4(.a(a_6__7),.q0(a_6__8),.q1(_w_1431));
  spl2 a_5__s_0(.a(_w_2540),.q0(a_5__0),.q1(_w_1430));
  bfr _b_934(.a(_w_1389),.q(_w_1390));
  bfr _b_1848(.a(_w_2303),.q(_w_2304));
  spl2 a_5__s_1(.a(a_5__1),.q0(a_5__2),.q1(_w_1429));
  spl2 a_5__s_4(.a(a_5__8),.q0(a_5__9),.q1(_w_1427));
  and_bb g277(.a(n271_0),.b(n276_0),.q(n277));
  spl2 g194_s_0(.a(n194),.q0(n194_0),.q1(n194_1));
  bfr _b_1318(.a(_w_1773),.q(_w_1774));
  and_bb g256(.a(n246_0),.b(n255_0),.q(n256));
  spl2 g65_s_0(.a(n65),.q0(n65_0),.q1(n65_1));
  and_bb g295(.a(n293_0),.b(n294_0),.q(n295));
  spl2 g91_s_0(.a(n91),.q0(n91_0),.q1(n91_1));
  bfr _b_1071(.a(_w_1526),.q(_w_1527));
  spl2 b_5__s_0(.a(_w_2541),.q0(b_5__0),.q1(b_5__1));
  bfr _b_1796(.a(_w_2251),.q(_w_2252));
  spl2 b_5__s_1(.a(b_5__0),.q0(b_5__2),.q1(b_5__3));
  spl4L b_5__s_2(.a(b_5__1),.q0(b_5__4),.q1(b_5__5),.q2(b_5__6),.q3(_w_1422));
  spl2 b_5__s_3(.a(b_5__7),.q0(b_5__8),.q1(b_5__9));
  bfr _b_1237(.a(_w_1692),.q(_w_1693));
  and_bb g203(.a(a_0__1),.b(b_3__8),.q(n203));
  spl2 b_5__s_4(.a(b_5__9),.q0(b_5__10),.q1(b_5__11));
  bfr _b_2037(.a(_w_2492),.q(_w_2493));
  bfr _b_1013(.a(_w_1468),.q(b_2__10));
  bfr _b_1027(.a(_w_1482),.q(n74_1));
  spl4L a_3__s_1(.a(a_3__2),.q0(a_3__3),.q1(a_3__4),.q2(a_3__5),.q3(_w_1419));
  spl2 a_0__s_2(.a(a_0__4),.q0(a_0__5),.q1(_w_1926));
  spl2 a_1__s_3(.a(a_1__7),.q0(a_1__8),.q1(_w_1901));
  spl2 g307_s_0(.a(n307),.q0(n307_0),.q1(n307_1));
  spl2 g123_s_0(.a(n123),.q0(n123_0),.q1(n123_1));
  spl2 a_3__s_2(.a(a_3__6),.q0(a_3__7),.q1(_w_1416));
  bfr _b_1330(.a(_w_1785),.q(n62));
  spl2 a_3__s_3(.a(a_3__8),.q0(a_3__9),.q1(_w_1413));
  bfr _b_1049(.a(_w_1504),.q(_w_1505));
  spl2 g36_s_0(.a(n36),.q0(n36_0),.q1(n36_1));
  spl2 b_1__s_3(.a(b_1__7),.q0(b_1__8),.q1(_w_1408));
  spl2 g30_s_0(.a(n30),.q0(n30_0),.q1(n30_1));
  spl2 g384_s_0(.a(n384),.q0(n384_0),.q1(n384_1));
  bfr _b_1245(.a(_w_1700),.q(_w_1701));
  and_bb g19(.a(n17_0),.b(n18_0),.q(_w_2000));
  spl2 g35_s_0(.a(n35),.q0(n35_0),.q1(n35_1));
  bfr _b_993(.a(_w_1448),.q(_w_1449));
  bfr _b_2012(.a(_w_2467),.q(_w_2468));
  spl2 g205_s_0(.a(n205),.q0(n205_0),.q1(n205_1));
  bfr _b_1509(.a(_w_1964),.q(_w_1965));
  spl2 g431_s_0(.a(n431),.q0(n431_0),.q1(_w_1384));
  bfr _b_1093(.a(_w_1548),.q(_w_1549));
  bfr _b_1960(.a(_w_2415),.q(_w_2416));
  spl2 g304_s_0(.a(n304),.q0(n304_0),.q1(n304_1));
  spl2 g363_s_0(.a(n363),.q0(n363_0),.q1(n363_1));
  bfr _b_1037(.a(_w_1492),.q(_w_1493));
  spl3L g255_s_0(.a(n255),.q0(n255_0),.q1(n255_1),.q2(n255_2));
  spl2 g186_s_0(.a(n186),.q0(n186_0),.q1(n186_1));
  spl2 g99_s_0(.a(n99),.q0(n99_0),.q1(n99_1));
  spl2 g109_s_0(.a(n109),.q0(n109_0),.q1(n109_1));
  spl2 g392_s_0(.a(n392),.q0(n392_0),.q1(n392_1));
  bfr _b_833(.a(_w_1288),.q(_w_1289));
  spl2 g165_s_0(.a(n165),.q0(n165_0),.q1(_w_1380));
  bfr _b_1452(.a(_w_1907),.q(_w_1908));
  bfr _b_1051(.a(_w_1506),.q(_w_1507));
  spl2 b_3__s_0(.a(_w_2549),.q0(_w_1379),.q1(b_3__1));
  spl2 g197_s_0(.a(n197),.q0(n197_0),.q1(n197_1));
  spl2 b_3__s_2(.a(b_3__5),.q0(b_3__6),.q1(_w_1377));
  spl2 b_3__s_3(.a(b_3__7),.q0(b_3__8),.q1(b_3__9));
  bfr _b_881(.a(_w_1336),.q(_w_1337));
  bfr _b_1080(.a(_w_1535),.q(n379_1));
  bfr _b_853(.a(_w_1308),.q(_w_1309));
  spl2 g24_s_0(.a(n24),.q0(n24_0),.q1(n24_1));
  bfr _b_1437(.a(_w_1892),.q(n104));
  spl2 g152_s_0(.a(n152),.q0(n152_0),.q1(n152_1));
  and_bi g52(.a(n51),.b(n50_0),.q(n52));
  and_bi g363(.a(n362),.b(n361_0),.q(n363));
  spl2 g390_s_0(.a(n390),.q0(n390_0),.q1(n390_1));
  bfr _b_1411(.a(_w_1866),.q(_w_1867));
  bfr _b_843(.a(_w_1298),.q(_w_1299));
  spl2 g38_s_0(.a(n38),.q0(n38_0),.q1(n38_1));
  and_bi g184(.a(n183),.b(n178_1),.q(n184));
  spl2 g41_s_0(.a(n41),.q0(n41_0),.q1(_w_1373));
  spl4L b_0__s_1(.a(b_0__1),.q0(b_0__2),.q1(b_0__3),.q2(b_0__4),.q3(_w_1372));
  bfr _b_1661(.a(_w_2116),.q(_w_2117));
  spl2 g242_s_0(.a(n242),.q0(n242_0),.q1(_w_1910));
  spl2 b_0__s_2(.a(b_0__5),.q0(b_0__6),.q1(_w_1367));
  bfr _b_878(.a(_w_1333),.q(_w_1334));
  spl2 b_0__s_3(.a(b_0__7),.q0(b_0__8),.q1(_w_1361));
  bfr _b_839(.a(_w_1294),.q(_w_1295));
  bfr _b_1572(.a(_w_2027),.q(_w_2028));
  spl2 g31_s_0(.a(n31),.q0(n31_0),.q1(_w_1357));
  spl2 a_7__s_0(.a(a_7_),.q0(a_7__0),.q1(_w_1353));
  or_bb g382(.a(n376_1),.b(n378_1),.q(_w_1654));
  spl2 a_7__s_3(.a(a_7__5),.q0(a_7__6),.q1(_w_1352));
  bfr _b_1896(.a(_w_2351),.q(_w_2352));
  bfr _b_1271(.a(_w_1726),.q(n275));
  and_bi g107(.a(n106),.b(n98_1),.q(n107));
  spl2 a_7__s_5(.a(a_7__9),.q0(a_7__10),.q1(_w_1349));
  spl2 g39_s_0(.a(n39),.q0(n39_0),.q1(n39_1));
  spl2 g193_s_0(.a(n193),.q0(n193_0),.q1(_w_2308));
  bfr _b_907(.a(_w_1362),.q(_w_1363));
  spl2 g114_s_0(.a(n114),.q0(n114_0),.q1(n114_1));
  spl2 g208_s_0(.a(n208),.q0(n208_0),.q1(n208_1));
  spl2 g154_s_0(.a(n154),.q0(n154_0),.q1(_w_1348));
  bfr _b_1202(.a(_w_1657),.q(_w_1658));
  and_bb g124(.a(n107_0),.b(n123_0),.q(n124));
  spl2 g170_s_0(.a(n170),.q0(n170_0),.q1(n170_1));
  bfr _b_1495(.a(_w_1950),.q(_w_1951));
  spl2 g124_s_0(.a(n124),.q0(n124_0),.q1(_w_1344));
  spl2 g130_s_0(.a(n130),.q0(n130_0),.q1(n130_1));
  spl2 g131_s_0(.a(n131),.q0(n131_0),.q1(_w_1340));
  spl2 g168_s_1(.a(n168_1),.q0(n168_2),.q1(n168_3));
  spl2 g204_s_0(.a(n204),.q0(n204_0),.q1(_w_1331));
  and_bi g450(.a(n449),.b(n437_1),.q(_w_2475));
  spl2 g100_s_0(.a(n100),.q0(n100_0),.q1(_w_1327));
  spl3L g240_s_0(.a(n240),.q0(n240_0),.q1(n240_1),.q2(n240_2));
  bfr _b_1409(.a(_w_1864),.q(_w_1865));
  spl2 g215_s_0(.a(n215),.q0(n215_0),.q1(_w_1322));
  bfr _b_1639(.a(_w_2094),.q(_w_2095));
  bfr _b_1366(.a(_w_1821),.q(_w_1822));
  spl2 g207_s_0(.a(n207),.q0(n207_0),.q1(n207_1));
  spl2 g321_s_0(.a(n321),.q0(n321_0),.q1(n321_1));
  spl2 g63_s_0(.a(n63),.q0(n63_0),.q1(_w_1317));
  or_bb g278(.a(n271_1),.b(n276_1),.q(_w_2025));
  spl2 g148_s_0(.a(n148),.q0(n148_0),.q1(n148_1));
  and_bb g231(.a(n228_0),.b(n230_0),.q(n231));
  spl2 g29_s_0(.a(n29),.q0(n29_0),.q1(n29_1));
  and_bb g71(.a(a_6__8),.b(b_2__9),.q(n71));
  spl2 g396_s_0(.a(n396),.q0(n396_0),.q1(n396_1));
  spl2 g160_s_0(.a(n160),.q0(n160_0),.q1(n160_1));
  spl2 g62_s_1(.a(n62_2),.q0(n62_3),.q1(_w_1315));
  spl2 g163_s_0(.a(n163),.q0(n163_0),.q1(n163_1));
  spl2 g167_s_0(.a(n167),.q0(n167_0),.q1(n167_1));
  bfr _b_1434(.a(_w_1889),.q(_w_1890));
  and_bi g186(.a(n185),.b(n173_1),.q(n186));
  spl2 g98_s_0(.a(n98),.q0(n98_0),.q1(n98_1));
  spl2 g177_s_0(.a(n177),.q0(n177_0),.q1(n177_1));
  and_bb g17(.a(a_1__11),.b(b_0__10),.q(n17));
  bfr _b_953(.a(_w_1408),.q(b_1__9));
  bfr _b_1650(.a(_w_2105),.q(_w_2106));
  spl2 g228_s_0(.a(n228),.q0(n228_0),.q1(n228_1));
  spl2 g178_s_0(.a(n178),.q0(n178_0),.q1(n178_1));
  spl2 g368_s_0(.a(n368),.q0(n368_0),.q1(n368_1));
  spl2 a_6__s_0(.a(a_6_),.q0(a_6__0),.q1(_w_1436));
  bfr _b_1084(.a(_w_1539),.q(_w_1540));
  bfr _b_1308(.a(_w_1763),.q(_w_1764));
  spl2 g181_s_0(.a(n181),.q0(n181_0),.q1(_w_1311));
  bfr _b_1223(.a(_w_1678),.q(_w_1679));
  spl2 g350_s_0(.a(n350),.q0(n350_0),.q1(n350_1));
  bfr _b_1062(.a(_w_1517),.q(n111_1));
  or_bb g417(.a(n324_3),.b(n403_1),.q(_w_2490));
  spl2 g17_s_0(.a(n17),.q0(n17_0),.q1(n17_1));
  bfr _b_917(.a(_w_1372),.q(b_0__5));
  bfr _b_2096(.a(_w_2551),.q(_w_2552));
  bfr _b_1243(.a(_w_1698),.q(_w_1699));
  and_bb g324(.a(a_7__10),.b(b_5__10),.q(n324));
  spl2 g190_s_0(.a(n190),.q0(n190_0),.q1(n190_1));
  spl2 g44_s_0(.a(n44),.q0(n44_0),.q1(n44_1));
  spl2 g25_s_0(.a(n25),.q0(n25_0),.q1(_w_2021));
  bfr _b_1088(.a(_w_1543),.q(_w_1544));
  spl2 g231_s_0(.a(n231),.q0(n231_0),.q1(n231_1));
  bfr _b_1563(.a(_w_2018),.q(_w_2019));
  spl2 g203_s_0(.a(n203),.q0(n203_0),.q1(_w_1300));
  spl2 g203_s_1(.a(n203_1),.q0(n203_2),.q1(n203_3));
  and_bi g28(.a(n27),.b(n25_0),.q(n28));
  spl2 g209_s_0(.a(n209),.q0(n209_0),.q1(n209_1));
  bfr _b_1753(.a(_w_2208),.q(_w_2209));
  bfr _b_1284(.a(_w_1739),.q(n120));
  bfr _b_1252(.a(_w_1707),.q(_w_1708));
  bfr _b_974(.a(_w_1429),.q(a_5__3));
  bfr _b_1758(.a(_w_2213),.q(_w_2214));
  spl2 g353_s_0(.a(n353),.q0(n353_0),.q1(n353_1));
  bfr _b_997(.a(_w_1452),.q(_w_1453));
  spl2 g212_s_0(.a(n212),.q0(n212_0),.q1(n212_1));
  bfr _b_1026(.a(_w_1481),.q(_w_1482));
  spl2 g216_s_0(.a(n216),.q0(n216_0),.q1(_w_1296));
  bfr _b_1772(.a(_w_2227),.q(n350));
  bfr _b_1326(.a(_w_1781),.q(_w_1782));
  bfr _b_1005(.a(_w_1460),.q(_w_1461));
  spl2 g220_s_0(.a(n220),.q0(n220_0),.q1(n220_1));
  spl2 g295_s_0(.a(n295),.q0(n295_0),.q1(_w_1292));
  and_bb g225(.a(a_1__4),.b(b_1__10),.q(n225));
  spl2 g222_s_0(.a(n222),.q0(n222_0),.q1(n222_1));
  spl2 g226_s_0(.a(n226),.q0(n226_0),.q1(n226_1));
  bfr _b_860(.a(_w_1315),.q(_w_1316));
  bfr _b_1485(.a(_w_1940),.q(_w_1941));
  spl2 g184_s_0(.a(n184),.q0(n184_0),.q1(n184_1));
  spl2 g134_s_0(.a(n134),.q0(n134_0),.q1(n134_1));
  and_bb g298(.a(n279_0),.b(n297_0),.q(n298));
  spl2 g230_s_0(.a(n230),.q0(n230_0),.q1(n230_1));
  bfr _b_854(.a(_w_1309),.q(_w_1310));
  bfr _b_1041(.a(_w_1496),.q(_w_1497));
  bfr _b_1390(.a(_w_1845),.q(_w_1846));
  spl2 g107_s_0(.a(n107),.q0(n107_0),.q1(n107_1));
  bfr _b_1953(.a(_w_2408),.q(n147));
  bfr _b_1828(.a(_w_2283),.q(n368));
  and_bb g98(.a(n95_0),.b(n97_0),.q(n98));
  spl2 g234_s_0(.a(n234),.q0(n234_0),.q1(n234_1));
  spl2 g235_s_0(.a(n235),.q0(n235_0),.q1(_w_1288));
  spl2 g151_s_0(.a(n151),.q0(n151_0),.q1(_w_2008));
  bfr _b_845(.a(_w_1300),.q(_w_1301));
  and_bi g347(.a(n346),.b(n345_0),.q(n347));
  spl2 g237_s_0(.a(n237),.q0(n237_0),.q1(n237_1));
  bfr _b_1423(.a(_w_1878),.q(_w_1879));
  and_bi g396(.a(n395),.b(n391_0),.q(_w_1734));
  spl3L g241_s_0(.a(n241),.q0(n241_0),.q1(n241_1),.q2(n241_2));
  bfr _b_834(.a(_w_1289),.q(_w_1290));
  bfr _b_1208(.a(_w_1663),.q(_w_1664));
  and_bb g351(.a(n348_0),.b(n350_0),.q(n351));
  spl2 g56_s_0(.a(n56),.q0(n56_0),.q1(_w_1409));
  bfr _b_835(.a(_w_1290),.q(_w_1291));
  bfr _b_1602(.a(_w_2057),.q(_w_2058));
  bfr _b_837(.a(_w_1292),.q(_w_1293));
  bfr _b_2073(.a(_w_2528),.q(_w_2529));
  bfr _b_1875(.a(_w_2330),.q(_w_2331));
  bfr _b_846(.a(_w_1301),.q(_w_1302));
  spl2 g309_s_0(.a(n309),.q0(n309_0),.q1(_w_1522));
  bfr _b_968(.a(_w_1423),.q(b_5__7));
  spl2 g68_s_0(.a(n68),.q0(n68_0),.q1(n68_1));
  bfr _b_838(.a(_w_1293),.q(_w_1294));
  and_bb g181(.a(n136_0),.b(n179_0),.q(n181));
  bfr _b_847(.a(_w_1302),.q(_w_1303));
  bfr _b_851(.a(_w_1306),.q(_w_1307));
  bfr _b_852(.a(_w_1307),.q(_w_1308));
  and_bb g68(.a(n65_0),.b(n67_0),.q(n68));
  bfr _b_855(.a(_w_1310),.q(n203_1));
  bfr _b_1791(.a(_w_2246),.q(_w_2247));
  bfr _b_849(.a(_w_1304),.q(_w_1305));
  bfr _b_856(.a(_w_1311),.q(_w_1312));
  bfr _b_1885(.a(_w_2340),.q(_w_2341));
  bfr _b_1029(.a(_w_1484),.q(_w_1485));
  spl4L b_6__s_1(.a(b_6__1),.q0(b_6__2),.q1(b_6__3),.q2(b_6__4),.q3(_w_2284));
  bfr _b_857(.a(_w_1312),.q(_w_1313));
  bfr _b_862(.a(_w_1317),.q(n63_1));
  bfr _b_1619(.a(_w_2074),.q(_w_2075));
  bfr _b_864(.a(_w_1319),.q(_w_1320));
  bfr _b_2031(.a(_w_2486),.q(_w_2487));
  bfr _b_1069(.a(_w_1524),.q(n309_1));
  bfr _b_866(.a(_w_1321),.q(n419_1));
  bfr _b_1802(.a(_w_2257),.q(_w_2258));
  bfr _b_1538(.a(_w_1993),.q(_w_1994));
  bfr _b_868(.a(_w_1323),.q(_w_1324));
  and_bi g293(.a(n292),.b(n291_0),.q(n293));
  or_bb g51(.a(n37_1),.b(n49_1),.q(_w_1792));
  bfr _b_869(.a(_w_1324),.q(_w_1325));
  bfr _b_870(.a(_w_1325),.q(_w_1326));
  bfr _b_1731(.a(_w_2186),.q(_w_2187));
  and_bb g153(.a(a_1__0),.b(b_4__5),.q(n153));
  or_bb g348(.a(n291_1),.b(n74_1),.q(n348));
  spl2 g224_s_0(.a(n224),.q0(n224_0),.q1(n224_1));
  bfr _b_876(.a(_w_1331),.q(_w_1332));
  bfr _b_1478(.a(_w_1933),.q(n94));
  bfr _b_877(.a(_w_1332),.q(_w_1333));
  bfr _b_879(.a(_w_1334),.q(_w_1335));
  bfr _b_883(.a(_w_1338),.q(_w_1339));
  or_bb g189(.a(n146_1),.b(n148_1),.q(_w_1667));
  bfr _b_884(.a(_w_1339),.q(n204_1));
  bfr _b_885(.a(_w_1340),.q(_w_1341));
  bfr _b_886(.a(_w_1341),.q(_w_1342));
  bfr _b_887(.a(_w_1342),.q(_w_1343));
  bfr _b_888(.a(_w_1343),.q(n131_1));
  bfr _b_1031(.a(_w_1486),.q(n47_1));
  bfr _b_1383(.a(_w_1838),.q(_w_1839));
  and_bi g416(.a(n415),.b(n409_1),.q(_w_2355));
  and_bb g87(.a(a_5__2),.b(b_1__6),.q(n87));
  spl2 g284_s_1(.a(n284_1),.q0(n284_2),.q1(_w_1404));
  bfr _b_892(.a(_w_1347),.q(n124_1));
  bfr _b_925(.a(_w_1380),.q(_w_1381));
  and_bb g29(.a(n26_0),.b(n28_0),.q(n29));
  bfr _b_1003(.a(_w_1458),.q(n76_1));
  bfr _b_893(.a(_w_1348),.q(n154_1));
  bfr _b_1469(.a(_w_1924),.q(_w_1925));
  bfr _b_895(.a(_w_1350),.q(_w_1351));
  bfr _b_896(.a(_w_1351),.q(a_7__11));
  bfr _b_897(.a(_w_1352),.q(a_7__7));
  bfr _b_901(.a(_w_1356),.q(a_7__1));
  bfr _b_1315(.a(_w_1770),.q(_w_1771));
  bfr _b_902(.a(_w_1357),.q(_w_1358));
  bfr _b_1882(.a(_w_2337),.q(_w_2338));
  bfr _b_1644(.a(_w_2099),.q(n326_1));
  and_bi g81(.a(n80),.b(n79_0),.q(n81));
  bfr _b_903(.a(_w_1358),.q(_w_1359));
  bfr _b_904(.a(_w_1359),.q(_w_1360));
  bfr _b_889(.a(_w_1344),.q(_w_1345));
  bfr _b_909(.a(_w_1364),.q(_w_1365));
  bfr _b_1105(.a(_w_1560),.q(_w_1561));
  bfr _b_972(.a(_w_1427),.q(_w_1428));
  bfr _b_910(.a(_w_1365),.q(_w_1366));
  bfr _b_911(.a(_w_1366),.q(b_0__9));
  or_bb g266(.a(n246_1),.b(n255_2),.q(_w_1884));
  bfr _b_913(.a(_w_1368),.q(_w_1369));
  bfr _b_916(.a(_w_1371),.q(b_0__7));
  spl2 g429_s_0(.a(n429),.q0(n429_0),.q1(n429_1));
  bfr _b_918(.a(_w_1373),.q(_w_1374));
  bfr _b_919(.a(_w_1374),.q(_w_1375));
  bfr _b_920(.a(_w_1375),.q(_w_1376));
  and_bi g279(.a(n278),.b(n277_0),.q(n279));
  spl2 g319_s_0(.a(n319),.q0(n319_0),.q1(n319_1));
  bfr _b_921(.a(_w_1376),.q(n41_1));
  bfr _b_923(.a(_w_1378),.q(b_3__7));
  bfr _b_927(.a(_w_1382),.q(_w_1383));
  bfr _b_1492(.a(_w_1947),.q(n441));
  bfr _b_1392(.a(_w_1847),.q(_w_1848));
  or_bb g323(.a(n318_1),.b(n322_1),.q(_w_2137));
  bfr _b_931(.a(_w_1386),.q(_w_1387));
  spl3L b_6__s_2(.a(b_6__5),.q0(b_6__6),.q1(b_6__7),.q2(b_6__8));
  bfr _b_932(.a(_w_1387),.q(_w_1388));
  bfr _b_933(.a(_w_1388),.q(_w_1389));
  or_bb g94(.a(n43_1),.b(n44_1),.q(_w_1933));
  bfr _b_848(.a(_w_1303),.q(_w_1304));
  bfr _b_1006(.a(_w_1461),.q(a_4__8));
  bfr _b_935(.a(_w_1390),.q(_w_1391));
  spl2 g289_s_0(.a(n289),.q0(n289_0),.q1(n289_1));
  spl2 g32_s_0(.a(n32),.q0(n32_0),.q1(n32_1));
  bfr _b_937(.a(_w_1392),.q(_w_1393));
  and_bi g172(.a(n171),.b(n165_0),.q(n172));
  or_bb g48(.a(n38_1),.b(n46_1),.q(_w_1665));
  bfr _b_938(.a(_w_1393),.q(_w_1394));
  bfr _b_939(.a(_w_1394),.q(_w_1395));
  bfr _b_1668(.a(_w_2123),.q(_w_2124));
  bfr _b_941(.a(_w_1396),.q(_w_1397));
  bfr _b_945(.a(_w_1400),.q(_w_1401));
  bfr _b_1505(.a(_w_1960),.q(s_12_));
  bfr _b_947(.a(_w_1402),.q(_w_1403));
  bfr _b_977(.a(_w_1432),.q(_w_1433));
  bfr _b_1382(.a(_w_1837),.q(_w_1838));
  bfr _b_948(.a(_w_1403),.q(n431_1));
  spl2 g436_s_0(.a(n436),.q0(n436_0),.q1(n436_1));
  bfr _b_949(.a(_w_1404),.q(_w_1405));
  bfr _b_2062(.a(_w_2517),.q(_w_2518));
  bfr _b_1667(.a(_w_2122),.q(s_9_));
  bfr _b_950(.a(_w_1405),.q(_w_1406));
  bfr _b_973(.a(_w_1428),.q(a_5__10));
  bfr _b_1766(.a(_w_2221),.q(n338));
  bfr _b_952(.a(_w_1407),.q(n284_3));
  spl2 g136_s_0(.a(n136),.q0(n136_0),.q1(n136_1));
  bfr _b_955(.a(_w_1410),.q(_w_1411));
  bfr _b_975(.a(_w_1430),.q(a_5__1));
  bfr _b_1015(.a(_w_1470),.q(_w_1471));
  spl2 g164_s_0(.a(n164),.q0(n164_0),.q1(n164_1));
  bfr _b_956(.a(_w_1411),.q(_w_1412));
  bfr _b_1209(.a(_w_1664),.q(n117_1));
  bfr _b_960(.a(_w_1415),.q(a_3__10));
  bfr _b_961(.a(_w_1416),.q(_w_1417));
  bfr _b_1353(.a(_w_1808),.q(_w_1809));
  spl2 g142_s_0(.a(n142),.q0(n142_0),.q1(n142_1));
  bfr _b_962(.a(_w_1417),.q(_w_1418));
  bfr _b_2017(.a(_w_2472),.q(_w_2473));
  bfr _b_963(.a(_w_1418),.q(a_3__8));
  and_bi g205(.a(n202),.b(n204_0),.q(n205));
  bfr _b_971(.a(_w_1426),.q(a_5__12));
  bfr _b_966(.a(_w_1421),.q(a_3__6));
  bfr _b_969(.a(_w_1424),.q(_w_1425));
  bfr _b_976(.a(_w_1431),.q(_w_1432));
  bfr _b_2010(.a(_w_2465),.q(_w_2466));
  bfr _b_1918(.a(_w_2373),.q(_w_2374));
  bfr _b_1685(.a(_w_2140),.q(_w_2141));
  bfr _b_979(.a(_w_1434),.q(_w_1435));
  bfr _b_1800(.a(_w_2255),.q(_w_2256));
  spl2 g419_s_0(.a(n419),.q0(n419_0),.q1(_w_1318));
  bfr _b_982(.a(_w_1437),.q(a_6__1));
  bfr _b_1197(.a(_w_1652),.q(n221));
  or_bb g362(.a(n323_1),.b(n360_1),.q(_w_2100));
  bfr _b_985(.a(_w_1440),.q(b_4__7));
  bfr _b_1930(.a(_w_2385),.q(n421));
  bfr _b_987(.a(_w_1442),.q(_w_1443));
  bfr _b_988(.a(_w_1443),.q(_w_1444));
  bfr _b_989(.a(_w_1444),.q(_w_1445));
  bfr _b_840(.a(_w_1295),.q(n295_1));
  bfr _b_991(.a(_w_1446),.q(_w_1447));
  bfr _b_992(.a(_w_1447),.q(_w_1448));
  spl2 g332_s_0(.a(n332),.q0(n332_0),.q1(n332_1));
  bfr _b_1001(.a(_w_1456),.q(_w_1457));
  bfr _b_994(.a(_w_1449),.q(_w_1450));
  bfr _b_995(.a(_w_1450),.q(_w_1451));
  and_bb g44(.a(a_2__6),.b(b_5__3),.q(n44));
  bfr _b_998(.a(_w_1453),.q(_w_1454));
  bfr _b_1002(.a(_w_1457),.q(_w_1458));
  spl2 a_5__s_5(.a(a_5__10),.q0(a_5__11),.q1(_w_1424));
  bfr _b_1007(.a(_w_1462),.q(_w_1463));
  bfr _b_1008(.a(_w_1463),.q(_w_1464));
  bfr _b_1009(.a(_w_1464),.q(a_4__6));
  bfr _b_1010(.a(_w_1465),.q(_w_1466));
  bfr _b_986(.a(_w_1441),.q(_w_1442));
  bfr _b_1011(.a(_w_1466),.q(_w_1467));
  bfr _b_1487(.a(_w_1942),.q(_w_1943));
  bfr _b_1012(.a(_w_1467),.q(_w_1468));
  bfr _b_1486(.a(_w_1941),.q(_w_1942));
  bfr _b_1014(.a(_w_1469),.q(_w_1470));
  bfr _b_1016(.a(_w_1471),.q(a_2__10));
  bfr _b_1331(.a(_w_1786),.q(n245));
  or_bb g239(.a(n235_1),.b(n238_0),.q(n239));
  bfr _b_946(.a(_w_1401),.q(_w_1402));
  bfr _b_1017(.a(_w_1472),.q(_w_1473));
  bfr _b_1019(.a(_w_1474),.q(a_2__1));
  bfr _b_1020(.a(_w_1475),.q(_w_1476));
  bfr _b_1054(.a(_w_1509),.q(n64_1));
  or_bb g159(.a(n152_1),.b(n157_1),.q(_w_1656));
  bfr _b_1022(.a(_w_1477),.q(_w_1478));
  and_bb g284(.a(a_6__4),.b(b_4__6),.q(n284));
  bfr _b_1032(.a(_w_1487),.q(_w_1488));
  bfr _b_1034(.a(_w_1489),.q(_w_1490));
  bfr _b_1035(.a(_w_1490),.q(n331_1));
  bfr _b_1036(.a(_w_1491),.q(_w_1492));
  bfr _b_1285(.a(_w_1740),.q(_w_1741));
  bfr _b_1038(.a(_w_1493),.q(_w_1494));
  bfr _b_1044(.a(_w_1499),.q(_w_1500));
  bfr _b_1046(.a(_w_1501),.q(b_1__11));
  bfr _b_1476(.a(_w_1931),.q(_w_1932));
  spl2 g43_s_0(.a(n43),.q0(n43_0),.q1(n43_1));
  spl2 g280_s_0(.a(n280),.q0(n280_0),.q1(n280_1));
  bfr _b_1048(.a(_w_1503),.q(_w_1504));
  bfr _b_1050(.a(_w_1505),.q(n145_1));
  or_bb g139(.a(n119_1),.b(n121_1),.q(_w_1905));
  bfr _b_954(.a(_w_1409),.q(_w_1410));
  bfr _b_936(.a(_w_1391),.q(_w_1392));
  bfr _b_1053(.a(_w_1508),.q(_w_1509));
  bfr _b_1055(.a(_w_1510),.q(_w_1511));
  bfr _b_1296(.a(_w_1751),.q(_w_1752));
  spl2 g378_s_0(.a(n378),.q0(n378_0),.q1(n378_1));
  bfr _b_1058(.a(_w_1513),.q(n175_1));
  bfr _b_1185(.a(_w_1640),.q(_w_1641));
  bfr _b_1059(.a(_w_1514),.q(_w_1515));
  bfr _b_1065(.a(_w_1520),.q(_w_1521));
  bfr _b_978(.a(_w_1433),.q(_w_1434));
  bfr _b_1107(.a(_w_1562),.q(_w_1563));
  bfr _b_1066(.a(_w_1521),.q(n156_1));
  bfr _b_1072(.a(_w_1527),.q(_w_1528));
  bfr _b_1184(.a(_w_1639),.q(n447));
  bfr _b_1074(.a(_w_1529),.q(_w_1530));
  bfr _b_1803(.a(_w_2258),.q(_w_2259));
  bfr _b_1075(.a(_w_1530),.q(_w_1531));
  bfr _b_1438(.a(_w_1893),.q(n340));
  bfr _b_1078(.a(_w_1533),.q(_w_1534));
  bfr _b_1081(.a(_w_1536),.q(_w_1537));
  bfr _b_1090(.a(_w_1545),.q(_w_1546));
  bfr _b_1094(.a(_w_1549),.q(_w_1550));
  bfr _b_900(.a(_w_1355),.q(_w_1356));
  bfr _b_1095(.a(_w_1550),.q(_w_1551));
  bfr _b_1096(.a(_w_1551),.q(_w_1552));
  bfr _b_1780(.a(_w_2235),.q(n36));
  bfr _b_1097(.a(_w_1552),.q(_w_1553));
  bfr _b_2022(.a(_w_2477),.q(_w_2478));
  bfr _b_1954(.a(_w_2409),.q(_w_2410));
  bfr _b_1099(.a(_w_1554),.q(_w_1555));
  bfr _b_1101(.a(_w_1556),.q(_w_1557));
  bfr _b_1941(.a(_w_2396),.q(_w_2397));
  bfr _b_1102(.a(_w_1557),.q(_w_1558));
  bfr _b_1104(.a(_w_1559),.q(_w_1560));
  bfr _b_1558(.a(_w_2013),.q(_w_2014));
  bfr _b_1108(.a(_w_1563),.q(_w_1564));
endmodule
